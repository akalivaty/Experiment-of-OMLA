//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1191, new_n1192, new_n1194, new_n1195,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n202), .A2(new_n203), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n203), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n210), .B(new_n217), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT64), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  NAND2_X1  g0040(.A1(new_n201), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n203), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n214), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n253), .B1(new_n250), .B2(new_n214), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n215), .A2(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n224), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n260), .A2(KEYINPUT11), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(new_n252), .B2(new_n254), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(G68), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n264), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n203), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT12), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n260), .A2(KEYINPUT11), .ZN(new_n273));
  AND4_X1   g0073(.A1(new_n261), .A2(new_n269), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n275), .A2(new_n278), .A3(new_n219), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n278), .A2(new_n281), .A3(G274), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n284), .B(new_n287), .C1(G232), .C2(new_n286), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G97), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n281), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT13), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n274), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n291), .B(KEYINPUT13), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT14), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n293), .A2(new_n300), .A3(G169), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n293), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n300), .B1(new_n293), .B2(G169), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n274), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n299), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n284), .A2(G1698), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT66), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(new_n219), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT69), .ZN(new_n311));
  INV_X1    g0111(.A(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT3), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n286), .A2(G232), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n311), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n284), .A2(KEYINPUT69), .A3(G232), .A4(new_n286), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n318), .B(new_n319), .C1(new_n226), .C2(new_n284), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n275), .B1(new_n310), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n275), .A2(new_n278), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n282), .B1(G244), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G190), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n266), .A2(G77), .A3(new_n268), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT15), .B(G87), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n258), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  INV_X1    g0130(.A(new_n256), .ZN(new_n331));
  OAI22_X1  g0131(.A1(new_n330), .A2(new_n331), .B1(new_n215), .B2(new_n224), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n255), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n270), .A2(new_n224), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n327), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(G200), .B2(new_n324), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n325), .A2(new_n302), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n335), .B1(new_n324), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n256), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT68), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n330), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n344), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n343), .B1(new_n348), .B2(new_n258), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n255), .B1(new_n201), .B2(new_n270), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n266), .A2(G50), .A3(new_n268), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n352), .B(KEYINPUT9), .ZN(new_n353));
  INV_X1    g0153(.A(G223), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n309), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n284), .A2(G222), .A3(new_n286), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n224), .B2(new_n284), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n275), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n282), .B1(G226), .B2(new_n322), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT65), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G200), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n353), .B(new_n362), .C1(new_n294), .C2(new_n361), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT10), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT70), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n363), .B(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n361), .A2(new_n339), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n352), .C1(G179), .C2(new_n361), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n307), .A2(new_n342), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n354), .A2(new_n286), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n285), .A2(G1698), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT71), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n313), .A2(new_n315), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n312), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n312), .A2(new_n220), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n275), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n281), .A2(G232), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n281), .A2(new_n380), .A3(KEYINPUT75), .A4(G232), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n282), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n379), .A2(new_n385), .A3(new_n294), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n379), .A2(new_n385), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(G200), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n345), .A2(new_n347), .A3(new_n268), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n265), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n346), .B1(new_n344), .B2(new_n330), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n264), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT74), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT74), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n394), .B1(new_n264), .B2(new_n391), .C1(new_n265), .C2(new_n389), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G58), .A2(G68), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT72), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(G58), .A3(G68), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n400), .A3(new_n211), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G20), .ZN(new_n402));
  INV_X1    g0202(.A(G159), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n402), .B1(new_n403), .B2(new_n331), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT7), .B1(new_n316), .B2(new_n215), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n406), .B(G20), .C1(new_n313), .C2(new_n315), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT73), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n406), .B1(new_n284), .B2(G20), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n316), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n203), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT73), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT16), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n375), .A2(new_n215), .A3(new_n376), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT7), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n375), .A2(new_n406), .A3(new_n215), .A4(new_n376), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(G68), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n331), .A2(new_n403), .ZN(new_n421));
  AOI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(new_n401), .C2(G20), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n255), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n388), .B(new_n396), .C1(new_n415), .C2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n421), .B1(new_n401), .B2(G20), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n413), .B2(KEYINPUT73), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n409), .B(new_n203), .C1(new_n411), .C2(new_n412), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n420), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n255), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n419), .B2(new_n422), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n431), .A2(new_n433), .B1(new_n393), .B2(new_n395), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n339), .B1(new_n379), .B2(new_n385), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(G179), .B2(new_n387), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT18), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n396), .B1(new_n415), .B2(new_n424), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  INV_X1    g0239(.A(new_n436), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n434), .A2(KEYINPUT17), .A3(new_n388), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n427), .A2(new_n437), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n370), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n281), .A2(G274), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n277), .A2(G1), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(new_n221), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n445), .A2(new_n446), .B1(new_n281), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G116), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n375), .A2(new_n376), .ZN(new_n451));
  NOR2_X1   g0251(.A1(G238), .A2(G1698), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n225), .B2(G1698), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n450), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n448), .B1(new_n454), .B2(new_n281), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT78), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(KEYINPUT78), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n302), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n455), .B(new_n457), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(G169), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT79), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n451), .A2(new_n215), .A3(G68), .ZN(new_n464));
  NOR2_X1   g0264(.A1(G97), .A2(G107), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n465), .A2(new_n220), .B1(new_n289), .B2(new_n215), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT19), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n258), .A2(KEYINPUT19), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n464), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n471), .A2(new_n255), .B1(new_n270), .B2(new_n328), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n267), .A2(G33), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n266), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n328), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n462), .A2(new_n463), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n460), .B(KEYINPUT79), .C1(G169), .C2(new_n461), .ZN(new_n479));
  INV_X1    g0279(.A(new_n461), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G200), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n475), .A2(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n472), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n461), .B2(G190), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n478), .A2(new_n479), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n451), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n227), .A2(G1698), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(G257), .B2(G1698), .ZN(new_n488));
  XOR2_X1   g0288(.A(KEYINPUT80), .B(G303), .Z(new_n489));
  OAI22_X1  g0289(.A1(new_n486), .A2(new_n488), .B1(new_n284), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n275), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT5), .B(G41), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n275), .B1(new_n446), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G270), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(G20), .B1(G33), .B2(G283), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G33), .B2(new_n469), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(new_n251), .C1(new_n215), .C2(G116), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT20), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G116), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n263), .A2(G20), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n500), .B(new_n502), .C1(new_n474), .C2(new_n501), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n492), .A2(new_n446), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n445), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n495), .A2(new_n503), .A3(G179), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n491), .A2(new_n506), .A3(new_n494), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n503), .A2(new_n508), .A3(KEYINPUT21), .A4(G169), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n503), .B1(G200), .B2(new_n508), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n294), .B2(new_n508), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n503), .A2(G169), .A3(new_n508), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n510), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G250), .A2(G1698), .ZN(new_n517));
  INV_X1    g0317(.A(G257), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(G1698), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n451), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G294), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n312), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n275), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n493), .A2(G264), .B1(new_n505), .B2(new_n445), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(KEYINPUT81), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT81), .B1(new_n525), .B2(new_n526), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n528), .A2(new_n529), .A3(new_n339), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(new_n526), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n302), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n226), .A2(KEYINPUT23), .A3(G20), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT23), .B1(new_n226), .B2(G20), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(G20), .B2(new_n449), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n284), .A2(new_n215), .A3(G87), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n451), .A2(KEYINPUT22), .A3(new_n215), .A4(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT24), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n542), .A3(new_n539), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n432), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n264), .A2(G107), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n545), .B(KEYINPUT25), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n474), .B2(new_n226), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n530), .A2(new_n532), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n221), .B2(new_n286), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n284), .ZN(new_n551));
  INV_X1    g0351(.A(G283), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n312), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n225), .A2(G1698), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT4), .B1(new_n451), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n275), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n493), .A2(G257), .B1(new_n505), .B2(new_n445), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n339), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n493), .A2(G257), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n506), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n557), .A2(KEYINPUT76), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n302), .A4(new_n556), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n474), .A2(new_n469), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n469), .A2(new_n226), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(new_n465), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n226), .A2(KEYINPUT6), .A3(G97), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n574));
  OAI21_X1  g0374(.A(G107), .B1(new_n405), .B2(new_n407), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n432), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n264), .A2(G97), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n568), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT77), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR4_X1   g0380(.A1(new_n568), .A2(new_n576), .A3(KEYINPUT77), .A4(new_n577), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n567), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n544), .A2(new_n547), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT81), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n531), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(G190), .B1(new_n585), .B2(new_n527), .ZN(new_n586));
  INV_X1    g0386(.A(new_n531), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n583), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n558), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G190), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n563), .A2(new_n564), .A3(new_n556), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G200), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n593), .A3(new_n578), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n548), .A2(new_n582), .A3(new_n589), .A4(new_n594), .ZN(new_n595));
  AND4_X1   g0395(.A1(new_n444), .A2(new_n485), .A3(new_n516), .A4(new_n595), .ZN(G372));
  OAI21_X1  g0396(.A(new_n306), .B1(new_n303), .B2(new_n304), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n338), .A2(new_n340), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n299), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n425), .A2(new_n426), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT17), .B1(new_n434), .B2(new_n388), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n437), .A2(new_n441), .A3(KEYINPUT82), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT82), .B1(new_n437), .B2(new_n441), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n367), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n607), .A2(new_n369), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT26), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n576), .A2(new_n577), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT77), .B1(new_n610), .B2(new_n568), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n578), .A2(new_n579), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n566), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n485), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n477), .A2(new_n472), .B1(new_n339), .B2(new_n455), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n460), .ZN(new_n616));
  INV_X1    g0416(.A(new_n483), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n455), .A2(G200), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n617), .B(new_n618), .C1(new_n480), .C2(new_n294), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n566), .A2(new_n578), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n619), .A2(new_n609), .A3(new_n616), .A4(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n548), .A2(new_n515), .A3(new_n510), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n582), .A2(new_n589), .A3(new_n619), .A4(new_n594), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n616), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n444), .B1(new_n614), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n608), .A2(new_n625), .ZN(G369));
  AND2_X1   g0426(.A1(new_n510), .A2(new_n515), .ZN(new_n627));
  INV_X1    g0427(.A(new_n263), .ZN(new_n628));
  OR3_X1    g0428(.A1(new_n628), .A2(KEYINPUT27), .A3(G20), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT27), .B1(new_n628), .B2(G20), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(G213), .ZN(new_n631));
  INV_X1    g0431(.A(G343), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n503), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n516), .B2(new_n634), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT83), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n548), .A2(new_n589), .ZN(new_n638));
  INV_X1    g0438(.A(new_n633), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n583), .A2(new_n639), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n638), .A2(new_n640), .B1(new_n548), .B2(new_n639), .ZN(new_n641));
  XOR2_X1   g0441(.A(new_n641), .B(KEYINPUT84), .Z(new_n642));
  NAND3_X1  g0442(.A1(new_n637), .A2(G330), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT85), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n548), .A2(new_n633), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n627), .A2(new_n633), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n645), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(G399));
  INV_X1    g0448(.A(new_n208), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(G41), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n465), .A2(new_n220), .A3(new_n501), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n650), .A2(new_n651), .A3(new_n267), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n213), .B2(new_n650), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT28), .Z(new_n654));
  INV_X1    g0454(.A(KEYINPUT29), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n655), .B(new_n639), .C1(new_n614), .C2(new_n624), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n478), .A2(new_n479), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n481), .A2(new_n484), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n609), .A3(new_n659), .A4(new_n613), .ZN(new_n660));
  INV_X1    g0460(.A(new_n594), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n613), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n548), .A2(new_n510), .A3(new_n515), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(new_n589), .A4(new_n619), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n619), .A2(new_n616), .A3(new_n620), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n660), .A2(new_n664), .A3(new_n616), .A4(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n655), .B1(new_n667), .B2(new_n639), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n657), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n595), .A2(new_n485), .A3(new_n516), .A4(new_n639), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n461), .A2(new_n495), .A3(new_n532), .A4(new_n590), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n587), .A2(new_n456), .A3(G179), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n592), .A2(new_n508), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n672), .A2(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n532), .A2(new_n495), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n677), .A2(KEYINPUT30), .A3(new_n461), .A4(new_n590), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n639), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT31), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n633), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(KEYINPUT86), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT86), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n679), .B2(KEYINPUT31), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n671), .A2(new_n680), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n670), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n654), .B1(new_n689), .B2(G1), .ZN(G364));
  NOR2_X1   g0490(.A1(new_n262), .A2(G20), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n267), .B1(new_n691), .B2(G45), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n650), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(G13), .A2(G33), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G20), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n214), .B1(G20), .B2(new_n339), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n451), .A2(new_n649), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT87), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n213), .A2(new_n277), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n703), .B(new_n704), .C1(new_n277), .C2(new_n245), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n649), .A2(new_n316), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n706), .A2(G355), .B1(new_n501), .B2(new_n649), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n701), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n297), .A2(G179), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(G20), .A3(G190), .ZN(new_n710));
  INV_X1    g0510(.A(G303), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n316), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n215), .A2(new_n302), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G200), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G190), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  XOR2_X1   g0516(.A(KEYINPUT33), .B(G317), .Z(new_n717));
  NOR2_X1   g0517(.A1(new_n714), .A2(new_n294), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G326), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n716), .A2(new_n717), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G179), .A2(G200), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n215), .B1(new_n722), .B2(G190), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n712), .B(new_n721), .C1(G294), .C2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n709), .A2(G20), .A3(new_n294), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT90), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n713), .B(KEYINPUT88), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n294), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI22_X1  g0535(.A1(G283), .A2(new_n731), .B1(new_n735), .B2(G322), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G190), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n722), .A2(G20), .A3(new_n294), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT89), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT89), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n739), .A2(G311), .B1(new_n744), .B2(G329), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n725), .A2(new_n736), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n731), .A2(G107), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n747), .B(new_n284), .C1(new_n220), .C2(new_n710), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT91), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n715), .A2(G68), .B1(new_n718), .B2(G50), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n224), .B2(new_n738), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(G58), .B2(new_n735), .ZN(new_n752));
  OR3_X1    g0552(.A1(new_n743), .A2(KEYINPUT32), .A3(new_n403), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n723), .B(KEYINPUT92), .Z(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G97), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT32), .B1(new_n743), .B2(new_n403), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n752), .A2(new_n753), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n746), .B1(new_n749), .B2(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n695), .B(new_n708), .C1(new_n758), .C2(new_n699), .ZN(new_n759));
  INV_X1    g0559(.A(new_n698), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n637), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n637), .A2(G330), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n695), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n637), .A2(G330), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n761), .B1(new_n763), .B2(new_n764), .ZN(G396));
  NOR2_X1   g0565(.A1(new_n699), .A2(new_n696), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n694), .B1(G77), .B2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT93), .Z(new_n769));
  INV_X1    g0569(.A(new_n710), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n284), .B1(new_n770), .B2(G107), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n771), .B1(new_n719), .B2(new_n711), .C1(new_n552), .C2(new_n716), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n739), .A2(G116), .B1(new_n744), .B2(G311), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n731), .A2(G87), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n773), .B(new_n774), .C1(new_n521), .C2(new_n734), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n772), .B(new_n775), .C1(G97), .C2(new_n754), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n451), .B1(new_n202), .B2(new_n723), .C1(new_n201), .C2(new_n710), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n731), .A2(G68), .ZN(new_n778));
  INV_X1    g0578(.A(G132), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n778), .B1(new_n779), .B2(new_n743), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n715), .A2(G150), .B1(new_n718), .B2(G137), .ZN(new_n781));
  INV_X1    g0581(.A(G143), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n781), .B1(new_n734), .B2(new_n782), .C1(new_n403), .C2(new_n738), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT34), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n777), .B(new_n780), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n776), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n699), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n769), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT95), .Z(new_n791));
  NOR2_X1   g0591(.A1(new_n335), .A2(new_n639), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT96), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n341), .B2(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n598), .B(KEYINPUT96), .C1(new_n335), .C2(new_n639), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n337), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n791), .B1(new_n697), .B2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT97), .Z(new_n798));
  OAI21_X1  g0598(.A(new_n639), .B1(new_n614), .B2(new_n624), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(new_n796), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n695), .B1(new_n800), .B2(new_n688), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n688), .B2(new_n800), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G384));
  OR2_X1    g0604(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n805), .A2(G116), .A3(new_n216), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT36), .Z(new_n808));
  NAND4_X1  g0608(.A1(new_n213), .A2(G77), .A3(new_n400), .A4(new_n398), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n267), .B(G13), .C1(new_n809), .C2(new_n241), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n305), .A2(new_n306), .A3(new_n639), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT101), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT39), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n438), .A2(new_n440), .ZN(new_n816));
  INV_X1    g0616(.A(new_n631), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n438), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT37), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n816), .A2(new_n818), .A3(new_n819), .A4(new_n425), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n390), .A2(new_n392), .ZN(new_n821));
  AOI21_X1  g0621(.A(KEYINPUT16), .B1(new_n419), .B2(new_n428), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n424), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n440), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n817), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n824), .A2(new_n825), .A3(new_n425), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n820), .B1(new_n826), .B2(new_n819), .ZN(new_n827));
  INV_X1    g0627(.A(new_n825), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n443), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT38), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n827), .A2(new_n829), .A3(KEYINPUT38), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n815), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n815), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n425), .B1(new_n434), .B2(new_n436), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n434), .A2(new_n631), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT37), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(KEYINPUT98), .A3(new_n820), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT98), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(KEYINPUT37), .C1(new_n836), .C2(new_n837), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT99), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n600), .B2(new_n601), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n427), .A2(KEYINPUT99), .A3(new_n442), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n837), .B1(new_n606), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n835), .B1(new_n848), .B2(new_n831), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n834), .B1(new_n849), .B2(KEYINPUT100), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT100), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n842), .B2(new_n847), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n852), .B2(new_n835), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n814), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n834), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n427), .A2(KEYINPUT99), .A3(new_n442), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT99), .B1(new_n427), .B2(new_n442), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT82), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n434), .A2(KEYINPUT18), .A3(new_n436), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n437), .A2(new_n441), .A3(KEYINPUT82), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n818), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n839), .A2(new_n841), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n831), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n833), .A2(new_n815), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(KEYINPUT100), .A3(new_n868), .ZN(new_n869));
  AND4_X1   g0669(.A1(new_n814), .A2(new_n853), .A3(new_n855), .A4(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n813), .B1(new_n854), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n796), .B(new_n639), .C1(new_n614), .C2(new_n624), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n341), .A2(new_n639), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n274), .A2(new_n639), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n307), .B(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n832), .A2(new_n833), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n877), .A2(new_n878), .B1(new_n606), .B2(new_n631), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT102), .B1(new_n871), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n869), .A2(new_n855), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT100), .B1(new_n867), .B2(new_n868), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT101), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n853), .A2(new_n814), .A3(new_n855), .A4(new_n869), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n812), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n877), .A2(new_n878), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n606), .A2(new_n631), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT102), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n444), .B1(new_n657), .B2(new_n668), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n608), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n891), .B(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(G330), .ZN(new_n895));
  INV_X1    g0695(.A(new_n875), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n307), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n796), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n682), .A2(KEYINPUT103), .A3(new_n683), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT103), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n679), .B2(KEYINPUT31), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n671), .A2(new_n680), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT40), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n867), .A2(new_n833), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT40), .B1(new_n904), .B2(new_n878), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n444), .A2(new_n902), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n895), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n910), .B2(new_n909), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n894), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n267), .B2(new_n691), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n894), .A2(new_n912), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n811), .B1(new_n914), .B2(new_n915), .ZN(G367));
  OAI21_X1  g0716(.A(new_n700), .B1(new_n208), .B2(new_n328), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n703), .B2(new_n239), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n284), .B1(new_n202), .B2(new_n710), .C1(new_n719), .C2(new_n782), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n731), .A2(G77), .ZN(new_n920));
  INV_X1    g0720(.A(G137), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n920), .B1(new_n921), .B2(new_n743), .C1(new_n738), .C2(new_n201), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n919), .B(new_n922), .C1(G159), .C2(new_n715), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n735), .A2(G150), .B1(new_n754), .B2(G68), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT105), .ZN(new_n925));
  INV_X1    g0725(.A(G317), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n486), .B1(new_n743), .B2(new_n926), .C1(new_n730), .C2(new_n469), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n718), .A2(G311), .B1(G107), .B2(new_n724), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT46), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n770), .A2(G116), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n933), .A2(new_n932), .B1(new_n715), .B2(G294), .ZN(new_n935));
  OAI221_X1 g0735(.A(new_n935), .B1(new_n734), .B2(new_n489), .C1(new_n552), .C2(new_n738), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n930), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n923), .A2(new_n925), .B1(new_n929), .B2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT47), .Z(new_n939));
  AOI211_X1 g0739(.A(new_n695), .B(new_n918), .C1(new_n939), .C2(new_n699), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n483), .A2(new_n633), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n619), .A2(new_n616), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n616), .A2(new_n941), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(new_n698), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n578), .A2(new_n639), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n566), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n662), .B2(new_n946), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n647), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT45), .Z(new_n951));
  NOR2_X1   g0751(.A1(new_n647), .A2(new_n949), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n644), .ZN(new_n955));
  INV_X1    g0755(.A(new_n644), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n951), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n642), .B(new_n646), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n762), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n689), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n650), .B(KEYINPUT41), .Z(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n693), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n642), .A2(new_n646), .A3(new_n949), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT42), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n948), .A2(new_n548), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n633), .B1(new_n968), .B2(new_n582), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n966), .B2(KEYINPUT42), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n942), .A2(new_n943), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n967), .A2(new_n970), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n644), .A2(new_n948), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n945), .B1(new_n965), .B2(new_n976), .ZN(G387));
  OAI22_X1  g0777(.A1(new_n201), .A2(new_n734), .B1(new_n738), .B2(new_n203), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n391), .B2(new_n715), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n754), .A2(new_n476), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n710), .A2(new_n224), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n981), .B(new_n486), .C1(G159), .C2(new_n718), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n731), .A2(G97), .B1(new_n744), .B2(G150), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n979), .A2(new_n980), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(KEYINPUT107), .B(G322), .Z(new_n985));
  AOI22_X1  g0785(.A1(G311), .A2(new_n715), .B1(new_n718), .B2(new_n985), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n734), .B2(new_n926), .C1(new_n489), .C2(new_n738), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT48), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n710), .A2(new_n521), .B1(new_n723), .B2(new_n552), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n987), .B2(new_n988), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(KEYINPUT49), .A3(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n486), .B1(new_n743), .B2(new_n720), .C1(new_n730), .C2(new_n501), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT108), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT49), .B1(new_n989), .B2(new_n991), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n984), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n699), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n706), .A2(new_n651), .B1(new_n226), .B2(new_n649), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n236), .A2(new_n277), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n330), .A2(G50), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n651), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1004), .B(new_n277), .C1(new_n203), .C2(new_n224), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n703), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n999), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n695), .B1(new_n1007), .B2(new_n700), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n998), .B(new_n1008), .C1(new_n642), .C2(new_n760), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n689), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n961), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n650), .B1(new_n961), .B2(new_n1010), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1009), .B1(new_n692), .B2(new_n961), .C1(new_n1011), .C2(new_n1012), .ZN(G393));
  INV_X1    g0813(.A(new_n650), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n961), .A2(new_n1010), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n958), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n1015), .B2(new_n958), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n958), .A2(new_n693), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n703), .A2(new_n248), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n701), .B1(G97), .B2(new_n649), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n695), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n451), .B1(new_n203), .B2(new_n710), .C1(new_n716), .C2(new_n201), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n774), .B1(new_n782), .B2(new_n743), .C1(new_n738), .C2(new_n330), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G77), .C2(new_n754), .ZN(new_n1024));
  INV_X1    g0824(.A(G150), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n734), .A2(new_n403), .B1(new_n1025), .B2(new_n719), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT51), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n316), .B1(new_n552), .B2(new_n710), .C1(new_n716), .C2(new_n489), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n744), .A2(new_n985), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n747), .B(new_n1029), .C1(new_n738), .C2(new_n521), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1028), .B(new_n1030), .C1(G116), .C2(new_n724), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n735), .A2(G311), .B1(G317), .B2(new_n718), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT52), .Z(new_n1033));
  AOI22_X1  g0833(.A1(new_n1024), .A2(new_n1027), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1021), .B1(new_n789), .B2(new_n1034), .C1(new_n949), .C2(new_n760), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1017), .A2(new_n1018), .A3(new_n1035), .ZN(G390));
  OAI21_X1  g0836(.A(new_n812), .B1(new_n874), .B2(new_n876), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n883), .A2(new_n884), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n906), .A2(new_n813), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n667), .A2(new_n639), .A3(new_n796), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n873), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT109), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1040), .A2(KEYINPUT109), .A3(new_n873), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1039), .B1(new_n1045), .B2(new_n876), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n897), .A2(new_n687), .A3(G330), .A4(new_n796), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n897), .A2(new_n902), .A3(G330), .A4(new_n796), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(KEYINPUT110), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n1038), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1049), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(KEYINPUT110), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n693), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n883), .A2(new_n696), .A3(new_n884), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n694), .B1(new_n391), .B2(new_n767), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n284), .B1(new_n716), .B2(new_n921), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G128), .B2(new_n718), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT54), .B(G143), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n739), .A2(new_n1063), .B1(new_n744), .B2(G125), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n754), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1061), .B(new_n1064), .C1(new_n403), .C2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n710), .A2(new_n1025), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT53), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n201), .B2(new_n730), .C1(new_n779), .C2(new_n734), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n735), .A2(G116), .B1(new_n744), .B2(G294), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n778), .C1(new_n469), .C2(new_n738), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n316), .B1(new_n710), .B2(new_n220), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G283), .B2(new_n718), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n226), .B2(new_n716), .C1(new_n1065), .C2(new_n224), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1066), .A2(new_n1069), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1059), .B1(new_n1075), .B2(new_n699), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1057), .A2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT115), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1056), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT113), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT112), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n444), .A2(G330), .A3(new_n902), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n892), .A2(new_n608), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT111), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT111), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n892), .A2(new_n608), .A3(new_n1086), .A4(new_n1083), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n687), .A2(G330), .A3(new_n796), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n876), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n874), .B1(new_n1090), .B2(new_n1049), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n902), .A2(G330), .A3(new_n796), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n876), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(new_n1047), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1091), .B1(new_n1045), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1088), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1082), .B1(new_n1055), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1053), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1038), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1100), .A2(new_n1096), .A3(new_n1082), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1081), .B(new_n650), .C1(new_n1097), .C2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1055), .A2(new_n1096), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1100), .A2(new_n1096), .A3(new_n1101), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT112), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1014), .B1(new_n1109), .B2(new_n1102), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(new_n1081), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1080), .B1(new_n1107), .B2(new_n1111), .ZN(G378));
  NAND2_X1  g0912(.A1(new_n1109), .A2(new_n1102), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1088), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n367), .A2(new_n369), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n352), .A2(new_n817), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1118), .B(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(KEYINPUT117), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n880), .B2(new_n890), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n909), .A2(G330), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n871), .A2(KEYINPUT102), .A3(new_n879), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n889), .B1(new_n885), .B2(new_n888), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1121), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1122), .A2(new_n1124), .A3(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1127), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1123), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1115), .A2(KEYINPUT57), .A3(new_n1129), .A4(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT57), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1129), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1088), .B1(new_n1109), .B2(new_n1102), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1137), .A3(new_n650), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1132), .A2(new_n693), .A3(new_n1129), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n694), .B1(G50), .B2(new_n767), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n735), .A2(G107), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT116), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n486), .A2(new_n276), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n731), .B2(G58), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n739), .A2(new_n476), .B1(new_n744), .B2(G283), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n981), .B1(G97), .B2(new_n715), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n501), .B2(new_n719), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G68), .B2(new_n754), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT58), .ZN(new_n1150));
  AOI21_X1  g0950(.A(G50), .B1(new_n312), .B2(new_n276), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1149), .A2(new_n1150), .B1(new_n1143), .B2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G128), .A2(new_n735), .B1(new_n739), .B2(G137), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n754), .A2(G150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n718), .A2(G125), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n715), .A2(G132), .B1(new_n770), .B2(new_n1063), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n312), .B(new_n276), .C1(new_n730), .C2(new_n403), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G124), .B2(new_n744), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1152), .B1(new_n1150), .B2(new_n1149), .C1(new_n1158), .C2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1140), .B1(new_n1163), .B2(new_n699), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1120), .B2(new_n697), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1139), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1138), .A2(new_n1166), .ZN(G375));
  OAI21_X1  g0967(.A(new_n694), .B1(G68), .B2(new_n767), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n739), .A2(G150), .B1(new_n744), .B2(G128), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n202), .B2(new_n730), .C1(new_n921), .C2(new_n734), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n486), .B1(G159), .B2(new_n770), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G132), .A2(new_n718), .B1(new_n715), .B2(new_n1063), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n1065), .C2(new_n201), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n735), .A2(G283), .B1(new_n744), .B2(G303), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1174), .B(new_n920), .C1(new_n226), .C2(new_n738), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n316), .B1(new_n710), .B2(new_n469), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G294), .B2(new_n718), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n980), .B(new_n1177), .C1(new_n501), .C2(new_n716), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1170), .A2(new_n1173), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1168), .B1(new_n1179), .B2(new_n699), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n897), .B2(new_n697), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1095), .A2(new_n692), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1182), .B2(KEYINPUT119), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(KEYINPUT119), .B2(new_n1182), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n963), .B(KEYINPUT118), .Z(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1096), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1088), .A2(new_n1095), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1189), .ZN(G381));
  OR2_X1    g0990(.A1(G393), .A2(G396), .ZN(new_n1191));
  OR4_X1    g0991(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1191), .ZN(new_n1192));
  OR4_X1    g0992(.A1(G387), .A2(new_n1192), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g0993(.A1(new_n632), .A2(G213), .ZN(new_n1194));
  OR3_X1    g0994(.A1(G375), .A2(G378), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(G407), .A2(G213), .A3(new_n1195), .ZN(G409));
  XNOR2_X1  g0996(.A(G393), .B(G396), .ZN(new_n1197));
  INV_X1    g0997(.A(G390), .ZN(new_n1198));
  AND2_X1   g0998(.A1(G387), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1199), .B2(KEYINPUT124), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(G387), .B(new_n1198), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1135), .A2(new_n1136), .A3(new_n1186), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1139), .A2(new_n1165), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(KEYINPUT120), .B1(new_n1208), .B2(G378), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1138), .A2(G378), .A3(new_n1166), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1115), .A2(new_n1129), .A3(new_n1132), .A4(new_n1185), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1166), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1113), .A2(new_n650), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT113), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1105), .B1(new_n1110), .B2(new_n1081), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1079), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT120), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1212), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1209), .A2(new_n1210), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT121), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT60), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1221), .B(new_n650), .C1(new_n1088), .C2(new_n1095), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1184), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n803), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(G384), .A3(new_n1184), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1219), .A2(new_n1194), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT122), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT63), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT122), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1219), .A2(new_n1232), .A3(new_n1194), .A4(new_n1228), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1219), .A2(new_n1194), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n632), .A2(G213), .A3(G2897), .ZN(new_n1237));
  AOI211_X1 g1037(.A(KEYINPUT123), .B(new_n1237), .C1(new_n1224), .C2(new_n1226), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT123), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1224), .A2(KEYINPUT123), .A3(new_n1226), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1237), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1238), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT61), .B1(new_n1236), .B2(new_n1244), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1205), .A2(new_n1234), .A3(new_n1235), .A4(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT62), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1229), .A2(KEYINPUT62), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1245), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1247), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1204), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1248), .A2(new_n1250), .A3(new_n1247), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1246), .B1(new_n1252), .B2(new_n1253), .ZN(G405));
  NAND2_X1  g1054(.A1(new_n1205), .A2(KEYINPUT126), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G375), .A2(new_n1216), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1210), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1228), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1228), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1204), .A2(new_n1256), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1255), .B(new_n1263), .ZN(G402));
endmodule


