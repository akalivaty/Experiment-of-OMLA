

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n539), .A2(G2104), .ZN(n887) );
  NOR2_X2 U554 ( .A1(n828), .A2(n827), .ZN(n829) );
  NOR2_X2 U555 ( .A1(n699), .A2(n698), .ZN(n705) );
  XNOR2_X1 U556 ( .A(n604), .B(KEYINPUT71), .ZN(n519) );
  INV_X1 U557 ( .A(n733), .ZN(n717) );
  XNOR2_X1 U558 ( .A(n725), .B(KEYINPUT30), .ZN(n726) );
  NOR2_X1 U559 ( .A1(n726), .A2(G168), .ZN(n727) );
  OR2_X2 U560 ( .A1(n688), .A2(n798), .ZN(n733) );
  XNOR2_X1 U561 ( .A(n723), .B(KEYINPUT90), .ZN(n774) );
  XNOR2_X1 U562 ( .A(KEYINPUT65), .B(G651), .ZN(n525) );
  XOR2_X1 U563 ( .A(KEYINPUT15), .B(n609), .Z(n981) );
  NAND2_X1 U564 ( .A1(G101), .A2(n887), .ZN(n540) );
  NOR2_X2 U565 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U566 ( .A1(G89), .A2(n653), .ZN(n520) );
  XOR2_X1 U567 ( .A(KEYINPUT4), .B(n520), .Z(n521) );
  XNOR2_X1 U568 ( .A(n521), .B(KEYINPUT73), .ZN(n523) );
  XOR2_X1 U569 ( .A(KEYINPUT0), .B(G543), .Z(n646) );
  NOR2_X2 U570 ( .A1(n646), .A2(n525), .ZN(n649) );
  NAND2_X1 U571 ( .A1(G76), .A2(n649), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U573 ( .A(KEYINPUT5), .B(n524), .ZN(n533) );
  NOR2_X1 U574 ( .A1(G543), .A2(n525), .ZN(n527) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(KEYINPUT66), .Z(n526) );
  XNOR2_X2 U576 ( .A(n527), .B(n526), .ZN(n652) );
  NAND2_X1 U577 ( .A1(G63), .A2(n652), .ZN(n529) );
  NOR2_X2 U578 ( .A1(G651), .A2(n646), .ZN(n656) );
  NAND2_X1 U579 ( .A1(G51), .A2(n656), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n531) );
  XOR2_X1 U581 ( .A(KEYINPUT6), .B(KEYINPUT74), .Z(n530) );
  XNOR2_X1 U582 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U584 ( .A(KEYINPUT7), .B(n534), .ZN(G168) );
  AND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  NAND2_X1 U586 ( .A1(G113), .A2(n897), .ZN(n536) );
  INV_X1 U587 ( .A(G2105), .ZN(n539) );
  NOR2_X1 U588 ( .A1(G2104), .A2(n539), .ZN(n894) );
  NAND2_X1 U589 ( .A1(G125), .A2(n894), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n544) );
  NOR2_X1 U591 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  XOR2_X1 U592 ( .A(KEYINPUT17), .B(n537), .Z(n625) );
  NAND2_X1 U593 ( .A1(G137), .A2(n625), .ZN(n538) );
  XNOR2_X1 U594 ( .A(n538), .B(KEYINPUT64), .ZN(n542) );
  XOR2_X1 U595 ( .A(KEYINPUT23), .B(n540), .Z(n541) );
  NAND2_X1 U596 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X2 U597 ( .A1(n544), .A2(n543), .ZN(G160) );
  XNOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .ZN(n545) );
  XNOR2_X1 U599 ( .A(n545), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U600 ( .A1(n653), .A2(G85), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G72), .A2(n649), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U603 ( .A1(G60), .A2(n652), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G47), .A2(n656), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U606 ( .A1(n551), .A2(n550), .ZN(G290) );
  XNOR2_X1 U607 ( .A(G2451), .B(G2446), .ZN(n561) );
  XOR2_X1 U608 ( .A(G2430), .B(KEYINPUT104), .Z(n553) );
  XNOR2_X1 U609 ( .A(G2454), .B(G2435), .ZN(n552) );
  XNOR2_X1 U610 ( .A(n553), .B(n552), .ZN(n557) );
  XOR2_X1 U611 ( .A(G2438), .B(KEYINPUT103), .Z(n555) );
  XNOR2_X1 U612 ( .A(G1348), .B(G1341), .ZN(n554) );
  XNOR2_X1 U613 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U614 ( .A(n557), .B(n556), .Z(n559) );
  XNOR2_X1 U615 ( .A(G2443), .B(G2427), .ZN(n558) );
  XNOR2_X1 U616 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U617 ( .A(n561), .B(n560), .ZN(n562) );
  AND2_X1 U618 ( .A1(n562), .A2(G14), .ZN(G401) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U620 ( .A(G57), .ZN(G237) );
  INV_X1 U621 ( .A(G132), .ZN(G219) );
  INV_X1 U622 ( .A(G82), .ZN(G220) );
  NAND2_X1 U623 ( .A1(G65), .A2(n652), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G53), .A2(n656), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n653), .A2(G91), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G78), .A2(n649), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n710) );
  INV_X1 U630 ( .A(n710), .ZN(G299) );
  NAND2_X1 U631 ( .A1(n653), .A2(G88), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G75), .A2(n649), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G62), .A2(n652), .ZN(n572) );
  NAND2_X1 U635 ( .A1(G50), .A2(n656), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U637 ( .A1(n574), .A2(n573), .ZN(G166) );
  NAND2_X1 U638 ( .A1(G64), .A2(n652), .ZN(n576) );
  NAND2_X1 U639 ( .A1(G52), .A2(n656), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n582) );
  NAND2_X1 U641 ( .A1(n653), .A2(G90), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G77), .A2(n649), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(KEYINPUT9), .B(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(KEYINPUT67), .B(n580), .ZN(n581) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(G171) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G102), .A2(n887), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G138), .A2(n625), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G114), .A2(n897), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G126), .A2(n894), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(G164) );
  NAND2_X1 U655 ( .A1(G7), .A2(G661), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n589), .B(KEYINPUT10), .ZN(n590) );
  XNOR2_X1 U657 ( .A(KEYINPUT68), .B(n590), .ZN(G223) );
  INV_X1 U658 ( .A(G223), .ZN(n830) );
  NAND2_X1 U659 ( .A1(n830), .A2(G567), .ZN(n591) );
  XOR2_X1 U660 ( .A(KEYINPUT11), .B(n591), .Z(G234) );
  NAND2_X1 U661 ( .A1(n653), .A2(G81), .ZN(n592) );
  XNOR2_X1 U662 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G68), .A2(n649), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U665 ( .A(KEYINPUT13), .B(n595), .Z(n599) );
  NAND2_X1 U666 ( .A1(G56), .A2(n652), .ZN(n596) );
  XNOR2_X1 U667 ( .A(n596), .B(KEYINPUT14), .ZN(n597) );
  XNOR2_X1 U668 ( .A(n597), .B(KEYINPUT69), .ZN(n598) );
  NOR2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n656), .A2(G43), .ZN(n600) );
  NAND2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n976) );
  INV_X1 U672 ( .A(G860), .ZN(n634) );
  OR2_X1 U673 ( .A1(n976), .A2(n634), .ZN(G153) );
  NAND2_X1 U674 ( .A1(n656), .A2(G54), .ZN(n603) );
  NAND2_X1 U675 ( .A1(G79), .A2(n649), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U677 ( .A1(G66), .A2(n652), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n519), .A2(n605), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n653), .A2(G92), .ZN(n606) );
  XOR2_X1 U680 ( .A(KEYINPUT70), .B(n606), .Z(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U682 ( .A1(n981), .A2(G868), .ZN(n610) );
  XOR2_X1 U683 ( .A(KEYINPUT72), .B(n610), .Z(n612) );
  NAND2_X1 U684 ( .A1(G868), .A2(G301), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(G284) );
  NOR2_X1 U686 ( .A1(G868), .A2(G299), .ZN(n614) );
  INV_X1 U687 ( .A(G868), .ZN(n671) );
  NOR2_X1 U688 ( .A1(G286), .A2(n671), .ZN(n613) );
  NOR2_X1 U689 ( .A1(n614), .A2(n613), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n634), .A2(G559), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n615), .A2(n981), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT76), .ZN(n617) );
  XNOR2_X1 U693 ( .A(KEYINPUT16), .B(n617), .ZN(G148) );
  NOR2_X1 U694 ( .A1(G559), .A2(n671), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n981), .A2(n618), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n619), .B(KEYINPUT77), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n976), .A2(G868), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(G282) );
  NAND2_X1 U699 ( .A1(G99), .A2(n887), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G111), .A2(n897), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n630) );
  NAND2_X1 U702 ( .A1(G123), .A2(n894), .ZN(n624) );
  XNOR2_X1 U703 ( .A(n624), .B(KEYINPUT18), .ZN(n628) );
  BUF_X1 U704 ( .A(n625), .Z(n889) );
  NAND2_X1 U705 ( .A1(G135), .A2(n889), .ZN(n626) );
  XNOR2_X1 U706 ( .A(n626), .B(KEYINPUT78), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n913) );
  XNOR2_X1 U709 ( .A(G2096), .B(n913), .ZN(n632) );
  INV_X1 U710 ( .A(G2100), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(G156) );
  NAND2_X1 U712 ( .A1(G559), .A2(n981), .ZN(n633) );
  XOR2_X1 U713 ( .A(n976), .B(n633), .Z(n668) );
  NAND2_X1 U714 ( .A1(n634), .A2(n668), .ZN(n641) );
  NAND2_X1 U715 ( .A1(G67), .A2(n652), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G55), .A2(n656), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n653), .A2(G93), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G80), .A2(n649), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n670) );
  XOR2_X1 U722 ( .A(n641), .B(n670), .Z(G145) );
  NAND2_X1 U723 ( .A1(G49), .A2(n656), .ZN(n643) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U726 ( .A1(n652), .A2(n644), .ZN(n645) );
  XOR2_X1 U727 ( .A(KEYINPUT79), .B(n645), .Z(n648) );
  NAND2_X1 U728 ( .A1(n646), .A2(G87), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(G288) );
  NAND2_X1 U730 ( .A1(G73), .A2(n649), .ZN(n651) );
  XNOR2_X1 U731 ( .A(KEYINPUT2), .B(KEYINPUT80), .ZN(n650) );
  XNOR2_X1 U732 ( .A(n651), .B(n650), .ZN(n661) );
  NAND2_X1 U733 ( .A1(G61), .A2(n652), .ZN(n655) );
  NAND2_X1 U734 ( .A1(G86), .A2(n653), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U736 ( .A1(G48), .A2(n656), .ZN(n657) );
  XNOR2_X1 U737 ( .A(KEYINPUT81), .B(n657), .ZN(n658) );
  NOR2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(G305) );
  XOR2_X1 U740 ( .A(KEYINPUT82), .B(KEYINPUT19), .Z(n662) );
  XNOR2_X1 U741 ( .A(G290), .B(n662), .ZN(n665) );
  XNOR2_X1 U742 ( .A(G166), .B(G299), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n663), .B(G288), .ZN(n664) );
  XNOR2_X1 U744 ( .A(n665), .B(n664), .ZN(n667) );
  XNOR2_X1 U745 ( .A(G305), .B(n670), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n667), .B(n666), .ZN(n839) );
  XOR2_X1 U747 ( .A(n839), .B(n668), .Z(n669) );
  NOR2_X1 U748 ( .A1(n671), .A2(n669), .ZN(n673) );
  AND2_X1 U749 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U750 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n675), .ZN(n677) );
  XOR2_X1 U754 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n676) );
  XNOR2_X1 U755 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U756 ( .A1(n678), .A2(G2072), .ZN(n679) );
  XNOR2_X1 U757 ( .A(n679), .B(KEYINPUT84), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U761 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G96), .A2(n682), .ZN(n835) );
  NAND2_X1 U763 ( .A1(n835), .A2(G2106), .ZN(n686) );
  NAND2_X1 U764 ( .A1(G69), .A2(G120), .ZN(n683) );
  NOR2_X1 U765 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U766 ( .A1(G108), .A2(n684), .ZN(n836) );
  NAND2_X1 U767 ( .A1(n836), .A2(G567), .ZN(n685) );
  NAND2_X1 U768 ( .A1(n686), .A2(n685), .ZN(n912) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U770 ( .A1(n912), .A2(n687), .ZN(n832) );
  NAND2_X1 U771 ( .A1(n832), .A2(G36), .ZN(G176) );
  INV_X1 U772 ( .A(G166), .ZN(G303) );
  XOR2_X1 U773 ( .A(KEYINPUT32), .B(KEYINPUT98), .Z(n741) );
  XNOR2_X1 U774 ( .A(KEYINPUT96), .B(KEYINPUT29), .ZN(n716) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n799) );
  INV_X1 U776 ( .A(n799), .ZN(n688) );
  NAND2_X1 U777 ( .A1(G160), .A2(G40), .ZN(n798) );
  NAND2_X1 U778 ( .A1(n717), .A2(G2072), .ZN(n689) );
  XNOR2_X1 U779 ( .A(n689), .B(KEYINPUT27), .ZN(n691) );
  XOR2_X1 U780 ( .A(G1956), .B(KEYINPUT92), .Z(n1003) );
  NOR2_X1 U781 ( .A1(n717), .A2(n1003), .ZN(n690) );
  NOR2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n693) );
  INV_X1 U783 ( .A(KEYINPUT93), .ZN(n692) );
  XNOR2_X1 U784 ( .A(n693), .B(n692), .ZN(n709) );
  NOR2_X1 U785 ( .A1(n709), .A2(n710), .ZN(n695) );
  INV_X1 U786 ( .A(KEYINPUT28), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n695), .B(n694), .ZN(n714) );
  INV_X1 U788 ( .A(G1996), .ZN(n941) );
  NOR2_X1 U789 ( .A1(n733), .A2(n941), .ZN(n696) );
  XNOR2_X1 U790 ( .A(n696), .B(KEYINPUT26), .ZN(n699) );
  AND2_X1 U791 ( .A1(n733), .A2(G1341), .ZN(n697) );
  OR2_X1 U792 ( .A1(n697), .A2(n976), .ZN(n698) );
  NAND2_X1 U793 ( .A1(n705), .A2(n981), .ZN(n700) );
  XNOR2_X1 U794 ( .A(n700), .B(KEYINPUT94), .ZN(n704) );
  NOR2_X1 U795 ( .A1(n717), .A2(G1348), .ZN(n702) );
  NOR2_X1 U796 ( .A1(G2067), .A2(n733), .ZN(n701) );
  NOR2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U799 ( .A1(n705), .A2(n981), .ZN(n706) );
  XNOR2_X1 U800 ( .A(n706), .B(KEYINPUT95), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U803 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U805 ( .A(n716), .B(n715), .ZN(n721) );
  NAND2_X1 U806 ( .A1(G1961), .A2(n733), .ZN(n719) );
  XOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .Z(n942) );
  NAND2_X1 U808 ( .A1(n717), .A2(n942), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n722) );
  NOR2_X1 U810 ( .A1(G301), .A2(n722), .ZN(n720) );
  NOR2_X1 U811 ( .A1(n721), .A2(n720), .ZN(n731) );
  AND2_X1 U812 ( .A1(G301), .A2(n722), .ZN(n728) );
  NAND2_X1 U813 ( .A1(n733), .A2(G8), .ZN(n723) );
  NOR2_X1 U814 ( .A1(n774), .A2(G1966), .ZN(n746) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n733), .ZN(n742) );
  NOR2_X1 U816 ( .A1(n746), .A2(n742), .ZN(n724) );
  NAND2_X1 U817 ( .A1(G8), .A2(n724), .ZN(n725) );
  NOR2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n729), .B(KEYINPUT31), .ZN(n730) );
  NOR2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U821 ( .A(n732), .B(KEYINPUT97), .ZN(n744) );
  NAND2_X1 U822 ( .A1(n744), .A2(G286), .ZN(n738) );
  NOR2_X1 U823 ( .A1(n774), .A2(G1971), .ZN(n735) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n736), .A2(G303), .ZN(n737) );
  NAND2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U828 ( .A1(n739), .A2(G8), .ZN(n740) );
  XNOR2_X1 U829 ( .A(n741), .B(n740), .ZN(n748) );
  NAND2_X1 U830 ( .A1(G8), .A2(n742), .ZN(n743) );
  NAND2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U832 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U833 ( .A1(n748), .A2(n747), .ZN(n753) );
  NAND2_X1 U834 ( .A1(G166), .A2(G8), .ZN(n749) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n749), .ZN(n750) );
  NOR2_X1 U836 ( .A1(n753), .A2(n750), .ZN(n751) );
  XNOR2_X1 U837 ( .A(n751), .B(KEYINPUT99), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n752), .A2(n774), .ZN(n769) );
  INV_X1 U839 ( .A(n753), .ZN(n756) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n760) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n754) );
  NOR2_X1 U842 ( .A1(n760), .A2(n754), .ZN(n971) );
  INV_X1 U843 ( .A(KEYINPUT33), .ZN(n759) );
  AND2_X1 U844 ( .A1(n971), .A2(n759), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n767) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n974) );
  INV_X1 U847 ( .A(n774), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n974), .A2(n757), .ZN(n758) );
  AND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n760), .A2(KEYINPUT33), .ZN(n761) );
  NOR2_X1 U851 ( .A1(n774), .A2(n761), .ZN(n763) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n966) );
  INV_X1 U853 ( .A(n966), .ZN(n762) );
  OR2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U855 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U858 ( .A(n770), .B(KEYINPUT100), .ZN(n819) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XNOR2_X1 U860 ( .A(n771), .B(KEYINPUT24), .ZN(n772) );
  XNOR2_X1 U861 ( .A(n772), .B(KEYINPUT91), .ZN(n773) );
  NOR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n817) );
  NAND2_X1 U863 ( .A1(G141), .A2(n889), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G117), .A2(n897), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n887), .A2(G105), .ZN(n777) );
  XOR2_X1 U867 ( .A(KEYINPUT38), .B(n777), .Z(n778) );
  NOR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n894), .A2(G129), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n881) );
  NOR2_X1 U871 ( .A1(G1996), .A2(n881), .ZN(n782) );
  XOR2_X1 U872 ( .A(KEYINPUT101), .B(n782), .Z(n923) );
  NAND2_X1 U873 ( .A1(G1996), .A2(n881), .ZN(n792) );
  NAND2_X1 U874 ( .A1(G131), .A2(n889), .ZN(n783) );
  XOR2_X1 U875 ( .A(KEYINPUT88), .B(n783), .Z(n788) );
  NAND2_X1 U876 ( .A1(G107), .A2(n897), .ZN(n785) );
  NAND2_X1 U877 ( .A1(G119), .A2(n894), .ZN(n784) );
  NAND2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U879 ( .A(KEYINPUT87), .B(n786), .Z(n787) );
  NOR2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n887), .A2(G95), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n882) );
  NAND2_X1 U883 ( .A1(G1991), .A2(n882), .ZN(n791) );
  NAND2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U885 ( .A(KEYINPUT89), .B(n793), .ZN(n820) );
  INV_X1 U886 ( .A(n820), .ZN(n917) );
  NOR2_X1 U887 ( .A1(G1986), .A2(G290), .ZN(n794) );
  NOR2_X1 U888 ( .A1(G1991), .A2(n882), .ZN(n914) );
  NOR2_X1 U889 ( .A1(n794), .A2(n914), .ZN(n795) );
  NOR2_X1 U890 ( .A1(n917), .A2(n795), .ZN(n796) );
  NOR2_X1 U891 ( .A1(n923), .A2(n796), .ZN(n797) );
  XNOR2_X1 U892 ( .A(KEYINPUT39), .B(n797), .ZN(n811) );
  NOR2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n821) );
  XNOR2_X1 U894 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  NAND2_X1 U895 ( .A1(G104), .A2(n887), .ZN(n801) );
  NAND2_X1 U896 ( .A1(G140), .A2(n889), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U898 ( .A(KEYINPUT34), .B(n802), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G116), .A2(n897), .ZN(n804) );
  NAND2_X1 U900 ( .A1(G128), .A2(n894), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U902 ( .A(KEYINPUT85), .B(n805), .ZN(n806) );
  XNOR2_X1 U903 ( .A(KEYINPUT35), .B(n806), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U905 ( .A(KEYINPUT36), .B(n809), .ZN(n902) );
  NOR2_X1 U906 ( .A1(n812), .A2(n902), .ZN(n810) );
  XNOR2_X1 U907 ( .A(n810), .B(KEYINPUT86), .ZN(n933) );
  NAND2_X1 U908 ( .A1(n821), .A2(n933), .ZN(n824) );
  NAND2_X1 U909 ( .A1(n811), .A2(n824), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n812), .A2(n902), .ZN(n813) );
  XNOR2_X1 U911 ( .A(n813), .B(KEYINPUT102), .ZN(n935) );
  NAND2_X1 U912 ( .A1(n814), .A2(n935), .ZN(n815) );
  NAND2_X1 U913 ( .A1(n815), .A2(n821), .ZN(n826) );
  INV_X1 U914 ( .A(n826), .ZN(n816) );
  OR2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n828) );
  XOR2_X1 U917 ( .A(G1986), .B(G290), .Z(n975) );
  NAND2_X1 U918 ( .A1(n820), .A2(n975), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n829), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U925 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT105), .B(n834), .Z(G188) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(n976), .B(KEYINPUT113), .ZN(n838) );
  XNOR2_X1 U936 ( .A(G171), .B(n981), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n841) );
  XNOR2_X1 U938 ( .A(G286), .B(n839), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  NOR2_X1 U940 ( .A1(G37), .A2(n842), .ZN(G397) );
  XOR2_X1 U941 ( .A(G2096), .B(KEYINPUT43), .Z(n844) );
  XNOR2_X1 U942 ( .A(G2090), .B(G2678), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n845), .B(KEYINPUT106), .Z(n847) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT42), .B(G2100), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2078), .B(G2084), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U951 ( .A(G1976), .B(G1956), .Z(n853) );
  XNOR2_X1 U952 ( .A(G1981), .B(G1971), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U954 ( .A(n854), .B(KEYINPUT41), .Z(n856) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1966), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U957 ( .A(G2474), .B(G1961), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U961 ( .A1(G124), .A2(n894), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n887), .A2(G100), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G136), .A2(n889), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G112), .A2(n897), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U968 ( .A1(n867), .A2(n866), .ZN(G162) );
  XNOR2_X1 U969 ( .A(G160), .B(n913), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n868), .B(G162), .ZN(n872) );
  XOR2_X1 U971 ( .A(KEYINPUT110), .B(KEYINPUT112), .Z(n870) );
  XNOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U974 ( .A(n872), .B(n871), .Z(n886) );
  NAND2_X1 U975 ( .A1(G103), .A2(n887), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G139), .A2(n889), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G115), .A2(n897), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G127), .A2(n894), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n877), .ZN(n878) );
  XNOR2_X1 U982 ( .A(KEYINPUT47), .B(n878), .ZN(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n918) );
  XNOR2_X1 U984 ( .A(n918), .B(n881), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U986 ( .A(G164), .B(n884), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n886), .B(n885), .ZN(n904) );
  NAND2_X1 U988 ( .A1(n887), .A2(G106), .ZN(n888) );
  XNOR2_X1 U989 ( .A(KEYINPUT108), .B(n888), .ZN(n892) );
  NAND2_X1 U990 ( .A1(n889), .A2(G142), .ZN(n890) );
  XOR2_X1 U991 ( .A(KEYINPUT109), .B(n890), .Z(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n893), .B(KEYINPUT45), .ZN(n896) );
  NAND2_X1 U994 ( .A1(G130), .A2(n894), .ZN(n895) );
  NAND2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n900) );
  NAND2_X1 U996 ( .A1(G118), .A2(n897), .ZN(n898) );
  XNOR2_X1 U997 ( .A(KEYINPUT107), .B(n898), .ZN(n899) );
  NOR2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(G395) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(G397), .A2(n907), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(n912), .A2(G401), .ZN(n908) );
  XOR2_X1 U1006 ( .A(KEYINPUT114), .B(n908), .Z(n909) );
  NOR2_X1 U1007 ( .A1(G395), .A2(n909), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(n912), .ZN(G319) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  INV_X1 U1012 ( .A(KEYINPUT55), .ZN(n938) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1014 ( .A(KEYINPUT116), .B(n915), .Z(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n931) );
  XOR2_X1 U1016 ( .A(G2072), .B(n918), .Z(n920) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(KEYINPUT50), .B(n921), .ZN(n926) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n924), .Z(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(G2084), .B(G160), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(KEYINPUT115), .B(n927), .ZN(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1030 ( .A(KEYINPUT52), .B(n936), .Z(n937) );
  NAND2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1032 ( .A1(n939), .A2(G29), .ZN(n1022) );
  XOR2_X1 U1033 ( .A(G2084), .B(G34), .Z(n940) );
  XNOR2_X1 U1034 ( .A(KEYINPUT54), .B(n940), .ZN(n959) );
  XNOR2_X1 U1035 ( .A(G2090), .B(G35), .ZN(n957) );
  XNOR2_X1 U1036 ( .A(G32), .B(n941), .ZN(n949) );
  XNOR2_X1 U1037 ( .A(n942), .B(G27), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(G2067), .B(G26), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(KEYINPUT119), .B(n945), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(G1991), .B(G25), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(n950), .B(KEYINPUT117), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(G28), .A2(n951), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(n952), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n960), .B(KEYINPUT120), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n962), .B(n961), .ZN(n964) );
  INV_X1 U1055 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n965), .ZN(n1020) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  XNOR2_X1 U1059 ( .A(G168), .B(G1966), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n968), .B(KEYINPUT57), .ZN(n989) );
  XNOR2_X1 U1062 ( .A(G1956), .B(KEYINPUT124), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(G299), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(G1971), .A2(G303), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n980) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(G1341), .B(n976), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n987) );
  XOR2_X1 U1071 ( .A(G1348), .B(n981), .Z(n982) );
  XNOR2_X1 U1072 ( .A(KEYINPUT122), .B(n982), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(G1961), .B(G301), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(n985), .B(KEYINPUT123), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n1018) );
  INV_X1 U1079 ( .A(G16), .ZN(n1016) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G21), .ZN(n998) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(G23), .B(G1976), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n995) );
  XOR2_X1 U1084 ( .A(G1986), .B(G24), .Z(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(KEYINPUT58), .B(n996), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1011) );
  XOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .Z(n999) );
  XNOR2_X1 U1089 ( .A(G4), .B(n999), .ZN(n1008) );
  XNOR2_X1 U1090 ( .A(G1981), .B(G6), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1002), .B(KEYINPUT126), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(n1003), .B(G20), .Z(n1004) );
  XNOR2_X1 U1095 ( .A(KEYINPUT125), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(n1009), .B(KEYINPUT60), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G5), .B(G1961), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

