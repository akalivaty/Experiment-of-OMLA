//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988;
  INV_X1    g000(.A(KEYINPUT40), .ZN(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT68), .B(G134gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G127gat), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G134gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n204), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n210), .B2(new_n209), .ZN(new_n212));
  INV_X1    g011(.A(G120gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT70), .B1(new_n213), .B2(G113gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n215));
  INV_X1    g014(.A(G113gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(G120gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(G113gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT71), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT71), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n214), .A2(new_n217), .A3(new_n221), .A4(new_n218), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT72), .B(KEYINPUT1), .Z(new_n224));
  INV_X1    g023(.A(G134gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G127gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(new_n208), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n223), .A2(KEYINPUT73), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT73), .B1(new_n223), .B2(new_n228), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n212), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(KEYINPUT80), .B(G162gat), .Z(new_n232));
  INV_X1    g031(.A(G155gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT2), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G155gat), .B(G162gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(G141gat), .B(G148gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT79), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT79), .ZN(new_n238));
  INV_X1    g037(.A(G148gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(G141gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n234), .A2(new_n235), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n235), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(KEYINPUT2), .B2(new_n236), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n231), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n241), .A2(new_n243), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n246), .B(new_n212), .C1(new_n229), .C2(new_n230), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n249), .B(KEYINPUT82), .Z(new_n250));
  OAI21_X1  g049(.A(KEYINPUT39), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT87), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n253), .B(KEYINPUT39), .C1(new_n248), .C2(new_n250), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n247), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n227), .B1(new_n220), .B2(new_n222), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT73), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(KEYINPUT4), .A3(new_n246), .A4(new_n212), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n257), .A2(new_n260), .A3(KEYINPUT83), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n237), .A2(new_n235), .A3(new_n240), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT2), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT80), .B(G162gat), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n268), .B2(G155gat), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n265), .B(new_n243), .C1(new_n266), .C2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT81), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n231), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n263), .A2(new_n264), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n255), .B1(new_n250), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT39), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n276), .A3(new_n250), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT0), .ZN(new_n279));
  XNOR2_X1  g078(.A(G57gat), .B(G85gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n202), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n284), .B(KEYINPUT76), .Z(new_n285));
  INV_X1    g084(.A(G169gat), .ZN(new_n286));
  INV_X1    g085(.A(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT26), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT26), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G183gat), .ZN(new_n294));
  INV_X1    g093(.A(G190gat), .ZN(new_n295));
  OAI22_X1  g094(.A1(new_n289), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT27), .B(G183gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n299), .B2(G190gat), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n298), .B(new_n295), .C1(KEYINPUT67), .C2(KEYINPUT28), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n296), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT25), .B1(new_n288), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n290), .A2(KEYINPUT65), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n290), .A2(KEYINPUT65), .ZN(new_n307));
  NOR4_X1   g106(.A1(new_n304), .A2(new_n305), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  OR2_X1    g108(.A1(new_n309), .A2(KEYINPUT66), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(new_n294), .B2(new_n295), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(KEYINPUT66), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n309), .ZN(new_n316));
  INV_X1    g115(.A(new_n290), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n288), .B2(new_n303), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT64), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n291), .A2(new_n319), .A3(KEYINPUT23), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT64), .B1(new_n288), .B2(new_n303), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n316), .A2(new_n318), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n302), .B1(new_n315), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n285), .B1(new_n325), .B2(KEYINPUT29), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(new_n325), .B2(new_n284), .ZN(new_n328));
  INV_X1    g127(.A(new_n284), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n314), .A2(new_n308), .B1(new_n322), .B2(new_n323), .ZN(new_n330));
  OAI211_X1 g129(.A(KEYINPUT77), .B(new_n329), .C1(new_n330), .C2(new_n302), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n326), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G197gat), .B(G204gat), .ZN(new_n333));
  INV_X1    g132(.A(G211gat), .ZN(new_n334));
  INV_X1    g133(.A(G218gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n333), .B1(KEYINPUT22), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G211gat), .B(G218gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n339), .B(KEYINPUT75), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n325), .A2(new_n285), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n284), .B1(new_n325), .B2(KEYINPUT29), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n346), .B(new_n347), .Z(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT78), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(new_n353), .A3(new_n350), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n349), .A2(new_n350), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n342), .A2(new_n345), .ZN(new_n357));
  INV_X1    g156(.A(new_n348), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n274), .A2(new_n250), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(new_n252), .A3(new_n254), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n362), .A2(KEYINPUT40), .A3(new_n281), .A4(new_n277), .ZN(new_n363));
  INV_X1    g162(.A(new_n281), .ZN(new_n364));
  INV_X1    g163(.A(new_n264), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT83), .B1(new_n257), .B2(new_n260), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n367));
  INV_X1    g166(.A(new_n250), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n273), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n273), .A2(new_n257), .A3(new_n260), .A4(new_n368), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n248), .A2(new_n250), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n371), .A2(KEYINPUT5), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n364), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n283), .A2(new_n360), .A3(new_n363), .A4(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT85), .B1(G228gat), .B2(G233gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n265), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n244), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n271), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n380), .B2(new_n340), .ZN(new_n381));
  NAND3_X1  g180(.A1(KEYINPUT85), .A2(G228gat), .A3(G233gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G22gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n381), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G78gat), .B(G106gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT31), .B(G50gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n384), .A2(KEYINPUT86), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n387), .B(KEYINPUT86), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n375), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n394));
  INV_X1    g193(.A(new_n369), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n263), .A3(new_n264), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n371), .A2(KEYINPUT5), .A3(new_n372), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(new_n281), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n374), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT6), .B(new_n364), .C1(new_n370), .C2(new_n373), .ZN(new_n400));
  INV_X1    g199(.A(new_n357), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT37), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n348), .A2(KEYINPUT38), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n343), .A2(new_n344), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n402), .B1(new_n405), .B2(new_n341), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n332), .A2(new_n340), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n403), .A2(new_n408), .B1(new_n401), .B2(new_n348), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n399), .A2(new_n400), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT88), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n399), .A2(new_n412), .A3(new_n400), .A4(new_n409), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT89), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n414), .B(new_n358), .C1(new_n401), .C2(new_n402), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n402), .B1(new_n342), .B2(new_n345), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT89), .B1(new_n416), .B2(new_n348), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n403), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT38), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT90), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(KEYINPUT90), .A3(KEYINPUT38), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n411), .A2(new_n413), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n393), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n325), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(new_n231), .ZN(new_n426));
  INV_X1    g225(.A(G227gat), .ZN(new_n427));
  INV_X1    g226(.A(G233gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT32), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT33), .B1(new_n426), .B2(new_n429), .ZN(new_n433));
  XNOR2_X1  g232(.A(G71gat), .B(G99gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT74), .ZN(new_n435));
  INV_X1    g234(.A(G15gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(G43gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT34), .B1(new_n426), .B2(new_n429), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n231), .B(new_n325), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT34), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n441), .B(new_n442), .C1(new_n427), .C2(new_n428), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n440), .B(new_n443), .C1(new_n433), .C2(new_n438), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n432), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n432), .A3(new_n446), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n448), .A2(KEYINPUT36), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT36), .B1(new_n448), .B2(new_n449), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n400), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n399), .B2(KEYINPUT84), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n374), .A2(new_n456), .A3(new_n394), .A4(new_n398), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n360), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n424), .B(new_n453), .C1(new_n458), .C2(new_n392), .ZN(new_n459));
  INV_X1    g258(.A(new_n449), .ZN(new_n460));
  NOR4_X1   g259(.A1(new_n460), .A2(new_n447), .A3(new_n389), .A4(new_n391), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n463));
  INV_X1    g262(.A(new_n360), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n399), .A2(new_n400), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n466), .A2(KEYINPUT35), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n463), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT91), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n459), .A2(new_n468), .A3(KEYINPUT91), .ZN(new_n472));
  XNOR2_X1  g271(.A(G113gat), .B(G141gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(G197gat), .ZN(new_n474));
  XOR2_X1   g273(.A(KEYINPUT11), .B(G169gat), .Z(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n476), .B(KEYINPUT12), .Z(new_n477));
  INV_X1    g276(.A(KEYINPUT96), .ZN(new_n478));
  XOR2_X1   g277(.A(G15gat), .B(G22gat), .Z(new_n479));
  INV_X1    g278(.A(G1gat), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT95), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n480), .A2(KEYINPUT94), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT16), .B1(new_n484), .B2(G1gat), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G8gat), .ZN(new_n488));
  INV_X1    g287(.A(G8gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n481), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n492));
  INV_X1    g291(.A(G50gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(G43gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(G43gat), .ZN(new_n495));
  INV_X1    g294(.A(G43gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(KEYINPUT93), .A3(G50gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT15), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n496), .A2(G50gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n501), .A3(KEYINPUT15), .ZN(new_n502));
  NAND2_X1  g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n504));
  INV_X1    g303(.A(G36gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n500), .A2(new_n502), .A3(new_n503), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(KEYINPUT92), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT92), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n511), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n512), .A3(new_n506), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n503), .ZN(new_n514));
  INV_X1    g313(.A(new_n502), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n491), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n488), .A2(new_n516), .A3(new_n509), .A4(new_n490), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n521), .B(KEYINPUT13), .Z(new_n522));
  AOI21_X1  g321(.A(new_n478), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n522), .ZN(new_n524));
  AOI211_X1 g323(.A(KEYINPUT96), .B(new_n524), .C1(new_n518), .C2(new_n519), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n517), .A2(KEYINPUT17), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n516), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n491), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n521), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n488), .A2(new_n490), .B1(new_n509), .B2(new_n516), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  OAI22_X1  g331(.A1(new_n523), .A2(new_n525), .B1(new_n532), .B2(KEYINPUT18), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(KEYINPUT18), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n477), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n522), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT96), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n478), .A3(new_n522), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n526), .A2(new_n528), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n521), .B(new_n518), .C1(new_n542), .C2(new_n491), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n477), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n540), .A2(new_n545), .A3(new_n546), .A4(new_n534), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n536), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n471), .A2(new_n472), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT104), .ZN(new_n550));
  OR2_X1    g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(KEYINPUT102), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT7), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT7), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(G85gat), .A3(G92gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G85gat), .ZN(new_n559));
  INV_X1    g358(.A(G92gat), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT8), .A2(new_n552), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n553), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT102), .ZN(new_n563));
  INV_X1    g362(.A(new_n552), .ZN(new_n564));
  NOR2_X1   g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n566), .A2(new_n553), .A3(new_n558), .A4(new_n561), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT103), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n550), .B1(new_n572), .B2(new_n541), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n541), .A3(new_n550), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT41), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n517), .B2(new_n570), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G190gat), .B(G218gat), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n576), .A2(new_n584), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n577), .A2(new_n578), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(KEYINPUT101), .Z(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n584), .B1(new_n576), .B2(new_n580), .ZN(new_n592));
  INV_X1    g391(.A(new_n580), .ZN(new_n593));
  AOI211_X1 g392(.A(new_n582), .B(new_n593), .C1(new_n574), .C2(new_n575), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G57gat), .ZN(new_n597));
  INV_X1    g396(.A(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G57gat), .A2(G64gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(KEYINPUT9), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  OR2_X1    g401(.A1(G71gat), .A2(G78gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT97), .ZN(new_n605));
  AND2_X1   g404(.A1(G57gat), .A2(G64gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(G57gat), .A2(G64gat), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n599), .A2(KEYINPUT97), .A3(new_n600), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(new_n602), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT9), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n602), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n602), .B2(new_n613), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n604), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G127gat), .B(G155gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n488), .B(new_n490), .C1(new_n618), .C2(new_n617), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT99), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G183gat), .B(G211gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT100), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n623), .B(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n596), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n612), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n634), .A2(new_n610), .A3(new_n609), .A4(new_n608), .ZN(new_n635));
  AOI221_X4 g434(.A(KEYINPUT102), .B1(new_n552), .B2(new_n551), .C1(new_n558), .C2(new_n561), .ZN(new_n636));
  AND4_X1   g435(.A1(new_n566), .A2(new_n553), .A3(new_n558), .A4(new_n561), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n604), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n617), .A2(new_n568), .A3(new_n569), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(KEYINPUT105), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n617), .A2(new_n643), .A3(new_n568), .A4(new_n569), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n640), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n638), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n640), .A2(new_n644), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n651), .B2(new_n649), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n641), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT10), .B1(new_n640), .B2(new_n644), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n655), .A2(KEYINPUT106), .A3(new_n650), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n645), .B(new_n648), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n645), .B1(new_n652), .B2(new_n642), .ZN(new_n658));
  INV_X1    g457(.A(new_n648), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n632), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n549), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n399), .A2(KEYINPUT84), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(new_n457), .A3(new_n400), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(new_n480), .ZN(G1324gat));
  NAND3_X1  g468(.A1(new_n549), .A2(new_n360), .A3(new_n664), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT16), .B(G8gat), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n549), .A2(KEYINPUT107), .A3(new_n360), .A4(new_n664), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR4_X1   g474(.A1(new_n670), .A2(KEYINPUT107), .A3(KEYINPUT42), .A4(new_n671), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT108), .B1(new_n670), .B2(G8gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n670), .A2(KEYINPUT108), .A3(G8gat), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n675), .A2(new_n676), .B1(new_n677), .B2(new_n679), .ZN(G1325gat));
  OAI21_X1  g479(.A(G15gat), .B1(new_n665), .B2(new_n453), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n460), .A2(new_n447), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n436), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n665), .B2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n665), .A2(new_n392), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n685), .B(new_n686), .Z(G1327gat));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  INV_X1    g487(.A(new_n468), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n667), .A2(new_n464), .ZN(new_n690));
  INV_X1    g489(.A(new_n392), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(KEYINPUT110), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n458), .B2(new_n392), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n424), .A2(new_n453), .A3(new_n692), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT111), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n452), .B1(new_n393), .B2(new_n423), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT111), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n697), .A2(new_n698), .A3(new_n694), .A4(new_n692), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n689), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n596), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n688), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n471), .A2(KEYINPUT44), .A3(new_n472), .A4(new_n596), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n662), .A2(new_n631), .ZN(new_n705));
  INV_X1    g504(.A(new_n548), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n667), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n701), .A2(new_n705), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT109), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n549), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n667), .A2(G29gat), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n710), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n549), .A2(KEYINPUT45), .A3(new_n712), .A4(new_n714), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n709), .A2(new_n716), .A3(new_n717), .ZN(G1328gat));
  OAI21_X1  g517(.A(G36gat), .B1(new_n708), .B2(new_n464), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n464), .A2(G36gat), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT46), .B1(new_n713), .B2(new_n721), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n713), .A2(KEYINPUT46), .A3(new_n721), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n719), .A2(new_n722), .A3(new_n723), .ZN(G1329gat));
  NOR2_X1   g523(.A1(new_n453), .A2(new_n496), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n704), .A2(new_n707), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n682), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n496), .B1(new_n713), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT47), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n726), .A2(new_n731), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1330gat));
  NAND4_X1  g532(.A1(new_n702), .A2(new_n691), .A3(new_n703), .A4(new_n707), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G50gat), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n691), .A2(new_n493), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n713), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n735), .B(KEYINPUT48), .C1(new_n713), .C2(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(G1331gat));
  INV_X1    g540(.A(new_n699), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT110), .B1(new_n690), .B2(new_n691), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n693), .B(new_n392), .C1(new_n667), .C2(new_n464), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n698), .B1(new_n745), .B2(new_n697), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n468), .B1(new_n742), .B2(new_n746), .ZN(new_n747));
  NOR4_X1   g546(.A1(new_n596), .A2(new_n662), .A3(new_n548), .A4(new_n631), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n667), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n597), .ZN(G1332gat));
  NOR2_X1   g550(.A1(new_n749), .A2(new_n464), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n756));
  INV_X1    g555(.A(new_n752), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT49), .B(G64gat), .Z(new_n758));
  OAI211_X1 g557(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT112), .B1(new_n760), .B2(new_n754), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1333gat));
  OR3_X1    g561(.A1(new_n749), .A2(G71gat), .A3(new_n727), .ZN(new_n763));
  OAI21_X1  g562(.A(G71gat), .B1(new_n749), .B2(new_n453), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1334gat));
  NOR2_X1   g566(.A1(new_n749), .A2(new_n392), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(G78gat), .Z(G1335gat));
  INV_X1    g568(.A(new_n631), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n662), .A2(new_n548), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n704), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n667), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n548), .A2(new_n770), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n747), .A2(new_n596), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n747), .A2(KEYINPUT51), .A3(new_n596), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n667), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n779), .A2(new_n559), .A3(new_n780), .A4(new_n661), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n773), .A2(new_n781), .ZN(G1336gat));
  NOR3_X1   g581(.A1(new_n464), .A2(new_n662), .A3(G92gat), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n702), .A2(new_n360), .A3(new_n703), .A4(new_n771), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n779), .A2(new_n783), .B1(G92gat), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n784), .A2(G92gat), .ZN(new_n788));
  INV_X1    g587(.A(new_n783), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n777), .B2(new_n778), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT52), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(G1337gat));
  OAI21_X1  g591(.A(G99gat), .B1(new_n772), .B2(new_n453), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n727), .A2(G99gat), .A3(new_n662), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1338gat));
  NOR3_X1   g595(.A1(new_n392), .A2(G106gat), .A3(new_n662), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT53), .B1(new_n779), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n702), .A2(new_n691), .A3(new_n703), .A4(new_n771), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT114), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n799), .A2(KEYINPUT114), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n799), .A2(G106gat), .ZN(new_n804));
  INV_X1    g603(.A(new_n797), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n805), .B1(new_n777), .B2(new_n778), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n803), .A2(new_n807), .ZN(G1339gat));
  NOR2_X1   g607(.A1(new_n529), .A2(new_n531), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n521), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n520), .A2(new_n522), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n476), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n547), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n661), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n652), .B2(new_n642), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n654), .B2(new_n656), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n815), .B(new_n641), .C1(new_n655), .C2(new_n650), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n818), .A2(new_n819), .A3(new_n659), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n818), .B2(new_n659), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n817), .B(KEYINPUT55), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n548), .A3(new_n657), .ZN(new_n823));
  INV_X1    g622(.A(new_n821), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n818), .A2(new_n819), .A3(new_n659), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT55), .B1(new_n826), .B2(new_n817), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n814), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n701), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n590), .A3(new_n595), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n827), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n822), .A2(new_n657), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n770), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n632), .A2(new_n706), .A3(new_n662), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT116), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n828), .A2(new_n701), .B1(new_n831), .B2(new_n833), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n839), .B(new_n836), .C1(new_n840), .C2(new_n770), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(new_n780), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n464), .A3(new_n461), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n706), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(new_n216), .ZN(G1340gat));
  NOR2_X1   g645(.A1(new_n844), .A2(new_n662), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(new_n213), .ZN(G1341gat));
  NOR2_X1   g647(.A1(new_n844), .A2(new_n631), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(new_n207), .ZN(G1342gat));
  NOR2_X1   g649(.A1(new_n844), .A2(new_n701), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n225), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n205), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(KEYINPUT56), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(KEYINPUT56), .B2(new_n853), .ZN(G1343gat));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n453), .A2(new_n691), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n360), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n706), .A2(G141gat), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n856), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n843), .A2(KEYINPUT121), .A3(new_n858), .A4(new_n860), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n453), .A2(new_n780), .A3(new_n464), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n838), .A2(new_n691), .A3(new_n841), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n871), .B1(new_n826), .B2(new_n817), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n814), .B1(new_n823), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n701), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n770), .B1(new_n874), .B2(new_n834), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT57), .B(new_n691), .C1(new_n875), .C2(new_n837), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT118), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n820), .A2(new_n821), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n651), .A2(new_n649), .ZN(new_n879));
  INV_X1    g678(.A(new_n650), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n642), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT54), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n880), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n642), .B1(new_n883), .B2(KEYINPUT106), .ZN(new_n884));
  INV_X1    g683(.A(new_n656), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n870), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n887), .A2(new_n548), .A3(new_n657), .A4(new_n822), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n596), .B1(new_n888), .B2(new_n814), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n830), .A2(new_n832), .A3(new_n827), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n631), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n392), .B1(new_n891), .B2(new_n836), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT57), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n866), .B1(new_n869), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G141gat), .B1(new_n896), .B2(new_n706), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT58), .B1(new_n864), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n877), .A2(new_n894), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n867), .A2(new_n868), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT119), .B(new_n865), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n877), .A3(new_n894), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n866), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G141gat), .B1(new_n906), .B2(new_n706), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT120), .B1(new_n859), .B2(new_n861), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT58), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n859), .A2(KEYINPUT120), .A3(new_n861), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n898), .B1(new_n907), .B2(new_n911), .ZN(G1344gat));
  NOR3_X1   g711(.A1(new_n859), .A2(G148gat), .A3(new_n662), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n239), .A2(KEYINPUT59), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n916), .B1(new_n905), .B2(new_n661), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n838), .A2(KEYINPUT57), .A3(new_n691), .A4(new_n841), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n661), .B(new_n866), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n918), .B1(new_n924), .B2(G148gat), .ZN(new_n925));
  OAI211_X1 g724(.A(KEYINPUT123), .B(new_n914), .C1(new_n917), .C2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n896), .A2(KEYINPUT119), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n903), .A2(new_n902), .A3(new_n866), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n661), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n925), .B1(new_n930), .B2(new_n915), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n927), .B1(new_n931), .B2(new_n913), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n926), .A2(new_n932), .ZN(G1345gat));
  NOR3_X1   g732(.A1(new_n906), .A2(new_n233), .A3(new_n631), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n859), .A2(new_n631), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n935), .A2(KEYINPUT124), .ZN(new_n936));
  AOI21_X1  g735(.A(G155gat), .B1(new_n935), .B2(KEYINPUT124), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1346gat));
  INV_X1    g737(.A(new_n859), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n268), .B1(new_n939), .B2(new_n596), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n701), .A2(new_n232), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n905), .B2(new_n941), .ZN(G1347gat));
  AND2_X1   g741(.A1(new_n842), .A2(new_n667), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n360), .A3(new_n461), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n944), .A2(G169gat), .A3(new_n706), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT125), .Z(new_n946));
  NOR2_X1   g745(.A1(new_n780), .A2(new_n464), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n682), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n392), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n950), .B1(new_n949), .B2(new_n948), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(new_n842), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G169gat), .B1(new_n953), .B2(new_n706), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n946), .A2(new_n954), .ZN(G1348gat));
  OAI21_X1  g754(.A(G176gat), .B1(new_n953), .B2(new_n662), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n661), .A2(new_n287), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n944), .B2(new_n957), .ZN(G1349gat));
  NOR3_X1   g757(.A1(new_n944), .A2(new_n299), .A3(new_n631), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n294), .B1(new_n952), .B2(new_n770), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n961), .B(new_n962), .ZN(G1350gat));
  AOI21_X1  g762(.A(new_n295), .B1(new_n952), .B2(new_n596), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT61), .Z(new_n965));
  NAND2_X1  g764(.A1(new_n596), .A2(new_n295), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n944), .B2(new_n966), .ZN(G1351gat));
  NOR2_X1   g766(.A1(new_n857), .A2(new_n464), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n943), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(G197gat), .B1(new_n970), .B2(new_n548), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n922), .A2(new_n923), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n453), .A2(new_n947), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n548), .A2(G197gat), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(G1352gat));
  NOR3_X1   g775(.A1(new_n969), .A2(G204gat), .A3(new_n662), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT62), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n972), .A2(new_n662), .A3(new_n973), .ZN(new_n979));
  INV_X1    g778(.A(G204gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(G1353gat));
  NAND3_X1  g780(.A1(new_n970), .A2(new_n334), .A3(new_n770), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n974), .A2(new_n770), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n335), .A3(new_n596), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n972), .A2(new_n701), .A3(new_n973), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n988), .B2(new_n335), .ZN(G1355gat));
endmodule


