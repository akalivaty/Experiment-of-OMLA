//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005;
  INV_X1    g000(.A(G1gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  INV_X1    g002(.A(G15gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G15gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(G1gat), .B1(new_n205), .B2(new_n207), .ZN(new_n210));
  OAI21_X1  g009(.A(G8gat), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n205), .A2(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(new_n202), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  INV_X1    g016(.A(G36gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT14), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT14), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G50gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G43gat), .ZN(new_n225));
  INV_X1    g024(.A(G43gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G50gat), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n223), .A2(KEYINPUT15), .A3(new_n225), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n227), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT15), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n225), .A2(new_n227), .A3(KEYINPUT15), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n222), .A2(KEYINPUT81), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(G29gat), .A3(G36gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n219), .A2(new_n234), .A3(new_n221), .A4(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n228), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n216), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n216), .A2(new_n238), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT83), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT83), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n216), .A2(new_n238), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n239), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT85), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n246), .B(KEYINPUT13), .Z(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OR3_X1    g047(.A1(new_n244), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n216), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT82), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n238), .A2(new_n251), .A3(KEYINPUT17), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT17), .B1(new_n238), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n241), .A2(new_n243), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT18), .A4(new_n246), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n245), .B1(new_n244), .B2(new_n248), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n249), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n254), .A2(new_n255), .A3(new_n246), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G141gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(G197gat), .ZN(new_n263));
  XOR2_X1   g062(.A(KEYINPUT11), .B(G169gat), .Z(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT12), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n258), .B(new_n261), .C1(KEYINPUT84), .C2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n249), .A2(new_n261), .A3(new_n256), .A4(new_n257), .ZN(new_n268));
  INV_X1    g067(.A(new_n266), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n249), .A2(new_n256), .A3(new_n257), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT84), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n268), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT34), .ZN(new_n275));
  INV_X1    g074(.A(G183gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT27), .B1(new_n276), .B2(KEYINPUT65), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT27), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(G183gat), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n277), .A2(new_n280), .A3(KEYINPUT66), .A4(new_n281), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT27), .B(G183gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n285), .A2(G190gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n279), .A2(G183gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n276), .A2(KEYINPUT27), .ZN(new_n293));
  AND4_X1   g092(.A1(new_n288), .A2(new_n290), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G169gat), .ZN(new_n297));
  INV_X1    g096(.A(G176gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT26), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT26), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n296), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n308), .A2(new_n309), .B1(G169gat), .B2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(new_n297), .A3(new_n298), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n276), .A2(new_n281), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(KEYINPUT24), .A3(new_n303), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n310), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n310), .A2(new_n314), .A3(new_n316), .A4(new_n318), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G134gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G127gat), .ZN(new_n326));
  INV_X1    g125(.A(G127gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G134gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(G113gat), .B2(G120gat), .ZN(new_n331));
  INV_X1    g130(.A(G113gat), .ZN(new_n332));
  INV_X1    g131(.A(G120gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n329), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n338));
  OAI21_X1  g137(.A(G120gat), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT1), .B1(new_n332), .B2(new_n333), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n326), .A3(new_n328), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n335), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n307), .A2(new_n324), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n329), .A2(new_n331), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n341), .B1(new_n332), .B2(new_n333), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n345), .A2(new_n339), .B1(new_n346), .B2(new_n329), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n305), .B1(new_n287), .B2(new_n295), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n320), .A2(new_n321), .B1(KEYINPUT64), .B2(KEYINPUT25), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G227gat), .ZN(new_n352));
  INV_X1    g151(.A(G233gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n275), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  AOI211_X1 g155(.A(KEYINPUT34), .B(new_n354), .C1(new_n344), .C2(new_n350), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(G15gat), .B(G43gat), .Z(new_n359));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n350), .A3(new_n354), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT33), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n363), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT32), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n365), .B1(new_n356), .B2(new_n357), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n367), .B2(new_n371), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT36), .ZN(new_n376));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(G197gat), .ZN(new_n378));
  INV_X1    g177(.A(G204gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G197gat), .A2(G204gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382));
  NAND2_X1  g181(.A1(G211gat), .A2(G218gat), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G211gat), .ZN(new_n385));
  INV_X1    g184(.A(G218gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT69), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n383), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n384), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G155gat), .ZN(new_n391));
  INV_X1    g190(.A(G162gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT71), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT71), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(G155gat), .B2(G162gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G148gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G141gat), .ZN(new_n399));
  INV_X1    g198(.A(G141gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(G148gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT2), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n391), .A3(new_n392), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n396), .ZN(new_n407));
  AND2_X1   g206(.A1(KEYINPUT72), .A2(G141gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(KEYINPUT72), .A2(G141gat), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n408), .A2(new_n409), .A3(new_n398), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n400), .A2(G148gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n405), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n390), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n387), .A2(new_n383), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n415), .B1(new_n384), .B2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n384), .A2(new_n419), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n413), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n412), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(new_n416), .B2(new_n417), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n377), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n416), .A2(KEYINPUT78), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n384), .A2(new_n389), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n384), .A2(new_n389), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n413), .B1(new_n430), .B2(KEYINPUT29), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n377), .B1(new_n431), .B2(new_n423), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n416), .A2(KEYINPUT78), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT79), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT31), .B(G50gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n206), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT79), .B1(new_n426), .B2(new_n434), .ZN(new_n442));
  INV_X1    g241(.A(new_n440), .ZN(new_n443));
  OAI21_X1  g242(.A(G22gat), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n435), .A2(new_n436), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n441), .A2(new_n446), .A3(new_n444), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT4), .B1(new_n423), .B2(new_n343), .ZN(new_n451));
  OR2_X1    g250(.A1(KEYINPUT72), .A2(G141gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(KEYINPUT72), .A2(G141gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(G148gat), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n399), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n455), .A2(new_n407), .B1(new_n397), .B2(new_n404), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n347), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n451), .A2(KEYINPUT75), .A3(new_n458), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n423), .A2(new_n343), .A3(KEYINPUT4), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT75), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT2), .B1(new_n399), .B2(new_n401), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n454), .A2(new_n399), .B1(new_n396), .B2(new_n406), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT3), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(new_n414), .A3(new_n343), .ZN(new_n468));
  NAND2_X1  g267(.A1(G225gat), .A2(G233gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(KEYINPUT5), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n459), .A2(new_n462), .A3(new_n468), .A4(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT76), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT74), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT73), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n457), .B1(new_n456), .B2(new_n347), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n468), .A2(new_n469), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n451), .A2(new_n458), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n480), .A2(KEYINPUT73), .A3(new_n469), .A4(new_n468), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n423), .A2(new_n343), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n345), .A2(new_n339), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n412), .A2(new_n405), .B1(new_n484), .B2(new_n335), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n470), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT5), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n474), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  AOI211_X1 g288(.A(KEYINPUT74), .B(new_n487), .C1(new_n479), .C2(new_n481), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n473), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G1gat), .B(G29gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT0), .ZN(new_n493));
  XNOR2_X1  g292(.A(G57gat), .B(G85gat), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n493), .B(new_n494), .Z(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n495), .B(new_n473), .C1(new_n489), .C2(new_n490), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n491), .A2(KEYINPUT6), .A3(new_n496), .ZN(new_n501));
  AND2_X1   g300(.A1(G226gat), .A2(G233gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(KEYINPUT29), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT70), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n307), .A2(new_n324), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT70), .B1(new_n348), .B2(new_n349), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n348), .A2(new_n349), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n502), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n390), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(new_n507), .A3(new_n502), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n503), .B1(new_n348), .B2(new_n349), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n430), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n516), .A2(KEYINPUT37), .ZN(new_n517));
  XNOR2_X1  g316(.A(G8gat), .B(G36gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(G64gat), .B(G92gat), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n518), .B(new_n519), .Z(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n516), .B2(KEYINPUT37), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT38), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n512), .A2(new_n515), .A3(new_n520), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n505), .B1(new_n307), .B2(new_n324), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT70), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n503), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n430), .B1(new_n528), .B2(new_n510), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n513), .A2(new_n430), .A3(new_n514), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n521), .A2(KEYINPUT37), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n513), .A2(new_n390), .A3(new_n514), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n534), .A2(KEYINPUT37), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n430), .B1(new_n508), .B2(new_n511), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT38), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n525), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n500), .A2(new_n501), .A3(new_n523), .A4(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT80), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT39), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n462), .A2(new_n468), .ZN(new_n542));
  INV_X1    g341(.A(new_n459), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n541), .B(new_n470), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n542), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n469), .B1(new_n545), .B2(new_n459), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n483), .A2(new_n485), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT39), .B1(new_n547), .B2(new_n470), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n495), .B(new_n544), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT40), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n540), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n546), .A2(new_n548), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n544), .A2(new_n495), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT80), .A4(KEYINPUT40), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n491), .A2(new_n496), .B1(new_n550), .B2(new_n549), .ZN(new_n556));
  OR3_X1    g355(.A1(new_n516), .A2(KEYINPUT30), .A3(new_n521), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n531), .A2(KEYINPUT30), .A3(new_n524), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n450), .B1(new_n539), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n558), .ZN(new_n561));
  INV_X1    g360(.A(new_n449), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n446), .B1(new_n441), .B2(new_n444), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n564), .B1(new_n501), .B2(new_n500), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n376), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n375), .A2(new_n561), .A3(new_n449), .A4(new_n448), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n500), .A2(new_n501), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT35), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n374), .ZN(new_n570));
  AND4_X1   g369(.A1(new_n372), .A2(new_n448), .A3(new_n570), .A4(new_n449), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT35), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n500), .A2(new_n501), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n561), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n274), .B1(new_n566), .B2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G134gat), .B(G162gat), .Z(new_n577));
  AND2_X1   g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n577), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT90), .B(KEYINPUT91), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(KEYINPUT92), .A3(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g384(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(G85gat), .A3(G92gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  AOI22_X1  g390(.A1(KEYINPUT8), .A2(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT93), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n595), .A3(new_n589), .ZN(new_n596));
  AND2_X1   g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT93), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n588), .A2(new_n599), .A3(new_n596), .A4(new_n592), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n603), .A2(new_n238), .B1(KEYINPUT41), .B2(new_n578), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT95), .Z(new_n605));
  XOR2_X1   g404(.A(G190gat), .B(G218gat), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n603), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT94), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(KEYINPUT94), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n609), .B(new_n610), .C1(new_n253), .C2(new_n252), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n607), .B1(new_n605), .B2(new_n611), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n583), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(new_n582), .A3(new_n612), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT9), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(G57gat), .A2(G64gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(G57gat), .A2(G64gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(G71gat), .A2(G78gat), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT86), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n626), .A3(new_n619), .ZN(new_n627));
  AND2_X1   g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT86), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n624), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  AND2_X1   g431(.A1(G57gat), .A2(G64gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(G57gat), .A2(G64gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n632), .A2(new_n635), .A3(new_n626), .A4(new_n621), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(KEYINPUT21), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n216), .B1(KEYINPUT21), .B2(new_n637), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT87), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT88), .ZN(new_n645));
  XNOR2_X1  g444(.A(G127gat), .B(G155gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT89), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n645), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G183gat), .B(G211gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n642), .B(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n618), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n596), .A2(new_n599), .A3(KEYINPUT96), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n603), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n637), .A2(new_n601), .A3(new_n602), .A4(new_n654), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT10), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n637), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n653), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n653), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n662), .A3(new_n657), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(G120gat), .B(G148gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT97), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n664), .A2(new_n668), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n652), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n576), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n573), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT98), .B(G1gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1324gat));
  INV_X1    g477(.A(new_n675), .ZN(new_n679));
  INV_X1    g478(.A(new_n561), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n679), .A2(KEYINPUT99), .A3(new_n680), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(G8gat), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT16), .B(G8gat), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n681), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n683), .B2(new_n684), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n685), .B(new_n688), .C1(new_n689), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g489(.A(G15gat), .B1(new_n675), .B2(new_n376), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n375), .A2(new_n204), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n675), .B2(new_n692), .ZN(G1326gat));
  INV_X1    g492(.A(new_n450), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n675), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT43), .B(G22gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n651), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n670), .A2(new_n671), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n615), .A2(new_n617), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n576), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n573), .A2(G29gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n709), .A2(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(KEYINPUT102), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n566), .A2(new_n575), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n618), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n704), .B1(new_n566), .B2(new_n575), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT44), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n703), .A2(new_n274), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n573), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n710), .A2(KEYINPUT45), .A3(new_n711), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n714), .A2(new_n724), .A3(new_n725), .ZN(G1328gat));
  OAI21_X1  g525(.A(G36gat), .B1(new_n723), .B2(new_n561), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n706), .A2(G36gat), .A3(new_n561), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT46), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1329gat));
  INV_X1    g529(.A(new_n376), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n722), .A2(G43gat), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n375), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n226), .B1(new_n706), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT47), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n732), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1330gat));
  AOI21_X1  g538(.A(new_n224), .B1(new_n722), .B2(new_n450), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n706), .A2(G50gat), .A3(new_n694), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(KEYINPUT103), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(KEYINPUT48), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n740), .B2(new_n741), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1331gat));
  AND4_X1   g547(.A1(new_n274), .A2(new_n715), .A3(new_n652), .A4(new_n701), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n568), .B(KEYINPUT104), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT105), .B(G57gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1332gat));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n680), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT49), .B(G64gat), .Z(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n754), .B2(new_n756), .ZN(G1333gat));
  NAND2_X1  g556(.A1(new_n749), .A2(new_n731), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n733), .A2(G71gat), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n758), .A2(G71gat), .B1(new_n749), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n749), .A2(new_n450), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n273), .A2(new_n700), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n701), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT106), .Z(new_n766));
  NAND3_X1  g565(.A1(new_n718), .A2(new_n720), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n590), .B1(new_n768), .B2(new_n568), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n719), .A2(new_n764), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT51), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n719), .A2(new_n774), .A3(new_n764), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n573), .A2(G85gat), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n773), .A2(new_n701), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n770), .A2(new_n771), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n777), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT107), .B1(new_n769), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1336gat));
  NAND4_X1  g580(.A1(new_n718), .A2(new_n680), .A3(new_n720), .A4(new_n766), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G92gat), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n773), .A2(new_n775), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n561), .A2(G92gat), .A3(new_n672), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT108), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n719), .A2(new_n764), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n719), .B2(new_n764), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n783), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n789), .B1(new_n794), .B2(KEYINPUT52), .ZN(new_n795));
  AOI211_X1 g594(.A(KEYINPUT109), .B(new_n784), .C1(new_n783), .C2(new_n793), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n788), .B1(new_n795), .B2(new_n796), .ZN(G1337gat));
  OR4_X1    g596(.A1(G99gat), .A2(new_n785), .A3(new_n733), .A4(new_n672), .ZN(new_n798));
  OAI21_X1  g597(.A(G99gat), .B1(new_n767), .B2(new_n376), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1338gat));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n768), .A2(new_n450), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n791), .A2(new_n792), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n694), .A2(G106gat), .A3(new_n672), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n802), .A2(G106gat), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n802), .A2(G106gat), .ZN(new_n806));
  INV_X1    g605(.A(new_n804), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n801), .B1(new_n785), .B2(new_n807), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n801), .A2(new_n805), .B1(new_n806), .B2(new_n808), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n674), .A2(new_n274), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n668), .B1(new_n661), .B2(KEYINPUT54), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT10), .ZN(new_n816));
  AND4_X1   g615(.A1(new_n637), .A2(new_n601), .A3(new_n602), .A4(new_n654), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n637), .A2(new_n654), .B1(new_n601), .B2(new_n602), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n659), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n815), .B1(new_n820), .B2(new_n653), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n662), .A3(new_n659), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n814), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n661), .A2(new_n822), .A3(new_n814), .A4(KEYINPUT54), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(KEYINPUT55), .B(new_n813), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n670), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n661), .A2(new_n822), .A3(KEYINPUT54), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT110), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n812), .B1(new_n829), .B2(new_n824), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(KEYINPUT55), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT111), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n669), .B1(new_n830), .B2(KEYINPUT55), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n813), .B1(new_n823), .B2(new_n825), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n832), .A2(new_n273), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n246), .B1(new_n254), .B2(new_n255), .ZN(new_n841));
  AOI211_X1 g640(.A(new_n247), .B(new_n239), .C1(new_n241), .C2(new_n243), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n265), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT112), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n845), .B(new_n265), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n844), .B(new_n846), .C1(new_n268), .C2(new_n269), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n840), .B1(new_n847), .B2(new_n672), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n258), .A2(new_n266), .A3(new_n261), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n844), .A2(new_n846), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n849), .A2(new_n850), .A3(KEYINPUT113), .A4(new_n701), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n618), .B1(new_n839), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n704), .A2(new_n847), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n832), .A2(new_n838), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n811), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n651), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n853), .A2(new_n811), .A3(new_n856), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n810), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(new_n750), .ZN(new_n861));
  INV_X1    g660(.A(new_n567), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n274), .A2(new_n338), .A3(new_n337), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n860), .A2(new_n571), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n573), .A2(new_n680), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n273), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n868), .A2(new_n869), .A3(G113gat), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n868), .B2(G113gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(G1340gat));
  NAND2_X1  g671(.A1(new_n701), .A2(new_n333), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT117), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n863), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n866), .A2(new_n701), .A3(new_n867), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(G120gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n876), .B2(G120gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(G1341gat));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n327), .A3(new_n700), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n866), .A2(new_n700), .A3(new_n867), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n327), .B2(new_n882), .ZN(G1342gat));
  NAND4_X1  g682(.A1(new_n860), .A2(new_n571), .A3(new_n618), .A4(new_n867), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G134gat), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n704), .A2(G134gat), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n860), .A2(new_n862), .A3(new_n750), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT56), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT119), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n889), .A2(KEYINPUT56), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n887), .A2(new_n891), .A3(new_n892), .ZN(G1343gat));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n731), .A2(new_n564), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n861), .A2(new_n400), .A3(new_n273), .A4(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n376), .A2(new_n867), .ZN(new_n897));
  OR2_X1    g696(.A1(KEYINPUT120), .A2(KEYINPUT55), .ZN(new_n898));
  NAND2_X1  g697(.A1(KEYINPUT120), .A2(KEYINPUT55), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n834), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n273), .A2(new_n833), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n850), .A2(new_n849), .A3(new_n701), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n618), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n651), .B1(new_n856), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n694), .B1(new_n904), .B2(new_n810), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT57), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n897), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n839), .A2(new_n852), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT114), .B(new_n855), .C1(new_n908), .C2(new_n618), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n651), .A3(new_n857), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n694), .B1(new_n910), .B2(new_n810), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n907), .B1(new_n911), .B2(new_n906), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n912), .A2(new_n273), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n452), .A2(new_n453), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n894), .B(new_n896), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n896), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n912), .B2(new_n273), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT58), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(G1344gat));
  AND2_X1   g719(.A1(new_n861), .A2(new_n895), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n398), .A3(new_n701), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n860), .A2(new_n450), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT57), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n618), .A2(new_n833), .A3(new_n836), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n847), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n928), .B1(new_n927), .B2(new_n926), .ZN(new_n929));
  INV_X1    g728(.A(new_n903), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n810), .B1(new_n931), .B2(new_n700), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n906), .A3(new_n450), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n672), .B1(new_n897), .B2(KEYINPUT121), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n925), .A2(new_n933), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n923), .B1(new_n936), .B2(G148gat), .ZN(new_n937));
  AOI211_X1 g736(.A(KEYINPUT59), .B(new_n398), .C1(new_n912), .C2(new_n701), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n922), .B1(new_n937), .B2(new_n938), .ZN(G1345gat));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n391), .A3(new_n700), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n912), .A2(new_n700), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n391), .ZN(G1346gat));
  AOI21_X1  g741(.A(G162gat), .B1(new_n921), .B2(new_n618), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n704), .A2(new_n392), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n912), .B2(new_n944), .ZN(G1347gat));
  AOI21_X1  g744(.A(new_n568), .B1(new_n910), .B2(new_n810), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n733), .A2(new_n450), .A3(new_n561), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n297), .A3(new_n273), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n750), .A2(new_n561), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n860), .A2(new_n273), .A3(new_n571), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G169gat), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n950), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n951), .B1(new_n950), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(G1348gat));
  AND3_X1   g756(.A1(new_n860), .A2(new_n571), .A3(new_n952), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n298), .B1(new_n958), .B2(new_n701), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n948), .A2(G176gat), .A3(new_n672), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n959), .A2(new_n960), .ZN(G1349gat));
  AOI21_X1  g760(.A(new_n276), .B1(new_n958), .B2(new_n700), .ZN(new_n962));
  AND4_X1   g761(.A1(new_n289), .A2(new_n946), .A3(new_n700), .A4(new_n947), .ZN(new_n963));
  OR3_X1    g762(.A1(new_n962), .A2(KEYINPUT60), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT60), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n281), .A3(new_n618), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n860), .A2(new_n571), .A3(new_n618), .A4(new_n952), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n968), .A2(new_n969), .A3(G190gat), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n968), .B2(G190gat), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n971), .A2(new_n972), .A3(KEYINPUT61), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n968), .A2(G190gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n974), .B1(new_n976), .B2(new_n970), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n967), .B1(new_n973), .B2(new_n977), .ZN(G1351gat));
  NOR3_X1   g777(.A1(new_n731), .A2(new_n561), .A3(new_n694), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n946), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n378), .A3(new_n273), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n750), .A2(new_n731), .A3(new_n561), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n933), .B(new_n982), .C1(new_n911), .C2(new_n906), .ZN(new_n983));
  OAI21_X1  g782(.A(KEYINPUT125), .B1(new_n983), .B2(new_n274), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G197gat), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n983), .A2(KEYINPUT125), .A3(new_n274), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(G1352gat));
  NAND3_X1  g786(.A1(new_n980), .A2(new_n379), .A3(new_n701), .ZN(new_n988));
  XOR2_X1   g787(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n988), .A2(new_n990), .ZN(new_n992));
  OAI21_X1  g791(.A(G204gat), .B1(new_n983), .B2(new_n672), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(G1353gat));
  NAND3_X1  g793(.A1(new_n980), .A2(new_n385), .A3(new_n700), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT63), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n996), .A2(KEYINPUT127), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n925), .A2(new_n700), .A3(new_n933), .A4(new_n982), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n385), .B1(KEYINPUT127), .B2(new_n996), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI211_X1 g799(.A(new_n999), .B(new_n997), .C1(new_n983), .C2(new_n651), .ZN(new_n1001));
  INV_X1    g800(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n995), .B1(new_n1000), .B2(new_n1002), .ZN(G1354gat));
  OAI21_X1  g802(.A(G218gat), .B1(new_n983), .B2(new_n704), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n980), .A2(new_n386), .A3(new_n618), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(G1355gat));
endmodule


