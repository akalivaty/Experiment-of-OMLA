//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n637,
    new_n638, new_n641, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(G137), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n471), .B1(new_n463), .B2(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT66), .B1(new_n472), .B2(new_n464), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G125), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n470), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n473), .B2(new_n479), .ZN(G160));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n474), .A2(new_n475), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT67), .ZN(new_n487));
  OR2_X1    g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n464), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT68), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n484), .B2(new_n464), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AOI211_X1 g069(.A(new_n483), .B(new_n487), .C1(G124), .C2(new_n494), .ZN(G162));
  NAND3_X1  g070(.A1(new_n490), .A2(KEYINPUT69), .A3(G126), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n464), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT70), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n500), .ZN(new_n503));
  INV_X1    g078(.A(new_n501), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n496), .A2(new_n499), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n464), .A2(G138), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n508), .B1(new_n488), .B2(new_n489), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n511));
  NOR3_X1   g086(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G138), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(G2105), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n514), .B1(new_n474), .B2(new_n475), .ZN(new_n515));
  AOI21_X1  g090(.A(KEYINPUT71), .B1(new_n515), .B2(KEYINPUT4), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n514), .B(new_n511), .C1(new_n475), .C2(new_n474), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT72), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n463), .A2(new_n520), .A3(new_n511), .A4(new_n514), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n507), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(G164));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G50), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n526), .A2(new_n527), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G62), .ZN(new_n539));
  NAND2_X1  g114(.A1(G75), .A2(G543), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT73), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n535), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n534), .A2(new_n542), .ZN(G303));
  INV_X1    g118(.A(G303), .ZN(G166));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  INV_X1    g121(.A(G51), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n526), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n529), .A2(new_n528), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n525), .A2(G89), .ZN(new_n550));
  NAND2_X1  g125(.A1(G63), .A2(G651), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n548), .A2(new_n552), .ZN(G168));
  AOI22_X1  g128(.A1(new_n538), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n535), .ZN(new_n555));
  INV_X1    g130(.A(G52), .ZN(new_n556));
  INV_X1    g131(.A(G90), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n526), .A2(new_n556), .B1(new_n532), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(G171));
  AOI22_X1  g134(.A1(new_n538), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n535), .ZN(new_n561));
  INV_X1    g136(.A(G43), .ZN(new_n562));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n526), .A2(new_n562), .B1(new_n532), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT74), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n538), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n549), .A2(KEYINPUT77), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G65), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  INV_X1    g154(.A(new_n532), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G91), .ZN(new_n581));
  INV_X1    g156(.A(G53), .ZN(new_n582));
  NAND2_X1  g157(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n526), .A2(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n530), .A2(new_n531), .ZN(new_n587));
  INV_X1    g162(.A(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n589), .A2(G53), .A3(new_n583), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n586), .B2(new_n590), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n579), .B(new_n581), .C1(new_n592), .C2(new_n594), .ZN(G299));
  INV_X1    g170(.A(G171), .ZN(G301));
  INV_X1    g171(.A(G168), .ZN(G286));
  INV_X1    g172(.A(G49), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n526), .A2(KEYINPUT78), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT78), .B1(new_n526), .B2(new_n598), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G74), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n535), .B1(new_n549), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(G87), .B2(new_n580), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(G288));
  NAND3_X1  g180(.A1(new_n538), .A2(new_n525), .A3(G86), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n525), .A2(G48), .A3(G543), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(KEYINPUT79), .A2(G73), .A3(G543), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(KEYINPUT79), .B1(G73), .B2(G543), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(G61), .B1(new_n529), .B2(new_n528), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n535), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(G305));
  AOI22_X1  g191(.A1(new_n580), .A2(G85), .B1(new_n589), .B2(G47), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n538), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n535), .B2(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT80), .B(G66), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n573), .B2(new_n574), .ZN(new_n622));
  AND2_X1   g197(.A1(G79), .A2(G543), .ZN(new_n623));
  OR3_X1    g198(.A1(new_n622), .A2(KEYINPUT81), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT81), .B1(new_n622), .B2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(G651), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n580), .A2(KEYINPUT10), .A3(G92), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  INV_X1    g203(.A(G92), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n532), .B2(new_n629), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n627), .A2(new_n630), .B1(G54), .B2(new_n589), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n620), .B1(new_n633), .B2(G868), .ZN(G284));
  OAI21_X1  g209(.A(new_n620), .B1(new_n633), .B2(G868), .ZN(G321));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NOR2_X1   g211(.A1(G286), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G299), .B(KEYINPUT82), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n636), .ZN(G280));
  XOR2_X1   g214(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n633), .B1(new_n641), .B2(G860), .ZN(G148));
  NAND2_X1  g217(.A1(new_n633), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G868), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g221(.A1(new_n463), .A2(new_n464), .ZN(new_n647));
  INV_X1    g222(.A(G135), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n464), .A2(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  OAI22_X1  g225(.A1(new_n647), .A2(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n494), .B2(G123), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n463), .A2(new_n467), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT12), .Z(new_n657));
  XOR2_X1   g232(.A(KEYINPUT13), .B(G2100), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n659), .ZN(G156));
  XOR2_X1   g235(.A(KEYINPUT15), .B(G2435), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT85), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(KEYINPUT14), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2451), .B(G2454), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1341), .B(G1348), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT86), .Z(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n676), .A2(G14), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G401));
  XOR2_X1   g254(.A(G2067), .B(G2678), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT87), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT88), .Z(new_n682));
  NOR2_X1   g257(.A1(G2072), .A2(G2078), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n442), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT17), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G2084), .B(G2090), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(KEYINPUT89), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n686), .B(new_n687), .C1(new_n682), .C2(new_n688), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT18), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n682), .A2(new_n687), .A3(new_n685), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2096), .B(G2100), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G227));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1971), .B(G1976), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT19), .ZN(new_n699));
  XOR2_X1   g274(.A(G1956), .B(G2474), .Z(new_n700));
  XOR2_X1   g275(.A(G1961), .B(G1966), .Z(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT20), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n700), .A2(new_n701), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n699), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n699), .B2(new_n705), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT90), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(G1991), .B(G1996), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n711), .A2(new_n712), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n697), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n711), .A2(new_n712), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n717), .A2(new_n696), .A3(new_n713), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(G229));
  MUX2_X1   g295(.A(G24), .B(G290), .S(G16), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT94), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G1986), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n485), .A2(G131), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT92), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n494), .A2(G119), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n464), .A2(G107), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G25), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT91), .Z(new_n736));
  AOI21_X1  g311(.A(new_n724), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT96), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n723), .B(new_n737), .C1(new_n738), .C2(KEYINPUT36), .ZN(new_n739));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G23), .ZN(new_n741));
  INV_X1    g316(.A(G288), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n740), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT33), .B(G1976), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n740), .A2(G22), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G166), .B2(new_n740), .ZN(new_n747));
  INV_X1    g322(.A(G1971), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G6), .A2(G16), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n615), .B2(G16), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT32), .B(G1981), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n745), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT95), .B(KEYINPUT34), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n733), .A2(new_n724), .A3(new_n736), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n739), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n738), .A2(KEYINPUT36), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n734), .A2(G33), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT102), .B(KEYINPUT25), .Z(new_n763));
  NAND3_X1  g338(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G139), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(new_n647), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(new_n464), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n762), .B1(new_n770), .B2(new_n734), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT103), .Z(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G2072), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT104), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(KEYINPUT104), .ZN(new_n775));
  NOR2_X1   g350(.A1(G171), .A2(new_n740), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G5), .B2(new_n740), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  NOR2_X1   g353(.A1(G16), .A2(G19), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n565), .B2(G16), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT98), .B(G1341), .Z(new_n781));
  AOI22_X1  g356(.A1(new_n777), .A2(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n772), .B2(G2072), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n774), .A2(new_n775), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n740), .A2(G20), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT23), .ZN(new_n787));
  INV_X1    g362(.A(G299), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n740), .ZN(new_n789));
  INV_X1    g364(.A(G1956), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT24), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G34), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n734), .B1(new_n792), .B2(G34), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT105), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G160), .B2(G29), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(G2084), .ZN(new_n799));
  NOR2_X1   g374(.A1(G27), .A2(G29), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G164), .B2(G29), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G2078), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n801), .A2(G2078), .B1(G2084), .B2(new_n798), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n791), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n740), .A2(G4), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n633), .B2(new_n740), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT97), .B(G1348), .Z(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n785), .A2(new_n806), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n734), .A2(G35), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT108), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G162), .B2(new_n734), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT29), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2090), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT30), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n818), .A2(G28), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n734), .B1(new_n818), .B2(G28), .ZN(new_n820));
  AND2_X1   g395(.A1(KEYINPUT31), .A2(G11), .ZN(new_n821));
  NOR2_X1   g396(.A1(KEYINPUT31), .A2(G11), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n819), .A2(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n740), .A2(G21), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G168), .B2(new_n740), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n823), .B1(new_n825), .B2(G1966), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n826), .B1(new_n654), .B2(new_n734), .C1(new_n778), .C2(new_n777), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(G1966), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT106), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT107), .Z(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT100), .B(KEYINPUT28), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT101), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n734), .A2(G26), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n833), .B(new_n834), .Z(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n836));
  INV_X1    g411(.A(G116), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(G2105), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n485), .B2(G140), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n491), .A2(new_n493), .ZN(new_n840));
  INV_X1    g415(.A(G128), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT99), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n844), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n835), .B1(new_n846), .B2(G29), .ZN(new_n847));
  INV_X1    g422(.A(G2067), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n734), .A2(G32), .ZN(new_n850));
  NAND3_X1  g425(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT26), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n467), .A2(G105), .ZN(new_n853));
  INV_X1    g428(.A(G141), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n852), .B(new_n853), .C1(new_n647), .C2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G129), .B2(new_n494), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n850), .B1(new_n856), .B2(new_n734), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT27), .ZN(new_n858));
  INV_X1    g433(.A(G1996), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NOR4_X1   g435(.A1(new_n817), .A2(new_n831), .A3(new_n849), .A4(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n760), .A2(new_n761), .A3(new_n812), .A4(new_n861), .ZN(G150));
  INV_X1    g437(.A(G150), .ZN(G311));
  NOR2_X1   g438(.A1(new_n632), .A2(new_n641), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT38), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n538), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(new_n535), .ZN(new_n867));
  INV_X1    g442(.A(G55), .ZN(new_n868));
  INV_X1    g443(.A(G93), .ZN(new_n869));
  OAI22_X1  g444(.A1(new_n526), .A2(new_n868), .B1(new_n532), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n565), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n865), .B(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  INV_X1    g449(.A(G860), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n871), .A2(new_n875), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(G145));
  XNOR2_X1  g455(.A(new_n654), .B(KEYINPUT109), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G160), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n882), .A2(G162), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(G162), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n846), .B(new_n856), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n523), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n769), .B2(new_n767), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n485), .A2(G142), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n464), .A2(G118), .ZN(new_n890));
  OAI21_X1  g465(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(G130), .B2(new_n494), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(new_n657), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n731), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n886), .B(G164), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n770), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n888), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n885), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n888), .A2(new_n897), .ZN(new_n900));
  INV_X1    g475(.A(new_n895), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n904), .A3(new_n898), .ZN(new_n905));
  INV_X1    g480(.A(new_n885), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n888), .A2(KEYINPUT110), .A3(new_n897), .A4(new_n895), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n903), .A2(new_n908), .A3(KEYINPUT40), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT40), .B1(new_n903), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(G395));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n632), .A2(G559), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n872), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n632), .A2(G299), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n592), .A2(new_n594), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n578), .A2(G651), .B1(G91), .B2(new_n580), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n916), .A2(new_n626), .A3(new_n917), .A4(new_n631), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(KEYINPUT41), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n915), .A2(new_n918), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(KEYINPUT111), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT111), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n919), .A2(new_n927), .A3(KEYINPUT41), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n643), .B(new_n872), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n912), .B(new_n922), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n926), .B2(new_n928), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT42), .B1(new_n932), .B2(new_n921), .ZN(new_n933));
  XOR2_X1   g508(.A(G290), .B(G303), .Z(new_n934));
  XNOR2_X1  g509(.A(G288), .B(new_n615), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n934), .B(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n931), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n931), .B2(new_n933), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n636), .B1(new_n867), .B2(new_n870), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(G295));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n940), .A2(new_n943), .A3(new_n941), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(new_n940), .B2(new_n941), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(G331));
  XNOR2_X1  g521(.A(G171), .B(G168), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n872), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT113), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n872), .B2(new_n947), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n928), .A3(new_n926), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n872), .A2(new_n947), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n919), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n948), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n937), .ZN(new_n956));
  INV_X1    g531(.A(G37), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n951), .A2(new_n936), .A3(new_n954), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n920), .A2(KEYINPUT114), .A3(new_n924), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT115), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n923), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n925), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n919), .A2(KEYINPUT115), .A3(KEYINPUT41), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n961), .A2(new_n963), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n948), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n952), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n949), .A2(new_n953), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n936), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n958), .A2(new_n957), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n960), .B1(new_n973), .B2(KEYINPUT43), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n959), .A2(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n971), .A2(new_n972), .A3(new_n977), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT44), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n976), .A2(new_n980), .ZN(G397));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n510), .B1(new_n509), .B2(new_n511), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n515), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n983), .A2(new_n984), .B1(new_n519), .B2(new_n521), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n506), .A2(new_n502), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT69), .B1(new_n490), .B2(G126), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n497), .A2(new_n498), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n982), .B1(new_n985), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n469), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n464), .B1(new_n476), .B2(new_n470), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(new_n478), .ZN(new_n995));
  AOI211_X1 g570(.A(KEYINPUT66), .B(new_n464), .C1(new_n476), .C2(new_n470), .ZN(new_n996));
  OAI211_X1 g571(.A(G40), .B(new_n993), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n731), .B(new_n724), .Z(new_n999));
  XNOR2_X1  g574(.A(new_n846), .B(new_n848), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n856), .B(G1996), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(KEYINPUT116), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G290), .A2(G1986), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1006), .B(new_n1007), .Z(new_n1008));
  OAI21_X1  g583(.A(new_n998), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1966), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n523), .B2(new_n982), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n991), .A2(G1384), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n985), .B2(new_n989), .ZN(new_n1013));
  INV_X1    g588(.A(G40), .ZN(new_n1014));
  AOI211_X1 g589(.A(new_n1014), .B(new_n469), .C1(new_n473), .C2(new_n479), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT121), .B(new_n1010), .C1(new_n1011), .C2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n997), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n1018));
  INV_X1    g593(.A(G2084), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(new_n982), .C1(new_n985), .C2(new_n989), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n997), .B1(new_n523), .B2(new_n1012), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n992), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT121), .B1(new_n1025), .B2(new_n1010), .ZN(new_n1026));
  OAI21_X1  g601(.A(G8), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT124), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT117), .B(G8), .Z(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G286), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n1031), .B(KEYINPUT123), .Z(new_n1032));
  INV_X1    g607(.A(KEYINPUT124), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1033), .B(G8), .C1(new_n1023), .C2(new_n1026), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1028), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT51), .B1(new_n1036), .B2(new_n1032), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1036), .A2(new_n1029), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1032), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(KEYINPUT62), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT62), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1032), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1027), .B2(KEYINPUT124), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1037), .B1(new_n1048), .B2(new_n1034), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1046), .B1(new_n1049), .B2(new_n1043), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  XOR2_X1   g626(.A(new_n1051), .B(KEYINPUT55), .Z(new_n1052));
  INV_X1    g627(.A(G2090), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n1054));
  AND4_X1   g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1015), .A4(new_n1021), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1971), .B1(new_n1024), .B2(new_n992), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1052), .B(G8), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(G1981), .B1(new_n608), .B2(new_n614), .ZN(new_n1058));
  INV_X1    g633(.A(G61), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n536), .B2(new_n537), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G73), .A2(G543), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT79), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n609), .ZN(new_n1064));
  OAI21_X1  g639(.A(G651), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1981), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n606), .A4(new_n607), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT49), .B1(new_n1058), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1058), .A2(KEYINPUT49), .A3(new_n1067), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1030), .B1(new_n990), .B2(new_n997), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT119), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n519), .A2(new_n521), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n516), .B2(new_n512), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1384), .B1(new_n1075), .B2(new_n507), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1029), .B1(new_n1076), .B2(new_n1015), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1058), .A2(KEYINPUT49), .A3(new_n1067), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(new_n1068), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n601), .A2(G1976), .A3(new_n604), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(new_n1030), .C1(new_n990), .C2(new_n997), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1073), .A2(new_n1081), .B1(KEYINPUT52), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  INV_X1    g660(.A(G1976), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1088), .B2(new_n1083), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1077), .A2(KEYINPUT118), .A3(new_n1082), .A4(new_n1087), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1057), .A2(new_n1084), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1025), .A2(new_n748), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1018), .A2(new_n1053), .A3(new_n1021), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1029), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1095), .A2(new_n1052), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n992), .A2(new_n803), .A3(new_n1015), .A4(new_n1013), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1054), .A2(new_n1015), .A3(new_n1021), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n778), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1024), .A2(new_n992), .A3(KEYINPUT53), .A4(new_n803), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AND4_X1   g678(.A1(G171), .A2(new_n1092), .A3(new_n1096), .A4(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1045), .A2(new_n1050), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1043), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1100), .A2(new_n790), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT57), .B1(new_n586), .B2(new_n590), .ZN(new_n1109));
  AOI22_X1  g684(.A1(G299), .A2(KEYINPUT57), .B1(new_n917), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1024), .A2(new_n992), .A3(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1107), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1076), .A2(new_n1116), .A3(new_n1015), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT122), .B1(new_n990), .B2(new_n997), .ZN(new_n1118));
  AOI21_X1  g693(.A(G2067), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n810), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1122), .A3(KEYINPUT60), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1125), .A3(new_n633), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n917), .A2(new_n1109), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n788), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1112), .ZN(new_n1130));
  AOI21_X1  g705(.A(G1956), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(KEYINPUT61), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1115), .A2(new_n1126), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT58), .B(G1341), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1136), .A2(new_n1137), .B1(new_n1025), .B2(G1996), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n565), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1120), .A2(new_n1122), .A3(KEYINPUT60), .A4(new_n632), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(KEYINPUT59), .A3(new_n565), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1114), .B1(new_n1145), .B2(new_n633), .ZN(new_n1146));
  OAI22_X1  g721(.A1(new_n1135), .A2(new_n1144), .B1(new_n1146), .B2(new_n1113), .ZN(new_n1147));
  XNOR2_X1  g722(.A(G171), .B(KEYINPUT54), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1013), .A2(KEYINPUT53), .A3(new_n803), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n465), .A2(G40), .A3(new_n468), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  OR3_X1    g728(.A1(new_n1152), .A2(new_n1153), .A3(new_n994), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(new_n1152), .B2(new_n994), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1151), .B1(new_n1011), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n992), .A2(KEYINPUT126), .A3(new_n1155), .A4(new_n1154), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1150), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1148), .B1(new_n1149), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1148), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1163), .A2(new_n1092), .A3(new_n1096), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1106), .A2(new_n1147), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT63), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1095), .B2(new_n1052), .ZN(new_n1168));
  OAI211_X1 g743(.A(G168), .B(new_n1030), .C1(new_n1023), .C2(new_n1026), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1057), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n742), .A2(new_n1086), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1073), .B2(new_n1081), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1067), .ZN(new_n1175));
  OR3_X1    g750(.A1(new_n1174), .A2(KEYINPUT120), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT120), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1176), .A2(new_n1077), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(G8), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1084), .B(new_n1091), .C1(new_n1180), .C2(new_n1052), .ZN(new_n1181));
  OAI21_X1  g756(.A(KEYINPUT63), .B1(new_n1181), .B2(new_n1169), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1172), .A2(new_n1178), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1166), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1009), .B1(new_n1105), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1004), .A2(new_n998), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n998), .A2(new_n1005), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT48), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n998), .A2(new_n859), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT46), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1000), .A2(new_n856), .ZN(new_n1194));
  INV_X1    g769(.A(new_n998), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT47), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1003), .A2(new_n724), .A3(new_n731), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(G2067), .B2(new_n846), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n998), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1191), .A2(new_n1197), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1186), .A2(new_n1187), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1009), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1049), .A2(new_n1164), .A3(new_n1043), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1183), .B1(new_n1205), .B2(new_n1147), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1045), .A2(new_n1050), .A3(new_n1104), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1204), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(KEYINPUT127), .B1(new_n1208), .B2(new_n1201), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1203), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g785(.A1(G227), .A2(new_n461), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1212), .B1(new_n675), .B2(new_n677), .ZN(new_n1213));
  AND2_X1   g787(.A1(new_n719), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n903), .A2(new_n908), .ZN(new_n1215));
  NAND3_X1  g789(.A1(new_n1214), .A2(new_n974), .A3(new_n1215), .ZN(G225));
  INV_X1    g790(.A(G225), .ZN(G308));
endmodule


