//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT81), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n204), .B1(G155gat), .B2(G162gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n207), .A2(G148gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT80), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT79), .B(G148gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n210), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT80), .A3(G141gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n203), .A2(new_n206), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n207), .A2(G148gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n206), .B1(new_n208), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n202), .A2(KEYINPUT78), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n202), .A2(KEYINPUT78), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT83), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT4), .ZN(new_n226));
  INV_X1    g025(.A(new_n223), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(new_n216), .B2(new_n217), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G113gat), .B(G120gat), .Z(new_n231));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(G127gat), .A2(G134gat), .ZN(new_n234));
  INV_X1    g033(.A(G134gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT67), .B(G127gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n233), .B(new_n234), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n231), .A2(new_n232), .A3(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n230), .A4(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n241), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT4), .B1(new_n224), .B2(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT5), .ZN(new_n247));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n244), .B1(new_n228), .B2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n247), .B(new_n248), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G1gat), .B(G29gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT0), .ZN(new_n255));
  XNOR2_X1  g054(.A(G57gat), .B(G85gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  OAI21_X1  g056(.A(new_n226), .B1(new_n224), .B2(new_n244), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n258), .B(new_n248), .C1(new_n249), .C2(new_n251), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n225), .A2(KEYINPUT4), .A3(new_n242), .A4(new_n230), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n248), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n224), .A2(new_n244), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n242), .A2(new_n228), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n253), .B(new_n257), .C1(new_n262), .C2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n257), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n260), .B2(new_n261), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n246), .A2(new_n252), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(KEYINPUT6), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n277));
  XOR2_X1   g076(.A(G197gat), .B(G204gat), .Z(new_n278));
  NAND2_X1  g077(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT22), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n280), .A2(new_n281), .B1(G211gat), .B2(G218gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n278), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n283), .A2(KEYINPUT74), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n284), .B1(new_n283), .B2(KEYINPUT74), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(G183gat), .B2(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n294), .A2(KEYINPUT65), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT24), .B1(new_n294), .B2(KEYINPUT65), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT23), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  INV_X1    g100(.A(G169gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n299), .B(new_n301), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n297), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT64), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n293), .B1(new_n308), .B2(new_n294), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n305), .B1(new_n309), .B2(new_n304), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n306), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n310), .A2(new_n307), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT27), .B(G183gat), .ZN(new_n313));
  INV_X1    g112(.A(G190gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(KEYINPUT28), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n313), .A2(KEYINPUT66), .ZN(new_n316));
  INV_X1    g115(.A(G183gat), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT66), .B1(new_n317), .B2(KEYINPUT27), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n314), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n315), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n321));
  INV_X1    g120(.A(new_n294), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n302), .A2(new_n303), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n323), .A2(KEYINPUT26), .A3(new_n298), .ZN(new_n324));
  AOI211_X1 g123(.A(new_n322), .B(new_n324), .C1(KEYINPUT26), .C2(new_n298), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n311), .A2(new_n312), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G226gat), .ZN(new_n328));
  INV_X1    g127(.A(G233gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(KEYINPUT29), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n326), .B(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n330), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n291), .B(new_n332), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n327), .A2(new_n335), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n334), .B2(new_n331), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n338), .B2(new_n291), .ZN(new_n339));
  XOR2_X1   g138(.A(G8gat), .B(G36gat), .Z(new_n340));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n342), .B(KEYINPUT77), .Z(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n336), .B(new_n342), .C1(new_n338), .C2(new_n291), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n277), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n277), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n276), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT69), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n242), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n244), .A2(KEYINPUT69), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n327), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n326), .A2(new_n244), .A3(KEYINPUT69), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n354), .A2(G227gat), .A3(G233gat), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT32), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT33), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G15gat), .B(G43gat), .Z(new_n360));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n362), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n356), .B(KEYINPUT32), .C1(new_n358), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT71), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n354), .A2(new_n355), .B1(G227gat), .B2(G233gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(KEYINPUT70), .A2(KEYINPUT34), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(G22gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT29), .B1(new_n228), .B2(new_n250), .ZN(new_n379));
  INV_X1    g178(.A(new_n291), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT84), .ZN(new_n382));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(new_n379), .B2(new_n380), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n283), .A2(new_n284), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n287), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n250), .B1(new_n387), .B2(KEYINPUT29), .ZN(new_n388));
  INV_X1    g187(.A(new_n230), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n228), .A2(new_n229), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n382), .A2(new_n383), .A3(new_n385), .A4(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n250), .B1(new_n291), .B2(KEYINPUT29), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n393), .A2(new_n224), .ZN(new_n394));
  OAI211_X1 g193(.A(G228gat), .B(G233gat), .C1(new_n394), .C2(new_n381), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT31), .B(G50gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n392), .B2(new_n395), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n378), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n377), .A3(new_n398), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n366), .A2(new_n367), .A3(new_n373), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n375), .A2(new_n401), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT35), .B1(new_n350), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT35), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n366), .A2(new_n374), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n373), .A2(new_n363), .A3(new_n365), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND4_X1   g209(.A1(new_n407), .A2(new_n410), .A3(new_n403), .A4(new_n401), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(new_n276), .A3(new_n349), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n401), .A2(new_n403), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n249), .A2(new_n251), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n263), .B1(new_n246), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT39), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n264), .A2(new_n265), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(new_n248), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n417), .B(new_n263), .C1(new_n246), .C2(new_n415), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n257), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT40), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n420), .A2(KEYINPUT40), .A3(new_n257), .A4(new_n421), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n272), .B1(new_n346), .B2(new_n348), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n414), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT38), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n342), .B1(new_n339), .B2(KEYINPUT37), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n336), .B(new_n431), .C1(new_n338), .C2(new_n291), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n429), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n380), .B(new_n332), .C1(new_n334), .C2(new_n335), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(KEYINPUT37), .C1(new_n338), .C2(new_n380), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(new_n432), .A3(new_n429), .A4(new_n343), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n436), .A2(new_n345), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n274), .A2(new_n275), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n438), .B2(KEYINPUT85), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n274), .A2(new_n440), .A3(new_n275), .A4(new_n437), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n428), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n414), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n350), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT72), .B1(new_n410), .B2(KEYINPUT36), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n375), .A2(KEYINPUT36), .A3(new_n404), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT72), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT36), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n408), .A2(new_n447), .A3(new_n448), .A4(new_n409), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n413), .B1(new_n442), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G43gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G50gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT15), .ZN(new_n455));
  INV_X1    g254(.A(G50gat), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(G43gat), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT87), .ZN(new_n458));
  AND2_X1   g257(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n458), .B(new_n456), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT15), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n453), .ZN(new_n464));
  NAND2_X1  g263(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n465));
  AOI21_X1  g264(.A(G50gat), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n454), .A2(KEYINPUT87), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n461), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT14), .B(G29gat), .ZN(new_n469));
  INV_X1    g268(.A(G36gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n472), .A2(new_n470), .A3(G29gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n457), .B1(new_n468), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n475), .A2(new_n457), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT17), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT17), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n457), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n473), .B1(new_n470), .B2(new_n469), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT15), .B1(new_n466), .B2(new_n458), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n459), .A2(new_n460), .ZN(new_n483));
  OAI211_X1 g282(.A(KEYINPUT87), .B(new_n454), .C1(new_n483), .C2(G50gat), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n481), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n479), .B(new_n480), .C1(new_n485), .C2(new_n457), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487));
  INV_X1    g286(.A(G1gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT16), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(G1gat), .B2(new_n487), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G8gat), .ZN(new_n492));
  INV_X1    g291(.A(G8gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n490), .B(new_n493), .C1(G1gat), .C2(new_n487), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n486), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n476), .A2(new_n477), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n495), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT18), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n497), .A2(KEYINPUT18), .A3(new_n498), .A4(new_n500), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n499), .B(new_n495), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n498), .B(KEYINPUT13), .Z(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(G197gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT11), .B(G169gat), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n510), .B(new_n511), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT12), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n501), .A2(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(new_n513), .A3(new_n504), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n452), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT101), .ZN(new_n520));
  XNOR2_X1  g319(.A(G183gat), .B(G211gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n521), .B(new_n522), .Z(new_n523));
  AND2_X1   g322(.A1(G71gat), .A2(G78gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(G71gat), .A2(G78gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT9), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT88), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n526), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n536));
  OR2_X1    g335(.A1(G57gat), .A2(G64gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(G57gat), .A2(G64gat), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n537), .B(new_n538), .C1(new_n524), .C2(new_n525), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n539), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n530), .A2(KEYINPUT89), .A3(new_n532), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n527), .A2(new_n531), .A3(new_n528), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n531), .B1(new_n527), .B2(new_n528), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n526), .A2(new_n534), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n546), .A2(new_n542), .A3(new_n547), .A4(new_n536), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n535), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT21), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n496), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT92), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n551), .ZN(new_n554));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G127gat), .B(G155gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT20), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n556), .A2(new_n558), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n553), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n553), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n556), .A2(new_n558), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n559), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n523), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n568));
  INV_X1    g367(.A(G99gat), .ZN(new_n569));
  INV_X1    g368(.A(G106gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT93), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(G85gat), .A3(G92gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT7), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n574), .A2(new_n577), .A3(G85gat), .A4(G92gat), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(KEYINPUT94), .A2(G92gat), .ZN(new_n580));
  INV_X1    g379(.A(G85gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(KEYINPUT94), .A2(G92gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n572), .A2(KEYINPUT8), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n568), .B(new_n573), .C1(new_n579), .C2(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n583), .A2(new_n584), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n573), .A2(new_n568), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n576), .A2(new_n578), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n571), .A2(KEYINPUT95), .A3(new_n572), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n586), .A2(new_n591), .A3(KEYINPUT96), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n594), .A2(new_n478), .A3(new_n486), .A4(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n586), .A2(new_n591), .A3(KEYINPUT96), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT96), .B1(new_n586), .B2(new_n591), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n499), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT41), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n596), .A2(new_n599), .A3(new_n605), .A4(new_n601), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n600), .A2(KEYINPUT41), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n604), .A2(KEYINPUT98), .A3(new_n606), .A4(new_n610), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n604), .A2(KEYINPUT97), .A3(new_n606), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n599), .A2(new_n601), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n605), .A4(new_n596), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n609), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n562), .A2(new_n565), .A3(new_n523), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n567), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G120gat), .B(G148gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT100), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n592), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n535), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n546), .A2(new_n542), .A3(new_n547), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT90), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n633), .B1(new_n635), .B2(new_n548), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n586), .A2(new_n591), .A3(KEYINPUT99), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n632), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n586), .A2(new_n591), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n636), .A2(new_n639), .A3(KEYINPUT99), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n630), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n597), .A2(new_n598), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(KEYINPUT10), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n629), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n638), .A2(new_n640), .A3(new_n628), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n627), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n550), .A2(new_n631), .A3(new_n592), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n636), .A3(new_n637), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT10), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n628), .B1(new_n651), .B2(new_n644), .ZN(new_n652));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  INV_X1    g452(.A(new_n627), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n520), .B1(new_n623), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n622), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n566), .ZN(new_n659));
  INV_X1    g458(.A(new_n656), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(KEYINPUT101), .A3(new_n621), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n519), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n276), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g465(.A(KEYINPUT16), .B(G8gat), .ZN(new_n667));
  INV_X1    g466(.A(new_n349), .ZN(new_n668));
  INV_X1    g467(.A(new_n662), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n452), .A2(new_n668), .A3(new_n518), .A4(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n667), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT103), .B1(new_n674), .B2(KEYINPUT42), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n670), .B(KEYINPUT102), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n676), .B(new_n677), .C1(new_n678), .C2(new_n667), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n670), .A2(new_n677), .A3(new_n667), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n678), .B2(G8gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n675), .A2(new_n679), .A3(new_n681), .ZN(G1325gat));
  AOI21_X1  g481(.A(G15gat), .B1(new_n663), .B2(new_n410), .ZN(new_n683));
  INV_X1    g482(.A(new_n450), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(G15gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT104), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n683), .B1(new_n663), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n663), .A2(new_n443), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NAND2_X1  g489(.A1(new_n567), .A2(new_n622), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n648), .ZN(new_n692));
  INV_X1    g491(.A(new_n655), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n613), .A2(new_n614), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n615), .A2(new_n619), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n452), .A2(new_n518), .A3(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n699), .A2(G29gat), .A3(new_n276), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT45), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n691), .B(KEYINPUT105), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n518), .A3(new_n660), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n452), .A2(new_n620), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n452), .B(new_n620), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n703), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n664), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G29gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n701), .A2(new_n713), .ZN(G1328gat));
  NOR3_X1   g513(.A1(new_n699), .A2(G36gat), .A3(new_n349), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n711), .A2(new_n668), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n470), .B2(new_n718), .ZN(G1329gat));
  NOR2_X1   g518(.A1(new_n450), .A2(new_n483), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n711), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n410), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n483), .B1(new_n699), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT47), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n721), .A2(new_n726), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1330gat));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n456), .B1(new_n711), .B2(new_n443), .ZN(new_n730));
  INV_X1    g529(.A(new_n699), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n443), .A2(new_n456), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT108), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n729), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n703), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n708), .A2(new_n709), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n704), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n705), .B1(new_n452), .B2(new_n620), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n443), .B(new_n737), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G50gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(KEYINPUT48), .A3(new_n734), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n743), .ZN(G1331gat));
  NOR3_X1   g543(.A1(new_n623), .A2(new_n518), .A3(new_n660), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n452), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n276), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT109), .B(G57gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1332gat));
  NOR2_X1   g548(.A1(new_n746), .A2(new_n349), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(G1333gat));
  INV_X1    g553(.A(new_n746), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(G71gat), .A3(new_n684), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n410), .B(KEYINPUT110), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n746), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(G71gat), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n755), .A2(new_n443), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n659), .A2(new_n518), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT111), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n656), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n707), .B2(new_n710), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(new_n664), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n452), .A2(new_n620), .A3(new_n765), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n452), .A2(KEYINPUT51), .A3(new_n620), .A4(new_n765), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n664), .A2(new_n581), .A3(new_n656), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT112), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n768), .A2(new_n581), .B1(new_n774), .B2(new_n776), .ZN(G1336gat));
  INV_X1    g576(.A(new_n580), .ZN(new_n778));
  INV_X1    g577(.A(new_n582), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n767), .B2(new_n668), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n349), .A2(G92gat), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n660), .B(new_n783), .C1(new_n771), .C2(new_n772), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n766), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n668), .B(new_n786), .C1(new_n739), .C2(new_n740), .ZN(new_n787));
  INV_X1    g586(.A(new_n780), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n656), .A3(new_n782), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n785), .A2(new_n792), .ZN(G1337gat));
  NAND4_X1  g592(.A1(new_n773), .A2(new_n569), .A3(new_n410), .A4(new_n656), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n767), .A2(new_n684), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n569), .ZN(G1338gat));
  AOI21_X1  g595(.A(new_n570), .B1(new_n767), .B2(new_n443), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n414), .A2(G106gat), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI211_X1 g598(.A(new_n660), .B(new_n799), .C1(new_n771), .C2(new_n772), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT53), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n443), .B(new_n786), .C1(new_n739), .C2(new_n740), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G106gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n773), .A2(new_n656), .A3(new_n798), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n806), .ZN(G1339gat));
  NOR3_X1   g606(.A1(new_n623), .A2(new_n518), .A3(new_n656), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n505), .A2(new_n506), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n498), .B1(new_n497), .B2(new_n500), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n512), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n517), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n641), .A2(new_n645), .A3(new_n629), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n815), .A2(new_n652), .A3(KEYINPUT54), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n817), .B(new_n628), .C1(new_n651), .C2(new_n644), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n627), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n814), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(new_n652), .A3(KEYINPUT54), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n627), .A4(new_n818), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n696), .A2(new_n813), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n812), .B1(new_n648), .B2(new_n655), .ZN(new_n824));
  AND4_X1   g623(.A1(new_n513), .A2(new_n503), .A3(new_n504), .A4(new_n507), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n513), .B1(new_n516), .B2(new_n504), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n655), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n646), .A2(new_n817), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n819), .B1(new_n828), .B2(new_n815), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n827), .B1(new_n829), .B2(KEYINPUT55), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n824), .B1(new_n830), .B2(new_n820), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n823), .B1(new_n831), .B2(new_n620), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n808), .B1(new_n702), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n443), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n276), .A2(new_n668), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n410), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(G113gat), .ZN(new_n837));
  INV_X1    g636(.A(new_n518), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n833), .A2(new_n276), .A3(new_n405), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n349), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n518), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n839), .B1(new_n837), .B2(new_n842), .ZN(G1340gat));
  INV_X1    g642(.A(G120gat), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n836), .A2(new_n844), .A3(new_n660), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n656), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n844), .B2(new_n846), .ZN(G1341gat));
  NOR3_X1   g646(.A1(new_n836), .A2(new_n236), .A3(new_n702), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n841), .A2(new_n659), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT113), .Z(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n850), .B2(new_n236), .ZN(G1342gat));
  NAND2_X1  g650(.A1(new_n349), .A2(new_n620), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT114), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n840), .A2(new_n854), .A3(new_n235), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n836), .B2(new_n621), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(G1343gat));
  NAND2_X1  g658(.A1(new_n450), .A2(new_n835), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n450), .A2(KEYINPUT115), .A3(new_n835), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n833), .B2(new_n414), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n832), .A2(new_n691), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT57), .B(new_n443), .C1(new_n867), .C2(new_n808), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n864), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G141gat), .B1(new_n870), .B2(new_n838), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n450), .A2(new_n443), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(new_n833), .A3(new_n276), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n873), .A2(new_n349), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n207), .A3(new_n518), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g676(.A1(new_n874), .A2(new_n212), .A3(new_n656), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n660), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n881), .B(new_n823), .C1(new_n831), .C2(new_n620), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n646), .A2(new_n647), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n883), .A2(new_n654), .B1(new_n515), .B2(new_n517), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n820), .A2(new_n822), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n824), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n620), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n620), .A2(new_n655), .A3(new_n813), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n820), .A2(new_n822), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT116), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n882), .A2(new_n891), .A3(new_n691), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n657), .A2(new_n838), .A3(new_n661), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n414), .B1(new_n894), .B2(KEYINPUT117), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT57), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n833), .A2(new_n865), .A3(new_n414), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n880), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n879), .B1(new_n900), .B2(G148gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n210), .A2(new_n879), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n869), .B2(new_n656), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n878), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT118), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n906), .B(new_n878), .C1(new_n901), .C2(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1345gat));
  OAI21_X1  g707(.A(G155gat), .B1(new_n870), .B2(new_n702), .ZN(new_n909));
  INV_X1    g708(.A(G155gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n874), .A2(new_n910), .A3(new_n659), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1346gat));
  OAI21_X1  g711(.A(G162gat), .B1(new_n870), .B2(new_n621), .ZN(new_n913));
  INV_X1    g712(.A(G162gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n873), .A2(new_n914), .A3(new_n854), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1347gat));
  NAND2_X1  g715(.A1(new_n276), .A2(new_n668), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n758), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n834), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n838), .ZN(new_n920));
  NOR4_X1   g719(.A1(new_n833), .A2(new_n664), .A3(new_n349), .A4(new_n405), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n302), .A3(new_n518), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT119), .Z(G1348gat));
  OAI21_X1  g723(.A(G176gat), .B1(new_n919), .B2(new_n660), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n303), .A3(new_n656), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1349gat));
  OAI21_X1  g726(.A(G183gat), .B1(new_n919), .B2(new_n702), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n921), .A2(new_n313), .A3(new_n659), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT60), .B1(new_n930), .B2(KEYINPUT120), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT120), .B1(new_n930), .B2(KEYINPUT121), .ZN(new_n932));
  MUX2_X1   g731(.A(KEYINPUT60), .B(new_n931), .S(new_n932), .Z(G1350gat));
  NAND3_X1  g732(.A1(new_n921), .A2(new_n314), .A3(new_n620), .ZN(new_n934));
  OAI21_X1  g733(.A(G190gat), .B1(new_n919), .B2(new_n621), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(KEYINPUT122), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(KEYINPUT122), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT61), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n872), .A2(new_n349), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n833), .A2(new_n664), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(KEYINPUT123), .B(G197gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n518), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n443), .A3(new_n897), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n899), .B1(new_n950), .B2(new_n865), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n951), .A2(KEYINPUT124), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(KEYINPUT124), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n684), .A2(new_n917), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n955), .A2(new_n838), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n948), .B1(new_n956), .B2(new_n947), .ZN(G1352gat));
  XNOR2_X1  g756(.A(KEYINPUT125), .B(G204gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n955), .B2(new_n660), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n945), .A2(new_n660), .A3(new_n958), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT62), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1353gat));
  OR3_X1    g761(.A1(new_n945), .A2(G211gat), .A3(new_n691), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n954), .A2(new_n659), .ZN(new_n964));
  OAI211_X1 g763(.A(KEYINPUT63), .B(G211gat), .C1(new_n951), .C2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n964), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n967), .B1(new_n898), .B2(new_n899), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n963), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g771(.A(KEYINPUT126), .B(new_n963), .C1(new_n966), .C2(new_n969), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1354gat));
  INV_X1    g773(.A(G218gat), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n955), .A2(new_n975), .A3(new_n621), .ZN(new_n976));
  AOI21_X1  g775(.A(G218gat), .B1(new_n946), .B2(new_n620), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT127), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n976), .A2(new_n978), .ZN(G1355gat));
endmodule


