

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  XNOR2_X2 U325 ( .A(n345), .B(n344), .ZN(n369) );
  XOR2_X2 U326 ( .A(G92GAT), .B(KEYINPUT73), .Z(n345) );
  XOR2_X1 U327 ( .A(KEYINPUT41), .B(n480), .Z(n555) );
  XNOR2_X1 U328 ( .A(n389), .B(n388), .ZN(n480) );
  XNOR2_X1 U329 ( .A(n379), .B(n378), .ZN(n381) );
  NOR2_X1 U330 ( .A1(n550), .A2(n555), .ZN(n390) );
  XNOR2_X1 U331 ( .A(n381), .B(n380), .ZN(n389) );
  XNOR2_X1 U332 ( .A(n347), .B(n346), .ZN(n348) );
  AND2_X1 U333 ( .A1(n416), .A2(n294), .ZN(n293) );
  XOR2_X1 U334 ( .A(KEYINPUT114), .B(n415), .Z(n294) );
  NOR2_X2 U335 ( .A1(n536), .A2(n458), .ZN(n568) );
  XOR2_X1 U336 ( .A(KEYINPUT36), .B(KEYINPUT104), .Z(n295) );
  XOR2_X1 U337 ( .A(n339), .B(n338), .Z(n296) );
  NOR2_X1 U338 ( .A1(n576), .A2(n414), .ZN(n415) );
  INV_X1 U339 ( .A(KEYINPUT32), .ZN(n376) );
  XNOR2_X1 U340 ( .A(n377), .B(n376), .ZN(n378) );
  INV_X1 U341 ( .A(n369), .ZN(n346) );
  XNOR2_X1 U342 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U343 ( .A(n567), .B(n295), .ZN(n588) );
  XNOR2_X1 U344 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U345 ( .A(KEYINPUT28), .B(n470), .Z(n534) );
  XNOR2_X1 U346 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U347 ( .A(n462), .B(n461), .ZN(G1349GAT) );
  XOR2_X1 U348 ( .A(G176GAT), .B(KEYINPUT85), .Z(n298) );
  XNOR2_X1 U349 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n309) );
  XOR2_X1 U351 ( .A(G99GAT), .B(G190GAT), .Z(n300) );
  XOR2_X1 U352 ( .A(G120GAT), .B(G71GAT), .Z(n383) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G127GAT), .Z(n403) );
  XNOR2_X1 U354 ( .A(n383), .B(n403), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U356 ( .A(n301), .B(G134GAT), .Z(n307) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n302), .B(KEYINPUT84), .ZN(n437) );
  XOR2_X1 U359 ( .A(G169GAT), .B(n437), .Z(n304) );
  NAND2_X1 U360 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U362 ( .A(G43GAT), .B(n305), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n314) );
  XOR2_X1 U365 ( .A(G183GAT), .B(KEYINPUT19), .Z(n311) );
  XNOR2_X1 U366 ( .A(KEYINPUT88), .B(KEYINPUT18), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n313) );
  XOR2_X1 U368 ( .A(KEYINPUT17), .B(KEYINPUT87), .Z(n312) );
  XOR2_X1 U369 ( .A(n313), .B(n312), .Z(n318) );
  XOR2_X2 U370 ( .A(n314), .B(n318), .Z(n536) );
  XOR2_X1 U371 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n316) );
  NAND2_X1 U372 ( .A1(G226GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U374 ( .A(n317), .B(G92GAT), .Z(n326) );
  INV_X1 U375 ( .A(n318), .ZN(n324) );
  XOR2_X1 U376 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n320) );
  XNOR2_X1 U377 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U379 ( .A(n321), .B(G211GAT), .Z(n323) );
  XNOR2_X1 U380 ( .A(G197GAT), .B(G204GAT), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n456) );
  XOR2_X1 U382 ( .A(n324), .B(n456), .Z(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U384 ( .A(G176GAT), .B(G64GAT), .Z(n380) );
  XOR2_X1 U385 ( .A(n327), .B(n380), .Z(n330) );
  XOR2_X1 U386 ( .A(G169GAT), .B(G8GAT), .Z(n354) );
  XNOR2_X1 U387 ( .A(G36GAT), .B(G190GAT), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n328), .B(KEYINPUT80), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n354), .B(n333), .ZN(n329) );
  XNOR2_X1 U390 ( .A(n330), .B(n329), .ZN(n524) );
  XOR2_X1 U391 ( .A(G29GAT), .B(G43GAT), .Z(n332) );
  XNOR2_X1 U392 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n355) );
  XNOR2_X1 U394 ( .A(n355), .B(n333), .ZN(n351) );
  XOR2_X1 U395 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n335) );
  XNOR2_X1 U396 ( .A(G218GAT), .B(KEYINPUT66), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U398 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n337) );
  XNOR2_X1 U399 ( .A(KEYINPUT68), .B(KEYINPUT65), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U401 ( .A(KEYINPUT11), .B(KEYINPUT78), .Z(n341) );
  NAND2_X1 U402 ( .A1(G232GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U404 ( .A(G106GAT), .B(n342), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n296), .B(n343), .ZN(n349) );
  XOR2_X1 U406 ( .A(G50GAT), .B(G162GAT), .Z(n450) );
  XOR2_X1 U407 ( .A(G134GAT), .B(KEYINPUT79), .Z(n429) );
  XNOR2_X1 U408 ( .A(n450), .B(n429), .ZN(n347) );
  XNOR2_X1 U409 ( .A(G99GAT), .B(G85GAT), .ZN(n344) );
  XOR2_X1 U410 ( .A(n351), .B(n350), .Z(n562) );
  INV_X1 U411 ( .A(n562), .ZN(n567) );
  XOR2_X1 U412 ( .A(G141GAT), .B(G197GAT), .Z(n353) );
  XNOR2_X1 U413 ( .A(G113GAT), .B(G15GAT), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n368) );
  XOR2_X1 U415 ( .A(n354), .B(G36GAT), .Z(n357) );
  XNOR2_X1 U416 ( .A(n355), .B(G50GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U418 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n359) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U421 ( .A(n361), .B(n360), .Z(n366) );
  XOR2_X1 U422 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n363) );
  XNOR2_X1 U423 ( .A(G22GAT), .B(G1GAT), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n364), .B(KEYINPUT29), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n576) );
  INV_X1 U428 ( .A(n576), .ZN(n550) );
  XNOR2_X1 U429 ( .A(n369), .B(KEYINPUT31), .ZN(n370) );
  AND2_X1 U430 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  NAND2_X1 U431 ( .A1(n370), .A2(n371), .ZN(n375) );
  INV_X1 U432 ( .A(n370), .ZN(n373) );
  INV_X1 U433 ( .A(n371), .ZN(n372) );
  NAND2_X1 U434 ( .A1(n373), .A2(n372), .ZN(n374) );
  NAND2_X1 U435 ( .A1(n375), .A2(n374), .ZN(n379) );
  XOR2_X1 U436 ( .A(G57GAT), .B(KEYINPUT13), .Z(n393) );
  XNOR2_X1 U437 ( .A(G204GAT), .B(n393), .ZN(n377) );
  XNOR2_X1 U438 ( .A(G106GAT), .B(G78GAT), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n382), .B(G148GAT), .ZN(n444) );
  XOR2_X1 U440 ( .A(n383), .B(n444), .Z(n387) );
  XOR2_X1 U441 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n385) );
  XNOR2_X1 U442 ( .A(KEYINPUT72), .B(KEYINPUT75), .ZN(n384) );
  XOR2_X1 U443 ( .A(n385), .B(n384), .Z(n386) );
  XNOR2_X1 U444 ( .A(n390), .B(KEYINPUT46), .ZN(n408) );
  XOR2_X1 U445 ( .A(G78GAT), .B(G211GAT), .Z(n392) );
  XNOR2_X1 U446 ( .A(G183GAT), .B(G71GAT), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n407) );
  XOR2_X1 U448 ( .A(G22GAT), .B(G155GAT), .Z(n451) );
  XOR2_X1 U449 ( .A(n393), .B(n451), .Z(n395) );
  NAND2_X1 U450 ( .A1(G231GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U452 ( .A(KEYINPUT82), .B(KEYINPUT12), .Z(n397) );
  XNOR2_X1 U453 ( .A(KEYINPUT81), .B(KEYINPUT15), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n405) );
  XOR2_X1 U456 ( .A(KEYINPUT14), .B(G64GAT), .Z(n401) );
  XNOR2_X1 U457 ( .A(G1GAT), .B(G8GAT), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U461 ( .A(n407), .B(n406), .Z(n558) );
  INV_X1 U462 ( .A(n558), .ZN(n584) );
  NOR2_X1 U463 ( .A1(n408), .A2(n584), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n409), .B(KEYINPUT113), .ZN(n410) );
  NOR2_X1 U465 ( .A1(n567), .A2(n410), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n411), .B(KEYINPUT47), .ZN(n416) );
  NOR2_X1 U467 ( .A1(n558), .A2(n588), .ZN(n412) );
  XNOR2_X1 U468 ( .A(KEYINPUT45), .B(n412), .ZN(n413) );
  NAND2_X1 U469 ( .A1(n413), .A2(n480), .ZN(n414) );
  XNOR2_X1 U470 ( .A(KEYINPUT48), .B(n293), .ZN(n532) );
  NOR2_X1 U471 ( .A1(n524), .A2(n532), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n417), .B(KEYINPUT54), .ZN(n440) );
  XOR2_X1 U473 ( .A(G57GAT), .B(G155GAT), .Z(n419) );
  XNOR2_X1 U474 ( .A(G127GAT), .B(G148GAT), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U476 ( .A(KEYINPUT93), .B(KEYINPUT95), .Z(n421) );
  XNOR2_X1 U477 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U479 ( .A(n423), .B(n422), .Z(n435) );
  XOR2_X1 U480 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n425) );
  XNOR2_X1 U481 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n433) );
  XOR2_X1 U483 ( .A(G85GAT), .B(G162GAT), .Z(n427) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(G120GAT), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U486 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U492 ( .A(G141GAT), .B(KEYINPUT3), .Z(n438) );
  XOR2_X1 U493 ( .A(KEYINPUT2), .B(n438), .Z(n449) );
  XOR2_X1 U494 ( .A(n439), .B(n449), .Z(n520) );
  NAND2_X1 U495 ( .A1(n440), .A2(n520), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n441), .B(KEYINPUT64), .ZN(n573) );
  XOR2_X1 U497 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n443) );
  XNOR2_X1 U498 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n448) );
  XOR2_X1 U500 ( .A(n444), .B(KEYINPUT92), .Z(n446) );
  NAND2_X1 U501 ( .A1(G228GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(n470) );
  NOR2_X1 U508 ( .A1(n573), .A2(n470), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n457), .B(KEYINPUT55), .ZN(n458) );
  INV_X1 U510 ( .A(n555), .ZN(n539) );
  NAND2_X1 U511 ( .A1(n568), .A2(n539), .ZN(n462) );
  XOR2_X1 U512 ( .A(G176GAT), .B(KEYINPUT56), .Z(n460) );
  XNOR2_X1 U513 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n459) );
  INV_X1 U514 ( .A(n520), .ZN(n472) );
  NOR2_X1 U515 ( .A1(n524), .A2(n536), .ZN(n463) );
  NOR2_X1 U516 ( .A1(n470), .A2(n463), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n464), .B(KEYINPUT25), .ZN(n467) );
  XOR2_X1 U518 ( .A(n524), .B(KEYINPUT27), .Z(n471) );
  NAND2_X1 U519 ( .A1(n470), .A2(n536), .ZN(n465) );
  XOR2_X1 U520 ( .A(n465), .B(KEYINPUT26), .Z(n571) );
  NAND2_X1 U521 ( .A1(n471), .A2(n571), .ZN(n466) );
  NAND2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U523 ( .A(KEYINPUT98), .B(n468), .Z(n469) );
  NOR2_X1 U524 ( .A1(n472), .A2(n469), .ZN(n475) );
  NAND2_X1 U525 ( .A1(n536), .A2(n534), .ZN(n473) );
  NAND2_X1 U526 ( .A1(n472), .A2(n471), .ZN(n531) );
  NOR2_X1 U527 ( .A1(n473), .A2(n531), .ZN(n474) );
  NOR2_X1 U528 ( .A1(n475), .A2(n474), .ZN(n493) );
  XOR2_X1 U529 ( .A(KEYINPUT16), .B(KEYINPUT83), .Z(n477) );
  NAND2_X1 U530 ( .A1(n584), .A2(n562), .ZN(n476) );
  XNOR2_X1 U531 ( .A(n477), .B(n476), .ZN(n478) );
  NOR2_X1 U532 ( .A1(n493), .A2(n478), .ZN(n479) );
  XOR2_X1 U533 ( .A(KEYINPUT99), .B(n479), .Z(n507) );
  INV_X1 U534 ( .A(n480), .ZN(n580) );
  NOR2_X1 U535 ( .A1(n580), .A2(n550), .ZN(n481) );
  XNOR2_X1 U536 ( .A(n481), .B(KEYINPUT76), .ZN(n497) );
  NAND2_X1 U537 ( .A1(n507), .A2(n497), .ZN(n490) );
  NOR2_X1 U538 ( .A1(n520), .A2(n490), .ZN(n483) );
  XNOR2_X1 U539 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U541 ( .A(G1GAT), .B(n484), .Z(G1324GAT) );
  NOR2_X1 U542 ( .A1(n524), .A2(n490), .ZN(n486) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1325GAT) );
  NOR2_X1 U545 ( .A1(n536), .A2(n490), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(n489), .ZN(G1326GAT) );
  NOR2_X1 U549 ( .A1(n534), .A2(n490), .ZN(n492) );
  XNOR2_X1 U550 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1327GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT105), .B(KEYINPUT37), .Z(n496) );
  NOR2_X1 U553 ( .A1(n493), .A2(n588), .ZN(n494) );
  NAND2_X1 U554 ( .A1(n494), .A2(n558), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n519) );
  NAND2_X1 U556 ( .A1(n497), .A2(n519), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n498), .B(KEYINPUT38), .ZN(n505) );
  NOR2_X1 U558 ( .A1(n505), .A2(n520), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n499), .B(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(n500), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n524), .A2(n505), .ZN(n501) );
  XOR2_X1 U562 ( .A(KEYINPUT106), .B(n501), .Z(n502) );
  XNOR2_X1 U563 ( .A(G36GAT), .B(n502), .ZN(G1329GAT) );
  NOR2_X1 U564 ( .A1(n505), .A2(n536), .ZN(n503) );
  XOR2_X1 U565 ( .A(KEYINPUT40), .B(n503), .Z(n504) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NOR2_X1 U567 ( .A1(n505), .A2(n534), .ZN(n506) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n506), .Z(G1331GAT) );
  XNOR2_X1 U569 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n511) );
  NOR2_X1 U570 ( .A1(n555), .A2(n576), .ZN(n518) );
  NAND2_X1 U571 ( .A1(n507), .A2(n518), .ZN(n515) );
  NOR2_X1 U572 ( .A1(n520), .A2(n515), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U576 ( .A1(n524), .A2(n515), .ZN(n512) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n536), .A2(n515), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n534), .A2(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n528) );
  NOR2_X1 U585 ( .A1(n520), .A2(n528), .ZN(n522) );
  XNOR2_X1 U586 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n528), .ZN(n525) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n536), .A2(n528), .ZN(n526) );
  XOR2_X1 U592 ( .A(KEYINPUT112), .B(n526), .Z(n527) );
  XNOR2_X1 U593 ( .A(G99GAT), .B(n527), .ZN(G1338GAT) );
  NOR2_X1 U594 ( .A1(n534), .A2(n528), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(n529), .Z(n530) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n538) );
  NOR2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U599 ( .A(n533), .B(KEYINPUT115), .Z(n549) );
  NAND2_X1 U600 ( .A1(n549), .A2(n534), .ZN(n535) );
  NOR2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n546), .A2(n576), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U605 ( .A1(n546), .A2(n539), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U607 ( .A(G120GAT), .B(n542), .Z(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n544) );
  NAND2_X1 U609 ( .A1(n546), .A2(n584), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n545), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n567), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n549), .A2(n571), .ZN(n561) );
  NOR2_X1 U616 ( .A1(n550), .A2(n561), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n557) );
  NOR2_X1 U622 ( .A1(n555), .A2(n561), .ZN(n556) );
  XOR2_X1 U623 ( .A(n557), .B(n556), .Z(G1345GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n561), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1346GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  NAND2_X1 U629 ( .A1(n576), .A2(n568), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT123), .Z(n566) );
  NAND2_X1 U632 ( .A1(n568), .A2(n584), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT58), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n578) );
  INV_X1 U638 ( .A(n571), .ZN(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n575) );
  INV_X1 U640 ( .A(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n589) );
  INV_X1 U642 ( .A(n589), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n585), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U647 ( .A1(n585), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(KEYINPUT126), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

