//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT66), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT67), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(G2105), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n465), .A3(KEYINPUT3), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n463), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n475), .A2(G137), .A3(new_n476), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n471), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  INV_X1    g058(.A(G100), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n484), .A2(new_n476), .A3(KEYINPUT70), .ZN(new_n485));
  AOI21_X1  g060(.A(KEYINPUT70), .B1(new_n484), .B2(new_n476), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G112), .B2(new_n476), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n475), .A2(new_n476), .A3(new_n480), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n475), .A2(G2105), .A3(new_n480), .ZN(new_n491));
  OAI221_X1 g066(.A(new_n487), .B1(new_n488), .B2(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  OR2_X1    g071(.A1(new_n476), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G126), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n491), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR4_X1   g078(.A1(new_n467), .A2(KEYINPUT4), .A3(new_n503), .A4(G2105), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n480), .A2(new_n472), .A3(new_n474), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n504), .B1(new_n507), .B2(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n506), .A2(new_n509), .A3(KEYINPUT4), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n502), .B1(new_n508), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n516), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT5), .B(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(new_n515), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n519), .A2(new_n518), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n513), .A2(new_n514), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n533), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n515), .A2(G52), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n542), .B2(new_n522), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n526), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(new_n515), .A2(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(new_n522), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n526), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  OAI211_X1 g134(.A(G53), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT74), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT75), .B1(new_n560), .B2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n515), .A2(new_n564), .A3(new_n565), .A4(G53), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n560), .A2(new_n567), .A3(KEYINPUT9), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n562), .A2(new_n563), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n534), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n522), .A2(KEYINPUT76), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n535), .A2(new_n524), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(G91), .A3(new_n576), .ZN(new_n577));
  AND4_X1   g152(.A1(new_n559), .A2(new_n569), .A3(new_n573), .A4(new_n577), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n577), .A2(new_n573), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n559), .B1(new_n579), .B2(new_n569), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n578), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND2_X1  g158(.A1(new_n515), .A2(G49), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT78), .Z(new_n585));
  NAND3_X1  g160(.A1(new_n574), .A2(G87), .A3(new_n576), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n534), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G48), .B2(new_n515), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n574), .A2(G86), .A3(new_n576), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT79), .Z(G305));
  INV_X1    g170(.A(new_n522), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G85), .B1(G47), .B2(new_n515), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n526), .B2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n534), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n515), .A2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n574), .A2(G92), .A3(new_n576), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n574), .A2(KEYINPUT10), .A3(G92), .A4(new_n576), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n600), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n600), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  AND4_X1   g189(.A1(new_n563), .A2(new_n562), .A3(new_n566), .A4(new_n568), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n577), .A2(new_n573), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT77), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n579), .A2(new_n559), .A3(new_n569), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n614), .B1(new_n619), .B2(G868), .ZN(G297));
  XOR2_X1   g195(.A(G297), .B(KEYINPUT80), .Z(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n611), .B1(new_n622), .B2(G860), .ZN(G148));
  INV_X1    g198(.A(new_n552), .ZN(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n611), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n626), .B1(new_n628), .B2(new_n625), .ZN(G323));
  XOR2_X1   g204(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n630));
  XNOR2_X1  g205(.A(G323), .B(new_n630), .ZN(G282));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n476), .ZN(new_n633));
  INV_X1    g208(.A(G135), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n633), .B1(new_n488), .B2(new_n634), .C1(new_n635), .C2(new_n491), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n637), .A2(new_n638), .A3(new_n642), .ZN(G156));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NOR2_X1   g235(.A1(G2072), .A2(G2078), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n444), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n663), .B2(KEYINPUT82), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(KEYINPUT82), .B2(new_n663), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n662), .B(KEYINPUT17), .ZN(new_n668));
  INV_X1    g243(.A(new_n660), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n665), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n667), .A2(new_n662), .A3(new_n669), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n669), .A3(new_n666), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT83), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT84), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n681), .A2(new_n683), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n679), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n687), .A2(new_n684), .A3(new_n679), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n685), .B1(new_n684), .B2(new_n679), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT86), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1981), .B(G1986), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(G229));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT90), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT32), .B(G1981), .Z(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G23), .ZN(new_n707));
  INV_X1    g282(.A(G288), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n706), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT33), .B(G1976), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n706), .A2(G22), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G166), .B2(new_n706), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1971), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n704), .A2(new_n705), .A3(new_n711), .A4(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n719));
  NOR2_X1   g294(.A1(G25), .A2(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(KEYINPUT88), .B1(G95), .B2(G2105), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g297(.A1(KEYINPUT88), .A2(G95), .A3(G2105), .ZN(new_n723));
  OAI221_X1 g298(.A(G2104), .B1(G107), .B2(new_n476), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT89), .Z(new_n725));
  INV_X1    g300(.A(new_n488), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G131), .ZN(new_n727));
  INV_X1    g302(.A(new_n491), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G119), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n725), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n720), .B1(new_n731), .B2(G29), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n706), .A2(G24), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G290), .B2(G16), .ZN(new_n737));
  INV_X1    g312(.A(G1986), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT92), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(KEYINPUT36), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n738), .B2(new_n737), .ZN(new_n741));
  INV_X1    g316(.A(new_n732), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n733), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n718), .A2(new_n719), .A3(new_n735), .A4(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n739), .B1(KEYINPUT91), .B2(KEYINPUT36), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NOR2_X1   g322(.A1(G168), .A2(new_n706), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n706), .B2(G21), .ZN(new_n749));
  INV_X1    g324(.A(G1966), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n706), .A2(G5), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G171), .B2(new_n706), .ZN(new_n752));
  OAI22_X1  g327(.A1(new_n749), .A2(new_n750), .B1(G1961), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n750), .B2(new_n749), .ZN(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n636), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT95), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n706), .A2(G19), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n552), .B2(new_n706), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1341), .Z(new_n760));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(G28), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n755), .B1(new_n761), .B2(G28), .ZN(new_n763));
  AND2_X1   g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  NOR2_X1   g339(.A1(KEYINPUT31), .A2(G11), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n762), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n752), .B2(G1961), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n754), .A2(new_n757), .A3(new_n760), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n755), .A2(G27), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT97), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n508), .A2(new_n510), .ZN(new_n771));
  INV_X1    g346(.A(new_n502), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n770), .B1(new_n773), .B2(G29), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n768), .B1(new_n443), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n443), .B2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n755), .A2(G35), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G162), .B2(new_n755), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT29), .B(G2090), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT26), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n783), .A2(new_n784), .B1(G105), .B2(new_n470), .ZN(new_n785));
  INV_X1    g360(.A(G141), .ZN(new_n786));
  INV_X1    g361(.A(G129), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n785), .B1(new_n488), .B2(new_n786), .C1(new_n787), .C2(new_n491), .ZN(new_n788));
  MUX2_X1   g363(.A(G32), .B(new_n788), .S(G29), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT27), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1996), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n706), .A2(G4), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n611), .B2(new_n706), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1348), .ZN(new_n794));
  INV_X1    g369(.A(G34), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(KEYINPUT24), .ZN(new_n796));
  AOI21_X1  g371(.A(G29), .B1(new_n795), .B2(KEYINPUT24), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(KEYINPUT94), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(KEYINPUT94), .B2(new_n797), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n482), .B2(new_n755), .ZN(new_n800));
  INV_X1    g375(.A(G2084), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT96), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n755), .A2(G33), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT25), .Z(new_n806));
  AND2_X1   g381(.A1(new_n464), .A2(new_n466), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n807), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n808));
  INV_X1    g383(.A(G139), .ZN(new_n809));
  OAI221_X1 g384(.A(new_n806), .B1(new_n808), .B2(new_n476), .C1(new_n488), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n804), .B1(new_n810), .B2(G29), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(new_n442), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n801), .B2(new_n800), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n442), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n794), .A2(new_n803), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n755), .A2(G26), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT28), .ZN(new_n817));
  OR2_X1    g392(.A1(G104), .A2(G2105), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n819));
  INV_X1    g394(.A(G140), .ZN(new_n820));
  INV_X1    g395(.A(G128), .ZN(new_n821));
  OAI221_X1 g396(.A(new_n819), .B1(new_n488), .B2(new_n820), .C1(new_n821), .C2(new_n491), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n822), .A2(KEYINPUT93), .A3(G29), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT93), .B1(new_n822), .B2(G29), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n817), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(G2067), .Z(new_n826));
  NAND4_X1  g401(.A1(new_n780), .A2(new_n791), .A3(new_n815), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n706), .A2(G20), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT23), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n619), .B2(new_n706), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1956), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n776), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n746), .A2(new_n747), .A3(new_n832), .ZN(G150));
  INV_X1    g408(.A(G150), .ZN(G311));
  AOI22_X1  g409(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  OR3_X1    g410(.A1(new_n835), .A2(KEYINPUT99), .A3(new_n526), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT99), .B1(new_n835), .B2(new_n526), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n596), .A2(G93), .B1(G55), .B2(new_n515), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n611), .A2(G559), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n839), .A2(new_n624), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n839), .A2(new_n624), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n844), .B(new_n847), .Z(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  INV_X1    g425(.A(G860), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n841), .B1(new_n850), .B2(new_n852), .ZN(G145));
  XNOR2_X1  g428(.A(G164), .B(new_n822), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n810), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n788), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n730), .B(new_n640), .ZN(new_n857));
  OR2_X1    g432(.A1(G106), .A2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n858), .B(G2104), .C1(G118), .C2(new_n476), .ZN(new_n859));
  INV_X1    g434(.A(G142), .ZN(new_n860));
  INV_X1    g435(.A(G130), .ZN(new_n861));
  OAI221_X1 g436(.A(new_n859), .B1(new_n488), .B2(new_n860), .C1(new_n861), .C2(new_n491), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n857), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n856), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n856), .A2(new_n865), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n636), .B(G160), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n495), .B(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n856), .B2(new_n863), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n856), .B2(new_n863), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g450(.A(G305), .B(G288), .ZN(new_n876));
  XNOR2_X1  g451(.A(G303), .B(G290), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT42), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n847), .B(new_n628), .Z(new_n881));
  OAI21_X1  g456(.A(new_n627), .B1(new_n578), .B2(new_n580), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n617), .A2(new_n618), .A3(new_n611), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(G299), .A2(KEYINPUT101), .A3(new_n611), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(KEYINPUT41), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n882), .A2(new_n892), .A3(new_n884), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n619), .A2(KEYINPUT102), .A3(new_n627), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n890), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n894), .B1(new_n885), .B2(new_n886), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(KEYINPUT103), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n889), .B1(new_n900), .B2(new_n881), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n880), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n901), .A2(new_n902), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(new_n879), .ZN(new_n907));
  OAI21_X1  g482(.A(G868), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n839), .A2(new_n625), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(G295));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n908), .A2(new_n911), .A3(new_n909), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n911), .B1(new_n908), .B2(new_n909), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(G331));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n915));
  OAI21_X1  g490(.A(G286), .B1(G171), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(G171), .A2(new_n915), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n916), .B(new_n917), .Z(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n847), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT109), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n916), .B(new_n917), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(new_n846), .A3(new_n845), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n888), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT103), .B1(new_n924), .B2(new_n898), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n891), .A2(new_n890), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n919), .A2(new_n922), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT108), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  AOI211_X1 g506(.A(new_n931), .B(new_n928), .C1(new_n925), .C2(new_n926), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n878), .B(new_n923), .C1(new_n930), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT110), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n929), .B1(new_n897), .B2(new_n899), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n931), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n927), .A2(KEYINPUT108), .A3(new_n929), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n878), .A4(new_n923), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n923), .B1(new_n930), .B2(new_n932), .ZN(new_n941));
  INV_X1    g516(.A(new_n878), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n934), .A2(new_n940), .A3(new_n943), .A4(new_n873), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n933), .B2(KEYINPUT110), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n888), .A2(new_n922), .A3(new_n919), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n920), .A2(new_n922), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n893), .A2(KEYINPUT41), .A3(new_n895), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n888), .A2(KEYINPUT41), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n942), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n946), .A2(new_n953), .A3(new_n954), .A4(new_n940), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n945), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n946), .A2(new_n954), .A3(new_n940), .A4(new_n943), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n946), .A2(new_n940), .A3(new_n953), .ZN(new_n960));
  OAI211_X1 g535(.A(KEYINPUT44), .B(new_n959), .C1(new_n960), .C2(new_n954), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(G397));
  INV_X1    g537(.A(KEYINPUT120), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n471), .A2(new_n481), .A3(G40), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT111), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n471), .A2(new_n481), .A3(new_n967), .A4(G40), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n773), .A2(new_n964), .A3(new_n966), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n708), .A2(G1976), .ZN(new_n970));
  INV_X1    g545(.A(G1976), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(G288), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n969), .A2(new_n970), .A3(G8), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1981), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n592), .A2(new_n593), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n515), .A2(G48), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n535), .A2(new_n524), .A3(G86), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n976), .B(new_n977), .C1(new_n978), .C2(new_n526), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G1981), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n975), .A2(new_n980), .A3(KEYINPUT49), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT49), .B1(new_n975), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n969), .A2(G8), .A3(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n969), .A2(new_n970), .A3(G8), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n973), .B(new_n984), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(G164), .B2(G1384), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n966), .A2(new_n968), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n506), .A2(new_n509), .A3(KEYINPUT4), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n509), .B1(new_n506), .B2(KEYINPUT4), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n991), .A2(new_n992), .A3(new_n504), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT45), .B(new_n964), .C1(new_n993), .C2(new_n502), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(new_n990), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1971), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n773), .A2(new_n998), .A3(new_n964), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1000));
  XOR2_X1   g575(.A(KEYINPUT114), .B(G2090), .Z(new_n1001));
  NAND4_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n990), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G8), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT116), .ZN(new_n1006));
  NAND3_X1  g581(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT115), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n987), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n995), .A2(new_n750), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n999), .A2(new_n1000), .A3(new_n801), .A4(new_n990), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(G286), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n997), .B2(new_n1002), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1018), .A2(KEYINPUT117), .A3(new_n1009), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT117), .B1(new_n1018), .B2(new_n1009), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1011), .B(new_n1016), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT118), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT63), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1003), .A2(G8), .A3(new_n1009), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1018), .A2(KEYINPUT117), .A3(new_n1009), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1029), .A2(new_n1030), .A3(new_n1011), .A4(new_n1016), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1029), .A2(new_n987), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G164), .A2(G1384), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1017), .B1(new_n1034), .B2(new_n990), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n984), .A2(new_n971), .A3(new_n708), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n975), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1033), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT119), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT63), .B1(new_n1021), .B2(KEYINPUT118), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1031), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n963), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1022), .A2(new_n1024), .A3(new_n1031), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1040), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(KEYINPUT120), .A3(new_n1032), .A4(new_n1038), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G286), .A2(G8), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT123), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1015), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1014), .B2(new_n1049), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1015), .A2(new_n1052), .A3(new_n1050), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(KEYINPUT62), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT62), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1029), .A2(new_n1011), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n995), .B2(G2078), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n999), .A2(new_n1000), .A3(new_n990), .ZN(new_n1062));
  INV_X1    g637(.A(G1961), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1060), .A2(G2078), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n989), .A2(new_n990), .A3(new_n994), .A4(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G171), .ZN(new_n1068));
  NOR4_X1   g643(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1070));
  INV_X1    g645(.A(new_n965), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n989), .A2(new_n1071), .A3(new_n994), .A4(new_n1065), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1061), .A2(G301), .A3(new_n1064), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT125), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1068), .A2(KEYINPUT125), .A3(new_n1073), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n985), .A2(new_n986), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n973), .A2(new_n984), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1079), .B(new_n1080), .C1(new_n1018), .C2(new_n1009), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1061), .A2(new_n1064), .A3(new_n1072), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT126), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT126), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1061), .A2(new_n1085), .A3(new_n1064), .A4(new_n1072), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(G171), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1061), .A2(G301), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1088), .A2(KEYINPUT54), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1017), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1091), .A2(KEYINPUT51), .A3(new_n1049), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1078), .A2(new_n1082), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n579), .A2(new_n569), .B1(KEYINPUT121), .B2(KEYINPUT57), .ZN(new_n1095));
  NOR2_X1   g670(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1956), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1062), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n989), .A2(new_n990), .A3(new_n994), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1099), .A2(new_n1097), .A3(new_n1101), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n969), .A2(G2067), .ZN(new_n1106));
  INV_X1    g681(.A(G1348), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n1062), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n627), .B1(new_n1108), .B2(KEYINPUT60), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1062), .A2(new_n1107), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1110), .B1(new_n1111), .B2(new_n1106), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1104), .A2(new_n1105), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  NOR4_X1   g688(.A1(new_n1111), .A2(new_n1110), .A3(new_n611), .A4(new_n1106), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n969), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n995), .B2(G1996), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1117), .A2(KEYINPUT59), .A3(new_n552), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT59), .B1(new_n1117), .B2(new_n552), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1114), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1105), .A2(KEYINPUT122), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1099), .A2(new_n1097), .A3(new_n1122), .A4(new_n1101), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1102), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1113), .B(new_n1120), .C1(KEYINPUT61), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1108), .A2(new_n627), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(new_n1102), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1094), .A2(KEYINPUT127), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1082), .A2(new_n1093), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(new_n1090), .A4(new_n1078), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1069), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1043), .A2(new_n1047), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n989), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1135), .A2(new_n990), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n822), .B(G2067), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT112), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n788), .B(G1996), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n730), .B(new_n734), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT113), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1136), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(G290), .B(G1986), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1136), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1134), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1136), .ZN(new_n1149));
  OR3_X1    g724(.A1(new_n1149), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT46), .B1(new_n1149), .B2(G1996), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1137), .A2(new_n788), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1150), .A2(new_n1151), .B1(new_n1136), .B2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT47), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1141), .A2(new_n731), .A3(new_n733), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n822), .A2(G2067), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1149), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1145), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1149), .A2(G1986), .A3(G290), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT48), .Z(new_n1160));
  AOI211_X1 g735(.A(new_n1154), .B(new_n1157), .C1(new_n1158), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1148), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g737(.A(G319), .B1(new_n657), .B2(new_n658), .ZN(new_n1164));
  NOR3_X1   g738(.A1(G229), .A2(G227), .A3(new_n1164), .ZN(new_n1165));
  AND3_X1   g739(.A1(new_n956), .A2(new_n874), .A3(new_n1165), .ZN(G308));
  NAND3_X1  g740(.A1(new_n956), .A2(new_n874), .A3(new_n1165), .ZN(G225));
endmodule


