//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n459), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n459), .A2(G137), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(new_n463), .B1(G101), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n464), .A2(new_n468), .ZN(G160));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n463), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(G124), .A2(new_n473), .B1(new_n474), .B2(G136), .ZN(new_n475));
  OAI221_X1 g050(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G162));
  XNOR2_X1  g053(.A(KEYINPUT69), .B(KEYINPUT4), .ZN(new_n479));
  OAI21_X1  g054(.A(G138), .B1(new_n470), .B2(new_n471), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT67), .B(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n463), .A2(new_n459), .A3(G138), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AND2_X1   g063(.A1(G126), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n470), .B2(new_n471), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(KEYINPUT68), .B(new_n489), .C1(new_n470), .C2(new_n471), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n485), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G62), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n503), .A2(new_n504), .B1(G75), .B2(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n502), .A2(KEYINPUT70), .A3(G62), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n497), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n499), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  INV_X1    g088(.A(new_n501), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n508), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n512), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n507), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(new_n511), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n502), .ZN(new_n525));
  OAI21_X1  g100(.A(G89), .B1(new_n516), .B2(new_n508), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n524), .A2(new_n528), .ZN(G168));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n530), .B(new_n531), .C1(new_n525), .C2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(new_n500), .B2(new_n501), .ZN(new_n534));
  INV_X1    g109(.A(new_n531), .ZN(new_n535));
  OAI21_X1  g110(.A(KEYINPUT71), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(G651), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n509), .A2(new_n510), .B1(new_n500), .B2(new_n501), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT72), .B(G90), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n538), .A2(new_n539), .B1(new_n511), .B2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n537), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n500), .B2(new_n501), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(KEYINPUT73), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(G56), .B1(new_n514), .B2(new_n515), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(new_n549), .A3(new_n545), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(G651), .A3(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n538), .A2(G81), .B1(new_n511), .B2(G43), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n511), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n525), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n564), .A2(G651), .B1(G91), .B2(new_n538), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n538), .A2(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n511), .A2(G49), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n511), .A2(G48), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n574), .B2(new_n497), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n538), .A2(KEYINPUT74), .A3(G86), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n517), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n576), .A2(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n511), .A2(G47), .ZN(new_n583));
  XNOR2_X1  g158(.A(KEYINPUT75), .B(G85), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n517), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n497), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n538), .A2(KEYINPUT10), .A3(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n517), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n591), .A2(new_n594), .B1(G54), .B2(new_n511), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n500), .B2(new_n501), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n598));
  AND2_X1   g173(.A1(G79), .A2(G543), .ZN(new_n599));
  OR3_X1    g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n597), .B2(new_n599), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n600), .A2(G651), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n590), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n590), .B1(new_n604), .B2(G868), .ZN(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n459), .A2(new_n467), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  AOI22_X1  g195(.A1(G123), .A2(new_n473), .B1(new_n474), .B2(G135), .ZN(new_n621));
  OAI221_X1 g196(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n463), .C2(G111), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT77), .Z(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n625), .A2(G2096), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(G2096), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT78), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(G14), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n641), .ZN(G401));
  XNOR2_X1  g220(.A(G2084), .B(G2090), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT79), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n648), .B(KEYINPUT17), .Z(new_n651));
  INV_X1    g226(.A(new_n649), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n646), .B(new_n650), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n646), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n649), .A2(new_n646), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n653), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(new_n666), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n663), .A2(new_n668), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT80), .B(KEYINPUT20), .Z(new_n671));
  OAI221_X1 g246(.A(new_n667), .B1(new_n669), .B2(new_n663), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n670), .B2(new_n671), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT81), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT82), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G229));
  NAND3_X1  g257(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT25), .Z(new_n684));
  NAND2_X1  g259(.A1(new_n474), .A2(G139), .ZN(new_n685));
  AOI22_X1  g260(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n684), .B(new_n685), .C1(new_n463), .C2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT90), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n689), .B2(G33), .ZN(new_n691));
  INV_X1    g266(.A(G2072), .ZN(new_n692));
  OAI21_X1  g267(.A(KEYINPUT92), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n691), .A2(KEYINPUT92), .A3(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT91), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n691), .A2(KEYINPUT91), .A3(new_n692), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n693), .A2(new_n694), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G5), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G171), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G1961), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT98), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(G1961), .ZN(new_n705));
  INV_X1    g280(.A(G34), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(KEYINPUT24), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n706), .B2(KEYINPUT24), .ZN(new_n708));
  AOI22_X1  g283(.A1(G160), .A2(G29), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(G2084), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(G2084), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n621), .A2(G29), .A3(new_n622), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT30), .B(G28), .ZN(new_n713));
  OR2_X1    g288(.A1(KEYINPUT31), .A2(G11), .ZN(new_n714));
  NAND2_X1  g289(.A1(KEYINPUT31), .A2(G11), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n713), .A2(new_n689), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n710), .A2(new_n711), .A3(new_n712), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n689), .A2(G27), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G164), .B2(new_n689), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G2078), .ZN(new_n720));
  NOR4_X1   g295(.A1(new_n704), .A2(new_n705), .A3(new_n717), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n689), .A2(G32), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n473), .A2(G129), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT93), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n467), .A2(G105), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT26), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n725), .B(new_n727), .C1(G141), .C2(new_n474), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT94), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n722), .B1(new_n731), .B2(new_n689), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT95), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n732), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G21), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G168), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT96), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT97), .B(G1966), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n721), .A2(new_n735), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n699), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT99), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n699), .A2(new_n741), .A3(KEYINPUT99), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n689), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n689), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT29), .Z(new_n748));
  INV_X1    g323(.A(G2090), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G4), .A2(G16), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT87), .Z(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n603), .B2(new_n700), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT88), .B(G1348), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n689), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n473), .A2(G128), .ZN(new_n758));
  OAI221_X1 g333(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n463), .C2(G116), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n474), .A2(G140), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G29), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n762), .A2(KEYINPUT89), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(KEYINPUT89), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n757), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n750), .B(new_n755), .C1(G2067), .C2(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n700), .A2(KEYINPUT83), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n700), .A2(KEYINPUT83), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n767), .A2(G20), .A3(new_n768), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT23), .Z(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G299), .B2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1956), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n765), .A2(G2067), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n772), .B(new_n773), .C1(new_n748), .C2(new_n749), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n767), .A2(new_n768), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(G19), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n554), .B2(new_n775), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1341), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n766), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n744), .A2(new_n745), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n689), .A2(G25), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n473), .A2(G119), .ZN(new_n783));
  OAI221_X1 g358(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n474), .A2(G131), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n782), .B1(new_n787), .B2(new_n689), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT35), .B(G1991), .Z(new_n789));
  XOR2_X1   g364(.A(new_n788), .B(new_n789), .Z(new_n790));
  NOR2_X1   g365(.A1(new_n775), .A2(G24), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n588), .B2(new_n775), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1986), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n775), .A2(G22), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n775), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1971), .ZN(new_n797));
  MUX2_X1   g372(.A(G6), .B(G305), .S(G16), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT84), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT32), .B(G1981), .Z(new_n800));
  AOI21_X1  g375(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n700), .A2(G23), .ZN(new_n802));
  INV_X1    g377(.A(G288), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n700), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT33), .B(G1976), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT85), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n801), .B(new_n807), .C1(new_n799), .C2(new_n800), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n794), .B1(new_n808), .B2(KEYINPUT34), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT86), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n781), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n781), .A3(new_n812), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n780), .B1(new_n814), .B2(new_n815), .ZN(G311));
  INV_X1    g391(.A(new_n780), .ZN(new_n817));
  INV_X1    g392(.A(new_n815), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n813), .ZN(G150));
  NAND2_X1  g394(.A1(G80), .A2(G543), .ZN(new_n820));
  INV_X1    g395(.A(G67), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n525), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G651), .ZN(new_n823));
  OAI211_X1 g398(.A(G55), .B(G543), .C1(new_n516), .C2(new_n508), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n517), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G860), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT37), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n604), .A2(G559), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n553), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n551), .A2(new_n552), .A3(new_n823), .A4(new_n827), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n832), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT100), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n836), .B2(new_n837), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n830), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT101), .Z(G145));
  XOR2_X1   g418(.A(G160), .B(new_n623), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n477), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n492), .A2(new_n493), .ZN(new_n846));
  INV_X1    g421(.A(new_n488), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT102), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n849));
  AOI211_X1 g424(.A(new_n849), .B(new_n488), .C1(new_n492), .C2(new_n493), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n485), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n729), .B(KEYINPUT94), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(new_n761), .ZN(new_n853));
  INV_X1    g428(.A(new_n761), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n731), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n688), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n688), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n851), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  INV_X1    g436(.A(new_n485), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT68), .B1(new_n459), .B2(new_n489), .ZN(new_n863));
  INV_X1    g438(.A(new_n493), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n847), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n849), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n494), .A2(KEYINPUT102), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n868), .A3(new_n857), .ZN(new_n869));
  AOI22_X1  g444(.A1(G130), .A2(new_n473), .B1(new_n474), .B2(G142), .ZN(new_n870));
  OAI221_X1 g445(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n463), .C2(G118), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n618), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n786), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT103), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n860), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n860), .B2(new_n869), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n845), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n860), .A2(new_n869), .A3(new_n874), .ZN(new_n879));
  INV_X1    g454(.A(new_n845), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n860), .A2(new_n869), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n879), .B(new_n880), .C1(new_n881), .C2(new_n875), .ZN(new_n882));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n878), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(G395));
  NAND2_X1  g461(.A1(new_n828), .A2(new_n607), .ZN(new_n887));
  NAND3_X1  g462(.A1(G290), .A2(new_n576), .A3(new_n581), .ZN(new_n888));
  NAND2_X1  g463(.A1(G305), .A2(new_n588), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(G166), .A2(G288), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n803), .B1(new_n507), .B2(new_n518), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n888), .A2(new_n891), .A3(new_n892), .A4(new_n889), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT42), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n894), .A2(KEYINPUT106), .A3(new_n895), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT106), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n896), .B1(new_n900), .B2(KEYINPUT42), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n613), .B(new_n835), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n561), .A2(new_n595), .A3(new_n602), .A4(new_n565), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n561), .A2(new_n565), .B1(new_n595), .B2(new_n602), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n902), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n904), .B2(new_n905), .ZN(new_n910));
  NAND2_X1  g485(.A1(G299), .A2(new_n603), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n903), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n907), .A2(KEYINPUT105), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(KEYINPUT105), .B2(new_n907), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n901), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n887), .B1(new_n916), .B2(new_n607), .ZN(G295));
  OAI21_X1  g492(.A(new_n887), .B1(new_n916), .B2(new_n607), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  NAND2_X1  g495(.A1(G301), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n537), .A2(KEYINPUT107), .A3(new_n540), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n828), .A2(new_n553), .ZN(new_n923));
  AOI22_X1  g498(.A1(new_n823), .A2(new_n827), .B1(new_n551), .B2(new_n552), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n921), .B(new_n922), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n537), .A2(KEYINPUT107), .A3(new_n540), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT107), .B1(new_n537), .B2(new_n540), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n834), .B(new_n833), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G286), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n925), .A2(new_n928), .A3(G168), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n906), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n910), .A2(new_n912), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n930), .B2(new_n931), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n931), .ZN(new_n937));
  AOI21_X1  g512(.A(G168), .B1(new_n925), .B2(new_n928), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n913), .B(new_n935), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n900), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n913), .B1(new_n937), .B2(new_n938), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n899), .A2(new_n944), .A3(new_n932), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n883), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n900), .B(KEYINPUT109), .C1(new_n936), .C2(new_n940), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n943), .A2(KEYINPUT43), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n899), .B1(new_n944), .B2(new_n932), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT44), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n943), .A2(new_n950), .A3(new_n947), .A4(new_n948), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n946), .B2(new_n951), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n919), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n949), .B2(new_n952), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT44), .B1(new_n955), .B2(new_n956), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n961), .A2(new_n962), .A3(KEYINPUT110), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n960), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT45), .B1(new_n851), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n464), .A2(new_n468), .A3(G40), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n852), .A2(G1996), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n761), .B(G2067), .Z(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n970), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT111), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n787), .A2(new_n789), .ZN(new_n978));
  OAI22_X1  g553(.A1(new_n977), .A2(new_n978), .B1(G2067), .B2(new_n761), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n976), .B(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n786), .B(new_n789), .Z(new_n982));
  NAND2_X1  g557(.A1(new_n970), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n969), .A2(G1986), .A3(G290), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT48), .Z(new_n986));
  AOI22_X1  g561(.A1(new_n970), .A2(new_n979), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n969), .B1(new_n731), .B2(new_n974), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT124), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n969), .B2(G1996), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n970), .A2(KEYINPUT46), .A3(new_n971), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n993), .B(new_n994), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT126), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n993), .B(new_n994), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n987), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT123), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT62), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n851), .A2(new_n1003), .A3(new_n965), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G2084), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n851), .A2(KEYINPUT112), .A3(new_n1003), .A4(new_n965), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n495), .A2(new_n965), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n967), .B1(new_n1009), .B2(KEYINPUT50), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT113), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n495), .A2(new_n1014), .A3(KEYINPUT45), .A4(new_n965), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n968), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n739), .B1(new_n1016), .B2(new_n966), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1011), .A2(new_n1017), .A3(G168), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G168), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT51), .B1(new_n1018), .B2(G8), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1002), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n868), .B2(G1384), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n1027), .B(G1384), .C1(new_n485), .C2(new_n494), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n967), .B1(new_n1029), .B2(new_n1014), .ZN(new_n1030));
  INV_X1    g605(.A(G2078), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .A4(new_n1013), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT119), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1015), .A2(new_n968), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n485), .B2(new_n494), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1014), .B1(new_n1035), .B2(KEYINPUT45), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1031), .A4(new_n1028), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1033), .A2(KEYINPUT53), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1006), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1041));
  INV_X1    g616(.A(G1961), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n851), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n967), .B1(new_n1009), .B2(new_n1027), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1031), .A3(new_n1045), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1041), .A2(new_n1042), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1040), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G171), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1006), .A2(new_n749), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1971), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G166), .A2(new_n1020), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT55), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(G8), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1003), .B1(new_n851), .B2(new_n965), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1035), .A2(new_n1003), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n968), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1057), .A2(new_n1059), .A3(G2090), .ZN(new_n1060));
  OAI21_X1  g635(.A(G8), .B1(new_n1060), .B2(new_n1051), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1055), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n851), .A2(new_n968), .A3(new_n965), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n803), .A2(G1976), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(G8), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(G288), .B2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1064), .A2(G8), .A3(new_n1065), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1981), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n576), .A2(new_n581), .A3(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n517), .A2(new_n579), .ZN(new_n1073));
  OAI21_X1  g648(.A(G1981), .B1(new_n575), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1072), .A2(KEYINPUT49), .A3(new_n1074), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1064), .A3(G8), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1067), .A2(new_n1070), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1056), .A2(new_n1063), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1049), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1018), .A2(G8), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1019), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G286), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1088), .A3(KEYINPUT62), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1026), .A2(new_n1083), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT63), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1086), .A2(G8), .A3(G168), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1082), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1020), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1080), .B1(new_n1094), .B2(new_n1055), .ZN(new_n1095));
  AND4_X1   g670(.A1(KEYINPUT63), .A2(new_n1086), .A3(G8), .A4(G168), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1062), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1095), .B(new_n1096), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1093), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1056), .A2(new_n1080), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1064), .A2(G8), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1079), .A2(new_n1068), .A3(new_n803), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(new_n1072), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1090), .A2(new_n1101), .A3(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1085), .A2(new_n1088), .A3(new_n1063), .A4(new_n1095), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1046), .A2(new_n1043), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT53), .B1(new_n1031), .B2(KEYINPUT121), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(KEYINPUT121), .B2(new_n1031), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n967), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1114), .B2(new_n967), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n1044), .A3(new_n1028), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1110), .A2(new_n1111), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1109), .B1(new_n1118), .B2(G301), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1047), .A2(new_n1117), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1048), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n1124), .B2(G301), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1108), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1956), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1044), .A2(new_n1045), .A3(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1128), .A2(KEYINPUT115), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT115), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n1133));
  XNOR2_X1  g708(.A(G299), .B(new_n1133), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1348), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1041), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1064), .A2(G2067), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1128), .A2(new_n1130), .A3(new_n1134), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1141), .A2(new_n604), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1135), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1134), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(KEYINPUT117), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1141), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT117), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1144), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n968), .B1(new_n1035), .B2(new_n1003), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1153));
  AOI21_X1  g728(.A(G1348), .B1(new_n1153), .B2(new_n1008), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1151), .B1(new_n1154), .B2(new_n1138), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n1139), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(new_n604), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1150), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n603), .A4(new_n1139), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1044), .A2(new_n971), .A3(new_n1045), .ZN(new_n1160));
  XOR2_X1   g735(.A(KEYINPUT58), .B(G1341), .Z(new_n1161));
  NAND2_X1  g736(.A1(new_n1064), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n553), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1141), .A2(KEYINPUT118), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1128), .A2(new_n1167), .A3(new_n1130), .A4(new_n1134), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1166), .A2(KEYINPUT61), .A3(new_n1168), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1159), .B(new_n1165), .C1(new_n1135), .C2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1143), .B1(new_n1158), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1049), .B1(G171), .B2(new_n1120), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n1123), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1126), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1107), .A2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n588), .B(G1986), .Z(new_n1176));
  NAND2_X1  g751(.A1(new_n970), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n981), .A2(new_n1177), .A3(new_n983), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1001), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  AOI211_X1 g755(.A(KEYINPUT123), .B(new_n1178), .C1(new_n1107), .C2(new_n1174), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1000), .B1(new_n1180), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n1184));
  INV_X1    g758(.A(G319), .ZN(new_n1185));
  NOR3_X1   g759(.A1(G401), .A2(G227), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g760(.A(new_n1186), .ZN(new_n1187));
  OAI21_X1  g761(.A(new_n1184), .B1(G229), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n681), .A2(KEYINPUT127), .A3(new_n1186), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AND3_X1   g764(.A1(new_n1190), .A2(new_n884), .A3(new_n957), .ZN(G308));
  NAND3_X1  g765(.A1(new_n1190), .A2(new_n884), .A3(new_n957), .ZN(G225));
endmodule


