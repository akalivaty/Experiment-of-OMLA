//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT67), .Z(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT33), .ZN(new_n206));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n207), .B1(KEYINPUT23), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G169gat), .ZN(new_n210));
  INV_X1    g009(.A(G176gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT23), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217));
  OR2_X1    g016(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(G190gat), .A3(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT25), .A4(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n213), .A2(new_n222), .B1(new_n207), .B2(KEYINPUT23), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n210), .A2(new_n211), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n223), .A2(new_n220), .A3(new_n226), .A4(KEYINPUT25), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n220), .A3(new_n226), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n221), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(G127gat), .B(G134gat), .Z(new_n233));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n233), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(G113gat), .B(G120gat), .Z(new_n238));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(new_n235), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n225), .A2(KEYINPUT26), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT26), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n207), .B1(new_n244), .B2(new_n208), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n246), .A2(KEYINPUT28), .A3(new_n213), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT28), .B1(new_n246), .B2(new_n213), .ZN(new_n248));
  OAI221_X1 g047(.A(new_n242), .B1(new_n243), .B2(new_n245), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n241), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n241), .B1(new_n232), .B2(new_n249), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n232), .A2(KEYINPUT66), .A3(new_n241), .A4(new_n249), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256));
  OAI211_X1 g055(.A(KEYINPUT32), .B(new_n206), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n253), .B2(new_n254), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT32), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n204), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n258), .A2(KEYINPUT33), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n253), .A2(new_n256), .A3(new_n254), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(KEYINPUT69), .A3(KEYINPUT34), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT34), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n253), .A2(new_n264), .A3(new_n256), .A4(new_n254), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT69), .B1(new_n262), .B2(KEYINPUT34), .ZN(new_n267));
  OAI221_X1 g066(.A(new_n257), .B1(new_n260), .B2(new_n261), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n266), .A2(new_n267), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT71), .A4(new_n272), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n266), .B2(new_n267), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(new_n270), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n275), .A2(new_n276), .B1(new_n279), .B2(KEYINPUT36), .ZN(new_n280));
  AND2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT75), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G155gat), .ZN(new_n284));
  INV_X1    g083(.A(G162gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n287));
  NAND2_X1  g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(KEYINPUT2), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n283), .A2(new_n289), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT2), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT2), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT74), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n288), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT73), .B1(new_n281), .B2(new_n282), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n302), .A3(new_n288), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n300), .A2(new_n292), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT3), .B1(new_n295), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n301), .A2(new_n303), .ZN(new_n307));
  XNOR2_X1  g106(.A(G141gat), .B(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n298), .A2(KEYINPUT74), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n296), .A2(KEYINPUT2), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n308), .B1(new_n288), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n306), .B(new_n294), .C1(new_n307), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n237), .A2(new_n240), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n305), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G225gat), .A2(G233gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT4), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n294), .B1(new_n307), .B2(new_n312), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(new_n314), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n300), .A2(new_n292), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n301), .A2(new_n303), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n322), .A4(new_n294), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n315), .A2(new_n316), .A3(new_n319), .A4(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(new_n314), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n322), .A2(new_n294), .A3(new_n237), .A4(new_n240), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n316), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n314), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n306), .B1(new_n322), .B2(new_n294), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n319), .B(new_n323), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n325), .A4(new_n316), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT76), .B1(new_n324), .B2(KEYINPUT5), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n331), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT0), .ZN(new_n341));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT6), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n331), .ZN(new_n346));
  INV_X1    g145(.A(new_n338), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n324), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n343), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(KEYINPUT6), .A3(new_n343), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G197gat), .B(G204gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT22), .ZN(new_n359));
  INV_X1    g158(.A(G211gat), .ZN(new_n360));
  INV_X1    g159(.A(G218gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G211gat), .B(G218gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n362), .B2(new_n358), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n232), .A2(new_n249), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n369), .B1(new_n232), .B2(new_n249), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n368), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n370), .ZN(new_n376));
  INV_X1    g175(.A(new_n368), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n232), .B2(new_n249), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n376), .B(new_n377), .C1(new_n370), .C2(new_n378), .ZN(new_n379));
  AOI211_X1 g178(.A(new_n354), .B(new_n357), .C1(new_n375), .C2(new_n379), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n375), .A2(new_n357), .A3(new_n379), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n380), .A2(KEYINPUT72), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT72), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n375), .A2(new_n379), .ZN(new_n384));
  INV_X1    g183(.A(new_n357), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(KEYINPUT30), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n375), .A2(new_n357), .A3(new_n379), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n385), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n354), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n353), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(KEYINPUT31), .B(G50gat), .Z(new_n393));
  INV_X1    g192(.A(G228gat), .ZN(new_n394));
  INV_X1    g193(.A(G233gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n313), .A2(new_n372), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n377), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n372), .B1(new_n366), .B2(new_n367), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(KEYINPUT77), .B(new_n372), .C1(new_n366), .C2(new_n367), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT3), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n295), .A2(new_n304), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n396), .B(new_n398), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G22gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n396), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n404), .B1(new_n306), .B2(new_n399), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n368), .B1(new_n313), .B2(new_n372), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n406), .B1(new_n405), .B2(new_n410), .ZN(new_n412));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n401), .A2(new_n402), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n404), .B1(new_n416), .B2(new_n306), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n396), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n410), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G22gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n413), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n393), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n414), .B1(new_n411), .B2(new_n412), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(new_n421), .A3(new_n413), .ZN(new_n425));
  INV_X1    g224(.A(new_n393), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n392), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n391), .A2(new_n387), .A3(new_n386), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n334), .A2(new_n329), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n326), .A2(new_n327), .A3(new_n316), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n432), .A2(KEYINPUT39), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n343), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n334), .A2(new_n435), .A3(new_n329), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT40), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n343), .A2(new_n349), .B1(new_n437), .B2(KEYINPUT78), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n431), .A2(new_n433), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n439), .A2(KEYINPUT40), .A3(new_n344), .A4(new_n436), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT79), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n434), .A2(KEYINPUT79), .A3(KEYINPUT40), .A4(new_n436), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n434), .A2(new_n436), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n446), .B2(KEYINPUT40), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n430), .A2(new_n438), .A3(new_n444), .A4(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n426), .B1(new_n424), .B2(new_n425), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n357), .B1(new_n375), .B2(new_n379), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n375), .A2(KEYINPUT37), .A3(new_n379), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n453), .A2(new_n357), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT38), .B1(new_n384), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n452), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n351), .A2(new_n457), .A3(new_n352), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT38), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(new_n357), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT80), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n460), .A2(new_n461), .B1(new_n455), .B2(new_n384), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n453), .A2(KEYINPUT80), .A3(new_n357), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n448), .B(new_n451), .C1(new_n458), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n429), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n280), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n351), .A2(new_n352), .B1(new_n354), .B2(new_n390), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n279), .A2(new_n451), .A3(new_n468), .A4(new_n389), .ZN(new_n469));
  INV_X1    g268(.A(new_n353), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT35), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n423), .A2(new_n471), .A3(new_n427), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n470), .A2(new_n472), .A3(new_n430), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n268), .A2(new_n271), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n469), .A2(KEYINPUT35), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G113gat), .B(G141gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT11), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(new_n210), .ZN(new_n479));
  INV_X1    g278(.A(G197gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT12), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT16), .ZN(new_n484));
  AOI21_X1  g283(.A(G1gat), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(KEYINPUT87), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(G8gat), .Z(new_n488));
  XOR2_X1   g287(.A(G43gat), .B(G50gat), .Z(new_n489));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT15), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT14), .ZN(new_n493));
  INV_X1    g292(.A(G29gat), .ZN(new_n494));
  INV_X1    g293(.A(G36gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT84), .B1(new_n494), .B2(new_n495), .ZN(new_n499));
  OR3_X1    g298(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT84), .ZN(new_n500));
  AND4_X1   g299(.A1(new_n492), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n489), .A2(new_n491), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n489), .A2(new_n491), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n502), .B1(new_n503), .B2(KEYINPUT83), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n496), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(KEYINPUT81), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n497), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT82), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n509), .A2(new_n510), .B1(G29gat), .B2(G36gat), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n503), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT17), .B(new_n505), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n488), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT86), .ZN(new_n517));
  INV_X1    g316(.A(new_n505), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n514), .B1(new_n511), .B2(new_n512), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT85), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT85), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n521), .B(new_n505), .C1(new_n513), .C2(new_n514), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n517), .B1(new_n523), .B2(KEYINPUT17), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT86), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n516), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n523), .A2(new_n488), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT18), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT88), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n488), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n523), .B(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n529), .B(KEYINPUT13), .Z(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n531), .B2(new_n533), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n482), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n531), .A2(new_n533), .ZN(new_n543));
  INV_X1    g342(.A(new_n482), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n543), .A2(new_n534), .A3(new_n540), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n476), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT89), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550));
  XNOR2_X1  g349(.A(G57gat), .B(G64gat), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G71gat), .B(G78gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT92), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n551), .A2(new_n552), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n558), .A2(new_n550), .A3(new_n554), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n554), .B1(new_n558), .B2(new_n550), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT92), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n536), .B1(new_n562), .B2(KEYINPUT21), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT93), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n555), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT91), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n571), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n565), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n564), .A3(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT96), .ZN(new_n583));
  OAI22_X1  g382(.A1(new_n583), .A2(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(KEYINPUT8), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(KEYINPUT95), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n588), .A2(new_n583), .A3(G85gat), .A4(G92gat), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n590), .A2(new_n591), .B1(new_n587), .B2(KEYINPUT95), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n586), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G99gat), .B(G106gat), .Z(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n586), .A2(new_n596), .A3(new_n589), .A4(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n515), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n599), .B1(new_n524), .B2(new_n526), .ZN(new_n600));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n523), .B2(new_n598), .ZN(new_n604));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605));
  OR3_X1    g404(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n600), .B2(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT94), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n612), .B1(new_n607), .B2(KEYINPUT97), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n606), .B(new_n607), .C1(KEYINPUT97), .C2(new_n612), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n582), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(G176gat), .B(G204gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n598), .A2(new_n555), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n595), .B(new_n597), .C1(new_n559), .C2(new_n560), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n598), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n561), .B2(new_n557), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n623), .A2(new_n626), .A3(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT98), .B1(new_n630), .B2(new_n622), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n632));
  INV_X1    g431(.A(new_n622), .ZN(new_n633));
  AOI211_X1 g432(.A(new_n632), .B(new_n633), .C1(new_n628), .C2(new_n629), .ZN(new_n634));
  OAI221_X1 g433(.A(new_n621), .B1(new_n622), .B2(new_n625), .C1(new_n631), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n622), .B(KEYINPUT99), .Z(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n628), .B2(new_n629), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n625), .A2(new_n622), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n620), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n617), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n549), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n470), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n430), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(G8gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT42), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT16), .B(G8gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  MUX2_X1   g449(.A(new_n648), .B(KEYINPUT42), .S(new_n650), .Z(G1325gat));
  NAND2_X1  g450(.A1(new_n275), .A2(new_n276), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n279), .A2(KEYINPUT36), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(G15gat), .B1(new_n642), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n474), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(G15gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n642), .B2(new_n657), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n451), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  NOR3_X1   g460(.A1(new_n582), .A2(new_n616), .A3(new_n640), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n549), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n494), .A3(new_n470), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n448), .A2(new_n451), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n462), .A2(new_n463), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT38), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n470), .A2(new_n668), .A3(new_n457), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n666), .A2(new_n669), .B1(new_n428), .B2(new_n392), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n654), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT101), .B1(new_n280), .B2(new_n466), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n469), .A2(KEYINPUT35), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n473), .A2(new_n474), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n672), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT102), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n672), .A2(new_n673), .A3(new_n679), .A4(new_n676), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n616), .A2(KEYINPUT44), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT44), .B1(new_n476), .B2(new_n616), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n640), .B(KEYINPUT100), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n547), .A2(new_n582), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G29gat), .B1(new_n688), .B2(new_n353), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n665), .A2(new_n689), .ZN(G1328gat));
  NAND3_X1  g489(.A1(new_n663), .A2(new_n495), .A3(new_n430), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT46), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n430), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n688), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(KEYINPUT104), .ZN(new_n697));
  OAI21_X1  g496(.A(G36gat), .B1(new_n696), .B2(KEYINPUT104), .ZN(new_n698));
  OAI221_X1 g497(.A(new_n694), .B1(KEYINPUT46), .B2(new_n691), .C1(new_n697), .C2(new_n698), .ZN(G1329gat));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  INV_X1    g499(.A(G43gat), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n663), .A2(new_n701), .A3(new_n474), .ZN(new_n702));
  INV_X1    g501(.A(new_n688), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n703), .B2(new_n280), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n700), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n280), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT105), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n701), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n702), .A2(new_n700), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(G1330gat));
  NAND3_X1  g509(.A1(new_n703), .A2(G50gat), .A3(new_n428), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n663), .A2(new_n428), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(G50gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g513(.A1(new_n678), .A2(new_n680), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n617), .A2(new_n546), .A3(new_n685), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n353), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT106), .B(G57gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1332gat));
  INV_X1    g519(.A(new_n717), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n695), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT107), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n724), .B(new_n725), .Z(G1333gat));
  NOR2_X1   g525(.A1(new_n717), .A2(new_n656), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(G71gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n721), .A2(G71gat), .A3(new_n280), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(KEYINPUT108), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(KEYINPUT108), .B2(new_n729), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n721), .A2(new_n428), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g533(.A1(new_n582), .A2(new_n546), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n640), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n682), .B2(new_n683), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n353), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n735), .B(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n475), .B1(new_n467), .B2(new_n671), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n616), .B1(new_n743), .B2(new_n673), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n742), .B1(new_n744), .B2(KEYINPUT110), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n614), .A2(new_n615), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT110), .B1(new_n677), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT51), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n677), .A2(KEYINPUT110), .A3(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n736), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n751), .A2(new_n752), .A3(new_n747), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n470), .A2(new_n590), .A3(new_n640), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n740), .B1(new_n754), .B2(new_n755), .ZN(G1336gat));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n685), .A2(G92gat), .A3(new_n695), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n749), .B2(new_n753), .ZN(new_n759));
  INV_X1    g558(.A(new_n737), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n684), .A2(new_n430), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n757), .B1(new_n763), .B2(KEYINPUT52), .ZN(new_n764));
  INV_X1    g563(.A(new_n758), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n752), .B1(new_n751), .B2(new_n747), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n736), .A4(new_n750), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n591), .B1(new_n738), .B2(new_n430), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n757), .B(KEYINPUT52), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n764), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n759), .A2(new_n762), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n759), .A2(new_n762), .A3(KEYINPUT112), .A4(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT113), .B1(new_n772), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT52), .B1(new_n768), .B2(new_n769), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT111), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n770), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n782), .A2(new_n783), .A3(new_n776), .A4(new_n777), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n784), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n739), .B2(new_n654), .ZN(new_n786));
  INV_X1    g585(.A(new_n640), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n656), .A2(G99gat), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n754), .B2(new_n788), .ZN(G1338gat));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  OAI21_X1  g589(.A(G106gat), .B1(new_n739), .B2(new_n451), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n685), .A2(G106gat), .A3(new_n451), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n791), .B1(new_n754), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n793), .B(new_n795), .ZN(G1339gat));
  XOR2_X1   g595(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n621), .B1(new_n637), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n628), .A2(new_n629), .A3(new_n636), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(KEYINPUT54), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n631), .B2(new_n634), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n802), .B(KEYINPUT115), .C1(new_n631), .C2(new_n634), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n635), .B1(new_n807), .B2(KEYINPUT55), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  AOI211_X1 g608(.A(new_n809), .B(new_n800), .C1(new_n805), .C2(new_n806), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT117), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n805), .A2(new_n806), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n799), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n809), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n807), .A2(KEYINPUT55), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n635), .A4(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n530), .B1(new_n527), .B2(new_n528), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(KEYINPUT118), .B(new_n530), .C1(new_n527), .C2(new_n528), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n537), .A2(new_n539), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n481), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n746), .A2(new_n826), .A3(new_n545), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n818), .A2(new_n828), .A3(KEYINPUT119), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n811), .A2(new_n817), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n827), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n545), .A2(new_n826), .A3(new_n640), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n831), .B2(new_n547), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n616), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n582), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n617), .A2(new_n546), .A3(new_n640), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n839), .A2(new_n353), .A3(new_n430), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n279), .A2(new_n451), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n547), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n656), .A2(new_n428), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n546), .A2(G113gat), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n844), .A2(G113gat), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT120), .ZN(G1340gat));
  INV_X1    g648(.A(G120gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n846), .A2(new_n850), .A3(new_n685), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n840), .A2(new_n842), .A3(new_n640), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(G1341gat));
  INV_X1    g652(.A(new_n582), .ZN(new_n854));
  OAI21_X1  g653(.A(G127gat), .B1(new_n846), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n854), .A2(G127gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n843), .B2(new_n856), .ZN(G1342gat));
  NOR3_X1   g656(.A1(new_n616), .A2(new_n841), .A3(G134gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT56), .Z(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n846), .B2(new_n616), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1343gat));
  AOI21_X1  g661(.A(KEYINPUT119), .B1(new_n818), .B2(new_n828), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n831), .A2(new_n827), .A3(new_n830), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n814), .A2(new_n635), .A3(new_n816), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n865), .B1(new_n542), .B2(new_n545), .ZN(new_n866));
  INV_X1    g665(.A(new_n834), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n863), .A2(new_n864), .B1(new_n868), .B2(new_n746), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n838), .B1(new_n869), .B2(new_n854), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT57), .B1(new_n870), .B2(new_n451), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n872), .B(new_n428), .C1(new_n837), .C2(new_n838), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n280), .A2(new_n353), .A3(new_n430), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n871), .A2(new_n546), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G141gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT121), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT58), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n280), .A2(new_n451), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n840), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n547), .A2(G141gat), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n882), .A2(new_n883), .B1(G141gat), .B2(new_n875), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n875), .B2(G141gat), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT122), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n879), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n884), .B1(new_n879), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(G1344gat));
  OR3_X1    g690(.A1(new_n881), .A2(G148gat), .A3(new_n787), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT123), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n838), .B(KEYINPUT124), .Z(new_n895));
  NOR2_X1   g694(.A1(new_n868), .A2(new_n746), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n827), .A2(new_n865), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n854), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT125), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n895), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n900), .A2(new_n872), .A3(new_n428), .A4(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT57), .B1(new_n839), .B2(new_n451), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n640), .A3(new_n874), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n894), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n894), .A2(G148gat), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n640), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n893), .B1(new_n907), .B2(new_n910), .ZN(G1345gat));
  NAND3_X1  g710(.A1(new_n882), .A2(new_n284), .A3(new_n582), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n909), .A2(new_n582), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n284), .ZN(G1346gat));
  NAND3_X1  g713(.A1(new_n882), .A2(new_n285), .A3(new_n746), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n909), .A2(new_n746), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n285), .ZN(G1347gat));
  OR2_X1    g716(.A1(new_n837), .A2(new_n838), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(KEYINPUT126), .A3(new_n353), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n839), .B2(new_n470), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n695), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n842), .A3(new_n546), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n470), .A2(new_n695), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n845), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n918), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n547), .A2(new_n210), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n923), .A2(new_n210), .B1(new_n926), .B2(new_n927), .ZN(G1348gat));
  INV_X1    g727(.A(new_n926), .ZN(new_n929));
  OAI21_X1  g728(.A(G176gat), .B1(new_n929), .B2(new_n685), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n922), .A2(new_n842), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n640), .A2(new_n211), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(G1349gat));
  NAND2_X1  g732(.A1(new_n926), .A2(new_n582), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT127), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n926), .A2(new_n936), .A3(new_n582), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(G183gat), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n582), .A2(new_n246), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n931), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n938), .B(new_n942), .C1(new_n931), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1350gat));
  AOI21_X1  g743(.A(new_n213), .B1(new_n926), .B2(new_n746), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT61), .Z(new_n946));
  NAND2_X1  g745(.A1(new_n746), .A2(new_n213), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n931), .B2(new_n947), .ZN(G1351gat));
  NAND2_X1  g747(.A1(new_n654), .A2(new_n924), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n905), .A2(G197gat), .A3(new_n546), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n922), .A2(new_n880), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n480), .B1(new_n952), .B2(new_n547), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n951), .A2(new_n953), .ZN(G1352gat));
  NAND3_X1  g753(.A1(new_n905), .A2(new_n686), .A3(new_n950), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G204gat), .ZN(new_n956));
  INV_X1    g755(.A(new_n952), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n787), .A2(G204gat), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n957), .A2(KEYINPUT62), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT62), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1353gat));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n360), .A3(new_n582), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n903), .A2(new_n582), .A3(new_n904), .A4(new_n950), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1354gat));
  NAND3_X1  g765(.A1(new_n957), .A2(new_n361), .A3(new_n746), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n905), .A2(new_n746), .A3(new_n950), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n361), .ZN(G1355gat));
endmodule


