//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AND2_X1   g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n202), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n211), .B(new_n215), .C1(G87), .C2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G50), .A2(G226), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(G68), .A2(G238), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n207), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n210), .B(new_n226), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT73), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT73), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n214), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n222), .A2(G1698), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n252), .A2(new_n254), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n253), .A2(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT65), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT65), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n254), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G303), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n258), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n227), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(new_n248), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT5), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n272), .A2(new_n274), .A3(new_n275), .A4(G45), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n276), .A2(new_n270), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n267), .A2(new_n271), .B1(G270), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  OR2_X1    g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G116), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n227), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(G1), .B2(new_n248), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G283), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n291), .B(new_n228), .C1(G33), .C2(new_n213), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n292), .B(new_n288), .C1(new_n228), .C2(G116), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT20), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n294), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n286), .B1(new_n290), .B2(new_n285), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n281), .A2(G169), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT21), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n281), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G179), .A3(new_n297), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n281), .A2(KEYINPUT21), .A3(G169), .A4(new_n297), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT73), .B(G33), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n305), .A2(G20), .A3(new_n285), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n228), .A2(G107), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT23), .ZN(new_n309));
  INV_X1    g0109(.A(G87), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(G20), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n261), .B2(new_n264), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n307), .B(new_n309), .C1(new_n313), .C2(KEYINPUT22), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n252), .A2(new_n254), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT22), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n315), .A2(new_n316), .A3(new_n312), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT86), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n254), .A2(new_n262), .A3(new_n263), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n263), .B1(new_n254), .B2(new_n262), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n311), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n306), .B1(new_n321), .B2(new_n316), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT86), .ZN(new_n323));
  INV_X1    g0123(.A(new_n315), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT22), .A3(new_n311), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n322), .A2(new_n323), .A3(new_n325), .A4(new_n309), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n318), .A2(KEYINPUT24), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT24), .ZN(new_n328));
  OAI211_X1 g0128(.A(KEYINPUT86), .B(new_n328), .C1(new_n314), .C2(new_n317), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n288), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n290), .B(KEYINPUT81), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G107), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n284), .A2(new_n221), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n333), .B(KEYINPUT25), .Z(new_n334));
  NAND3_X1  g0134(.A1(new_n330), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  OR2_X1    g0135(.A1(G250), .A2(G1698), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n214), .A2(G1698), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n252), .A2(new_n254), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n305), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G294), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n271), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT87), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n342), .A2(new_n343), .B1(G264), .B2(new_n277), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(KEYINPUT87), .A3(new_n271), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n280), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G169), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n277), .A2(G264), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n342), .A2(new_n280), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n335), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT88), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT88), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n335), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n304), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n279), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n220), .B(new_n255), .C1(new_n261), .C2(new_n264), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT71), .ZN(new_n362));
  AOI21_X1  g0162(.A(G1698), .B1(new_n261), .B2(new_n264), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(new_n363), .B2(G226), .ZN(new_n364));
  OAI211_X1 g0164(.A(G226), .B(new_n255), .C1(new_n319), .C2(new_n320), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(KEYINPUT71), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n359), .B(new_n361), .C1(new_n364), .C2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n358), .B1(new_n367), .B2(new_n271), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n270), .A2(new_n357), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT64), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G238), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n368), .B2(new_n372), .ZN(new_n374));
  OAI21_X1  g0174(.A(G200), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n228), .A2(G33), .ZN(new_n376));
  XOR2_X1   g0176(.A(new_n376), .B(KEYINPUT67), .Z(new_n377));
  INV_X1    g0177(.A(G68), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n377), .A2(G77), .B1(G20), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G50), .ZN(new_n380));
  NOR2_X1   g0180(.A1(G20), .A2(G33), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n379), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n288), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT11), .ZN(new_n385));
  INV_X1    g0185(.A(new_n284), .ZN(new_n386));
  OR3_X1    g0186(.A1(new_n386), .A2(KEYINPUT12), .A3(G68), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT12), .B1(new_n386), .B2(G68), .ZN(new_n388));
  INV_X1    g0188(.A(new_n282), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(new_n288), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n387), .A2(new_n388), .B1(G68), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n358), .ZN(new_n394));
  INV_X1    g0194(.A(new_n359), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n363), .A2(new_n362), .A3(G226), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n365), .A2(KEYINPUT71), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n395), .B(new_n360), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n372), .B(new_n394), .C1(new_n398), .C2(new_n270), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(G190), .A3(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n375), .A2(new_n393), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n265), .A2(G238), .A3(G1698), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n221), .B2(new_n265), .ZN(new_n406));
  INV_X1    g0206(.A(new_n265), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n407), .A2(new_n220), .A3(G1698), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n271), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n371), .A2(G244), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n394), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G200), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G20), .A2(G77), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT15), .B(G87), .Z(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  OR2_X1    g0215(.A1(KEYINPUT8), .A2(G58), .ZN(new_n416));
  NAND2_X1  g0216(.A1(KEYINPUT8), .A2(G58), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n413), .B1(new_n415), .B2(new_n376), .C1(new_n382), .C2(new_n418), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n288), .B1(G77), .B2(new_n390), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n284), .A2(new_n202), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G190), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n412), .B(new_n423), .C1(new_n424), .C2(new_n411), .ZN(new_n425));
  INV_X1    g0225(.A(G169), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n411), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n409), .A2(new_n348), .A3(new_n394), .A4(new_n410), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n422), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n400), .A2(new_n401), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n432), .A2(G169), .B1(KEYINPUT72), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n435));
  AOI211_X1 g0235(.A(new_n426), .B(new_n435), .C1(new_n400), .C2(new_n401), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n400), .A2(G179), .A3(new_n401), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n434), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n404), .B(new_n431), .C1(new_n441), .C2(new_n393), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT66), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n418), .B(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT75), .A3(new_n282), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n418), .A2(new_n443), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT66), .B1(new_n416), .B2(new_n417), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n282), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT75), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n445), .A2(new_n450), .A3(new_n289), .ZN(new_n451));
  INV_X1    g0251(.A(new_n444), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n284), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n261), .A2(new_n228), .A3(new_n264), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT7), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n262), .B1(new_n305), .B2(KEYINPUT3), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G68), .ZN(new_n462));
  XNOR2_X1  g0262(.A(G58), .B(G68), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n463), .A2(G20), .B1(G159), .B2(new_n381), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n455), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(G20), .B1(new_n252), .B2(new_n254), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n457), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(G68), .B1(new_n466), .B2(new_n457), .ZN(new_n469));
  OAI211_X1 g0269(.A(KEYINPUT16), .B(new_n464), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n288), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n454), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G223), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n255), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n255), .A2(G226), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n252), .A2(new_n254), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G87), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n271), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT76), .ZN(new_n480));
  INV_X1    g0280(.A(new_n370), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n358), .B1(new_n481), .B2(G232), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT76), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(new_n483), .A3(new_n271), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n480), .A2(new_n348), .A3(new_n482), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n479), .A2(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n426), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n472), .A2(KEYINPUT18), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT77), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT18), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n451), .A2(new_n453), .ZN(new_n492));
  INV_X1    g0292(.A(new_n288), .ZN(new_n493));
  INV_X1    g0293(.A(new_n464), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n315), .A2(new_n228), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n378), .B1(new_n495), .B2(KEYINPUT7), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n496), .B2(new_n467), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n493), .B1(new_n497), .B2(KEYINPUT16), .ZN(new_n498));
  INV_X1    g0298(.A(new_n455), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n378), .B1(new_n458), .B2(new_n460), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n494), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n492), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n485), .A2(new_n487), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n491), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT77), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n472), .A2(new_n488), .A3(new_n505), .A4(KEYINPUT18), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n490), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n501), .A2(new_n288), .A3(new_n470), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n480), .A2(new_n424), .A3(new_n482), .A4(new_n484), .ZN(new_n509));
  INV_X1    g0309(.A(G200), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n486), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n508), .A2(new_n512), .A3(new_n454), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT78), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT17), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n502), .A2(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(new_n516), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n507), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT79), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n371), .A2(G226), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n473), .A2(G1698), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(G222), .B2(G1698), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n270), .B1(new_n265), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(G77), .B2(new_n265), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n522), .A2(new_n526), .A3(new_n348), .A4(new_n394), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT69), .ZN(new_n528));
  XNOR2_X1  g0328(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n390), .A2(G50), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n201), .A2(new_n228), .ZN(new_n531));
  INV_X1    g0331(.A(G150), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n382), .A2(new_n532), .ZN(new_n533));
  AOI211_X1 g0333(.A(new_n531), .B(new_n533), .C1(new_n444), .C2(new_n377), .ZN(new_n534));
  OAI221_X1 g0334(.A(new_n530), .B1(G50), .B2(new_n386), .C1(new_n534), .C2(new_n493), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n522), .A2(new_n394), .A3(new_n526), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n426), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT68), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n537), .A3(KEYINPUT68), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n529), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n535), .A2(KEYINPUT9), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n386), .A2(G50), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n533), .B1(new_n444), .B2(new_n377), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n228), .B2(new_n201), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n544), .B1(new_n546), .B2(new_n288), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT9), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(new_n530), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n536), .A2(G200), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT70), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT70), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n536), .A2(new_n553), .A3(G200), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n554), .C1(new_n424), .C2(new_n536), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT10), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n554), .B1(new_n424), .B2(new_n536), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n543), .A2(new_n549), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT10), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .A4(new_n552), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n542), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT79), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n507), .A2(new_n519), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n521), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n442), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n301), .A2(G190), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n297), .B1(new_n281), .B2(G200), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT85), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G238), .A2(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n212), .B2(G1698), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(new_n252), .A3(new_n254), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n339), .A2(G116), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n270), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(G45), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n270), .B(G250), .C1(G1), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n577), .A2(new_n279), .A3(G1), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n348), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G169), .B2(new_n581), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT84), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n252), .A2(new_n228), .A3(G68), .A4(new_n254), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n228), .B1(new_n359), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G87), .B2(new_n205), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n587), .B1(new_n376), .B2(new_n213), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n288), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n386), .A2(new_n414), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n592), .A2(KEYINPUT82), .A3(new_n594), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n414), .B(KEYINPUT83), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n288), .B(new_n284), .C1(new_n275), .C2(G33), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT81), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n290), .A2(KEYINPUT81), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n585), .B1(new_n599), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT82), .B1(new_n592), .B2(new_n594), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n596), .B(new_n593), .C1(new_n591), .C2(new_n288), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n606), .B(new_n585), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n584), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n290), .B(new_n603), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n608), .A2(new_n609), .B1(new_n613), .B2(new_n310), .ZN(new_n614));
  OR3_X1    g0414(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n424), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n581), .A2(new_n510), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n461), .A2(G107), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n382), .A2(new_n202), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT80), .ZN(new_n624));
  NAND2_X1  g0424(.A1(KEYINPUT6), .A2(G97), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n624), .B1(new_n625), .B2(G107), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n221), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(G97), .ZN(new_n627));
  XOR2_X1   g0427(.A(G97), .B(G107), .Z(new_n628));
  OAI211_X1 g0428(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(KEYINPUT6), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G20), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n621), .A2(new_n623), .A3(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n288), .B1(G97), .B2(new_n331), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n252), .A2(G244), .A3(new_n255), .A4(new_n254), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT4), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(KEYINPUT4), .B(new_n255), .C1(new_n319), .C2(new_n320), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(new_n212), .ZN(new_n637));
  OAI211_X1 g0437(.A(G250), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n291), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n271), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n277), .A2(G257), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n280), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G200), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n284), .A2(new_n213), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n640), .A2(G190), .A3(new_n280), .A4(new_n641), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n632), .A2(new_n643), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n331), .A2(G97), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n221), .B1(new_n458), .B2(new_n460), .ZN(new_n648));
  INV_X1    g0448(.A(new_n630), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n648), .A2(new_n622), .A3(new_n649), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n647), .B(new_n644), .C1(new_n650), .C2(new_n493), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n642), .A2(new_n426), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n640), .A2(new_n348), .A3(new_n280), .A4(new_n641), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n646), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n350), .ZN(new_n656));
  OAI22_X1  g0456(.A1(new_n346), .A2(G190), .B1(G200), .B2(new_n656), .ZN(new_n657));
  AND4_X1   g0457(.A1(new_n332), .A2(new_n657), .A3(new_n330), .A4(new_n334), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n620), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n356), .A2(new_n566), .A3(new_n571), .A4(new_n659), .ZN(G372));
  NAND2_X1  g0460(.A1(new_n556), .A2(new_n561), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT89), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n429), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n427), .A2(KEYINPUT89), .A3(new_n422), .A4(new_n428), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(G169), .B1(new_n373), .B2(new_n374), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n435), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n432), .A2(KEYINPUT72), .A3(new_n433), .A4(G169), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n437), .A4(new_n439), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n665), .B1(new_n669), .B2(new_n392), .ZN(new_n670));
  INV_X1    g0470(.A(new_n517), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n514), .A2(new_n515), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n516), .B1(new_n513), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n670), .A2(new_n403), .A3(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n504), .A2(new_n489), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n661), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n542), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n566), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT84), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n610), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n618), .B1(new_n683), .B2(new_n584), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT26), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n583), .B1(new_n682), .B2(new_n610), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT26), .ZN(new_n688));
  NOR4_X1   g0488(.A1(new_n687), .A2(new_n654), .A3(new_n618), .A4(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n612), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n612), .A2(new_n654), .A3(new_n619), .A4(new_n646), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n304), .B1(new_n351), .B2(new_n335), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n691), .A2(new_n692), .A3(new_n658), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n679), .B1(new_n680), .B2(new_n694), .ZN(G369));
  INV_X1    g0495(.A(new_n304), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n571), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n283), .A2(G20), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n275), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G213), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G343), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n297), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n304), .A2(new_n705), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G330), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  INV_X1    g0511(.A(new_n704), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n352), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT92), .Z(new_n714));
  NAND2_X1  g0514(.A1(new_n353), .A2(new_n355), .ZN(new_n715));
  INV_X1    g0515(.A(new_n658), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n335), .A2(new_n704), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n715), .B(new_n716), .C1(KEYINPUT91), .C2(new_n717), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n717), .A2(KEYINPUT91), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n714), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n711), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n352), .A2(new_n704), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n696), .A2(new_n704), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT93), .Z(G399));
  INV_X1    g0526(.A(new_n208), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(G1), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(new_n230), .B2(new_n729), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n335), .A2(new_n351), .A3(new_n354), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n354), .B1(new_n335), .B2(new_n351), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n696), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n659), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n687), .B1(new_n686), .B2(KEYINPUT95), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n612), .A2(new_n685), .A3(new_n619), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n688), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT95), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n684), .A2(KEYINPUT26), .A3(new_n685), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n737), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(KEYINPUT29), .A3(new_n712), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n712), .B1(new_n690), .B2(new_n693), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT29), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n356), .A2(new_n659), .A3(new_n571), .A4(new_n712), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n281), .A2(new_n615), .A3(new_n348), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n640), .A2(new_n641), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n750), .A2(KEYINPUT30), .A3(new_n656), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n656), .A2(new_n581), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(new_n642), .A3(new_n348), .A4(new_n281), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n750), .A2(new_n656), .A3(new_n751), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT30), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n752), .B(new_n754), .C1(new_n757), .C2(KEYINPUT94), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n757), .A2(KEYINPUT94), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n704), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n757), .A2(new_n752), .A3(new_n754), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n749), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n745), .A2(new_n748), .B1(G330), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n733), .B1(new_n766), .B2(G1), .ZN(G364));
  AOI21_X1  g0567(.A(new_n711), .B1(new_n709), .B2(new_n708), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n698), .A2(G45), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT96), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(KEYINPUT96), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(G1), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n729), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT97), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n768), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n775), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT98), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  OR2_X1    g0580(.A1(KEYINPUT99), .A2(G169), .ZN(new_n781));
  NAND2_X1  g0581(.A1(KEYINPUT99), .A2(G169), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n781), .A2(G20), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n268), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT100), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n780), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n324), .A2(new_n727), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n231), .A2(new_n577), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n789), .C1(new_n246), .C2(new_n577), .ZN(new_n790));
  INV_X1    g0590(.A(G355), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n265), .A2(new_n208), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n790), .B1(G116), .B2(new_n208), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n708), .A2(new_n780), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n228), .A2(new_n348), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n795), .A2(G190), .A3(new_n510), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n424), .A2(new_n510), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n797), .A2(G58), .B1(new_n800), .B2(G50), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n228), .A2(G179), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G190), .A2(G200), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  OAI21_X1  g0605(.A(KEYINPUT32), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n424), .A2(G179), .A3(G200), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n228), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n801), .B(new_n806), .C1(new_n213), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n510), .A2(G190), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n802), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT101), .Z(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G107), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n795), .A2(new_n803), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n407), .B1(G77), .B2(new_n816), .ZN(new_n817));
  OR3_X1    g0617(.A1(new_n804), .A2(KEYINPUT32), .A3(new_n805), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n798), .A2(new_n802), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G87), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n814), .A2(new_n817), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n795), .A2(new_n810), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n809), .B(new_n822), .C1(G68), .C2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n813), .A2(G283), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G326), .A2(new_n800), .B1(new_n816), .B2(G311), .ZN(new_n827));
  INV_X1    g0627(.A(G322), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT102), .B(KEYINPUT33), .ZN(new_n829));
  INV_X1    g0629(.A(G317), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n829), .B(new_n830), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n827), .B1(new_n828), .B2(new_n796), .C1(new_n831), .C2(new_n823), .ZN(new_n832));
  INV_X1    g0632(.A(G294), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n808), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n804), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(G329), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n407), .B(new_n836), .C1(new_n266), .C2(new_n819), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n826), .A2(new_n832), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n786), .B1(new_n825), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n777), .B1(new_n794), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n776), .A2(new_n840), .ZN(G396));
  NOR2_X1   g0641(.A1(new_n423), .A2(new_n712), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n430), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n663), .A2(new_n664), .A3(new_n842), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n712), .B(new_n847), .C1(new_n690), .C2(new_n693), .ZN(new_n848));
  INV_X1    g0648(.A(new_n746), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n846), .B(KEYINPUT106), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n765), .A2(G330), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT107), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n775), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(KEYINPUT107), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n779), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n786), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT103), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n777), .B1(new_n860), .B2(new_n202), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n813), .A2(G87), .ZN(new_n862));
  XOR2_X1   g0662(.A(KEYINPUT104), .B(G283), .Z(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n862), .B1(new_n833), .B2(new_n796), .C1(new_n823), .C2(new_n864), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n808), .A2(new_n213), .B1(new_n815), .B2(new_n285), .ZN(new_n866));
  INV_X1    g0666(.A(G311), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n407), .B1(new_n221), .B2(new_n819), .C1(new_n867), .C2(new_n804), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n266), .B2(new_n799), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n812), .A2(new_n378), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G50), .B2(new_n820), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n808), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n873), .A2(KEYINPUT105), .B1(G58), .B2(new_n874), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n797), .A2(G143), .B1(new_n824), .B2(G150), .ZN(new_n876));
  INV_X1    g0676(.A(G137), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n876), .B1(new_n877), .B2(new_n799), .C1(new_n805), .C2(new_n815), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT34), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n835), .A2(G132), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT105), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n315), .B1(new_n872), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n875), .A2(new_n879), .A3(new_n880), .A4(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n870), .A2(new_n883), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n861), .B1(new_n785), .B2(new_n884), .C1(new_n847), .C2(new_n779), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n857), .A2(new_n885), .ZN(G384));
  INV_X1    g0686(.A(KEYINPUT40), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n393), .A2(new_n712), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n404), .B(new_n889), .C1(new_n441), .C2(new_n393), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n669), .A2(new_n392), .A3(new_n704), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n846), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n497), .A2(new_n455), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n454), .B1(new_n895), .B2(new_n471), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n502), .A2(new_n512), .B1(new_n896), .B2(new_n488), .ZN(new_n897));
  INV_X1    g0697(.A(new_n702), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n894), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n503), .B1(new_n508), .B2(new_n454), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n508), .A2(new_n512), .A3(new_n454), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT109), .B1(new_n502), .B2(new_n702), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT109), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n472), .A2(new_n904), .A3(new_n898), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(KEYINPUT110), .B(KEYINPUT37), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n900), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n899), .B1(new_n507), .B2(new_n519), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n893), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n899), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n520), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n897), .A2(new_n899), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n915));
  INV_X1    g0715(.A(new_n901), .ZN(new_n916));
  INV_X1    g0716(.A(new_n905), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n904), .B1(new_n472), .B2(new_n898), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n513), .B(new_n916), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n915), .B1(new_n919), .B2(new_n907), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n913), .A2(new_n920), .A3(KEYINPUT38), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n911), .A2(KEYINPUT111), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT111), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n913), .A2(new_n920), .A3(new_n923), .A4(KEYINPUT38), .ZN(new_n924));
  OAI211_X1 g0724(.A(KEYINPUT31), .B(new_n704), .C1(new_n758), .C2(new_n759), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n749), .A2(new_n762), .A3(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n892), .A2(new_n922), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n888), .B(new_n403), .C1(new_n669), .C2(new_n392), .ZN(new_n928));
  INV_X1    g0728(.A(new_n891), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n926), .B(new_n847), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT113), .B1(new_n917), .B2(new_n918), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n907), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n919), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n905), .B(new_n903), .C1(new_n674), .C2(new_n676), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n906), .A2(new_n907), .A3(new_n932), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n893), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n887), .B1(new_n938), .B2(new_n921), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n887), .A2(new_n927), .B1(new_n931), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT114), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n566), .A2(new_n926), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(G330), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n745), .A2(new_n566), .A3(new_n748), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n679), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n669), .A2(new_n392), .A3(new_n712), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT112), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT112), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n669), .A2(new_n950), .A3(new_n392), .A4(new_n712), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n924), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT39), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n938), .A2(new_n955), .A3(new_n921), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n953), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n429), .A2(new_n704), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n848), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n890), .A2(new_n891), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n960), .A2(new_n922), .A3(new_n924), .A4(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n676), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n898), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n957), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n947), .B(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n275), .B2(new_n698), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n285), .B1(new_n629), .B2(KEYINPUT35), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n970), .B(new_n229), .C1(KEYINPUT35), .C2(new_n629), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT36), .ZN(new_n972));
  OAI21_X1  g0772(.A(G77), .B1(new_n219), .B2(new_n378), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n973), .A2(new_n230), .B1(G50), .B2(new_n378), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(G1), .A3(new_n283), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT108), .Z(new_n976));
  NAND3_X1  g0776(.A1(new_n969), .A2(new_n972), .A3(new_n976), .ZN(G367));
  NAND2_X1  g0777(.A1(new_n720), .A2(new_n723), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n685), .A2(new_n704), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n651), .A2(new_n704), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n646), .A2(new_n654), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n978), .A2(KEYINPUT42), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n654), .B1(new_n715), .B2(new_n981), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n712), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT42), .B1(new_n978), .B2(new_n983), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n614), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n684), .B1(new_n989), .B2(new_n712), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n687), .A2(new_n614), .A3(new_n704), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT115), .Z(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n988), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n995), .B1(new_n988), .B2(new_n996), .ZN(new_n998));
  OR4_X1    g0798(.A1(new_n721), .A2(new_n997), .A3(new_n998), .A4(new_n983), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n997), .A2(new_n998), .B1(new_n721), .B2(new_n983), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n728), .B(KEYINPUT41), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n724), .A2(new_n982), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT45), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT44), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n724), .A2(new_n1006), .A3(new_n982), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1006), .B1(new_n724), .B2(new_n982), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(KEYINPUT116), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT116), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1010), .B(new_n1006), .C1(new_n724), .C2(new_n982), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1005), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n721), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n720), .B(new_n723), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(new_n711), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n766), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1005), .A2(new_n1009), .A3(new_n721), .A4(new_n1011), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1014), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1002), .B1(new_n1020), .B2(new_n766), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n999), .B(new_n1000), .C1(new_n1021), .C2(new_n772), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n992), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n777), .B1(new_n1023), .B2(new_n780), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n788), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n787), .B1(new_n208), .B2(new_n415), .C1(new_n239), .C2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n808), .A2(new_n378), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n796), .A2(new_n532), .B1(new_n811), .B2(new_n202), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G58), .C2(new_n820), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n824), .A2(G159), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n407), .B1(G137), .B2(new_n835), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G143), .A2(new_n800), .B1(new_n816), .B2(G50), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n820), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT46), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n819), .B2(new_n285), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(new_n830), .C2(new_n804), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n324), .B(new_n1037), .C1(G294), .C2(new_n824), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n797), .A2(G303), .B1(new_n800), .B2(G311), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n864), .A2(new_n815), .B1(new_n808), .B2(new_n221), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT117), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n811), .A2(new_n213), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1033), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT47), .Z(new_n1045));
  OAI211_X1 g0845(.A(new_n1024), .B(new_n1026), .C1(new_n785), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1022), .A2(new_n1046), .ZN(G387));
  OAI211_X1 g0847(.A(new_n714), .B(new_n780), .C1(new_n719), .C2(new_n718), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n797), .A2(G317), .B1(new_n824), .B2(G311), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n266), .B2(new_n815), .C1(new_n828), .C2(new_n799), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT48), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n833), .B2(new_n819), .C1(new_n808), .C2(new_n864), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n324), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n835), .A2(G326), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n811), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(G116), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n600), .A2(new_n808), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n444), .B2(new_n824), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n378), .B2(new_n815), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G159), .B2(new_n800), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n813), .A2(G97), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n819), .A2(new_n202), .B1(new_n804), .B2(new_n532), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G50), .B2(new_n797), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n324), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n785), .B1(new_n1059), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n788), .B1(new_n236), .B2(new_n577), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n730), .B2(new_n792), .ZN(new_n1070));
  OR3_X1    g0870(.A1(new_n418), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT50), .B1(new_n418), .B2(G50), .ZN(new_n1072));
  AOI21_X1  g0872(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n730), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n727), .A2(new_n221), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n777), .B(new_n1068), .C1(new_n787), .C2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1016), .A2(new_n772), .B1(new_n1048), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n728), .B1(new_n1016), .B2(new_n766), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1018), .B2(new_n1080), .ZN(G393));
  AOI21_X1  g0881(.A(new_n777), .B1(new_n983), .B2(new_n780), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n787), .B1(new_n213), .B2(new_n208), .C1(new_n243), .C2(new_n1025), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n816), .A2(G294), .B1(new_n820), .B2(new_n863), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1084), .B(new_n407), .C1(new_n266), .C2(new_n823), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n796), .A2(new_n867), .B1(new_n799), .B2(new_n830), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n814), .B(new_n1087), .C1(new_n285), .C2(new_n808), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1085), .B(new_n1088), .C1(G322), .C2(new_n835), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G50), .A2(new_n824), .B1(new_n835), .B2(G143), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n418), .B2(new_n815), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n796), .A2(new_n805), .B1(new_n799), .B2(new_n532), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT51), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1092), .A2(new_n1093), .B1(G77), .B2(new_n874), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n862), .A2(new_n324), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1091), .B(new_n1096), .C1(G68), .C2(new_n820), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1089), .A2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT118), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1082), .B(new_n1083), .C1(new_n785), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n773), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n729), .B1(new_n1101), .B2(new_n1017), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1020), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(G390));
  NAND3_X1  g0905(.A1(new_n566), .A2(G330), .A3(new_n926), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n677), .A2(new_n945), .A3(new_n1106), .A4(new_n678), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n765), .A2(G330), .A3(new_n847), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n403), .B1(new_n669), .B2(new_n392), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n441), .A2(new_n393), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1109), .A2(new_n889), .B1(new_n1110), .B2(new_n704), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n961), .A2(G330), .A3(new_n847), .A4(new_n926), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n960), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n926), .A2(new_n850), .A3(G330), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1111), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n744), .A2(new_n712), .A3(new_n847), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(new_n959), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n892), .A2(G330), .A3(new_n765), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1107), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n952), .B1(new_n921), .B2(new_n938), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1119), .B2(new_n1111), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n848), .A2(new_n959), .B1(new_n890), .B2(new_n891), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n954), .B(new_n956), .C1(new_n952), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1120), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1113), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1122), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  AND4_X1   g0931(.A1(new_n678), .A2(new_n677), .A3(new_n945), .A4(new_n1106), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1112), .A2(new_n1113), .B1(new_n848), .B2(new_n959), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n954), .A2(new_n956), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1125), .A2(new_n952), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1111), .B1(new_n959), .B2(new_n1118), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n938), .A2(new_n921), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n953), .A2(new_n1139), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1136), .A2(new_n1137), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1113), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1135), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1131), .A2(new_n1144), .A3(new_n728), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n954), .A2(new_n858), .A3(new_n956), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n800), .A2(G283), .B1(new_n835), .B2(G294), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n213), .B2(new_n815), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1149), .B(new_n871), .C1(G77), .C2(new_n874), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n824), .A2(G107), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n407), .A2(new_n821), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT119), .Z(new_n1153));
  NAND2_X1  g0953(.A1(new_n797), .A2(G116), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(G128), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n799), .A2(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n808), .A2(new_n805), .B1(new_n380), .B2(new_n811), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(G137), .C2(new_n824), .ZN(new_n1159));
  XOR2_X1   g0959(.A(KEYINPUT54), .B(G143), .Z(new_n1160));
  NAND2_X1  g0960(.A1(new_n816), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n819), .A2(new_n532), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT53), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n797), .A2(G132), .B1(new_n835), .B2(G125), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1164), .A2(new_n265), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1159), .A2(new_n1161), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n785), .B1(new_n1155), .B2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n777), .B(new_n1167), .C1(new_n452), .C2(new_n860), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1146), .A2(new_n772), .B1(new_n1147), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1145), .A2(new_n1169), .ZN(G378));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1136), .A2(new_n952), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n922), .A2(new_n924), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n964), .B1(new_n1173), .B2(new_n1125), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n661), .A2(new_n678), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT124), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n535), .A2(new_n898), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n562), .A2(KEYINPUT124), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1178), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT124), .B1(new_n661), .B2(new_n678), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1176), .B(new_n542), .C1(new_n556), .C2(new_n561), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1185));
  AND3_X1   g0985(.A1(new_n1180), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1180), .B2(new_n1184), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1172), .A2(new_n1174), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n922), .A2(new_n924), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n887), .B1(new_n1190), .B2(new_n930), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n939), .A2(new_n926), .A3(new_n892), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1191), .A2(G330), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n957), .B2(new_n966), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1189), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1189), .A2(new_n1195), .B1(G330), .B2(new_n940), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1107), .B1(new_n1146), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1171), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1189), .A2(new_n1195), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1193), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1189), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1207), .A3(KEYINPUT57), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1201), .A2(new_n728), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n777), .B1(new_n1194), .B2(new_n858), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n796), .A2(new_n221), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1027), .B1(G283), .B2(new_n835), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G97), .A2(new_n824), .B1(new_n1057), .B2(G58), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT121), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n315), .B(new_n269), .C1(new_n202), .C2(new_n819), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1212), .B(new_n1213), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1211), .B(new_n1216), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n285), .B2(new_n799), .C1(new_n600), .C2(new_n815), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT58), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n874), .A2(G150), .B1(new_n800), .B2(G125), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT123), .Z(new_n1223));
  NAND2_X1  g1023(.A1(new_n820), .A2(new_n1160), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1224), .A2(KEYINPUT122), .B1(G132), .B2(new_n824), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(new_n1156), .C2(new_n796), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G137), .B2(new_n816), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(KEYINPUT122), .B2(new_n1224), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G159), .A2(new_n1057), .B1(new_n835), .B2(G124), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n248), .A3(new_n269), .A4(new_n1230), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1220), .B(new_n1221), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n250), .A2(KEYINPUT3), .A3(G33), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G50), .B1(new_n1234), .B2(new_n269), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT120), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n786), .B1(new_n1233), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n859), .A2(new_n380), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1210), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1206), .B2(new_n772), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1209), .A2(new_n1240), .ZN(G375));
  NOR2_X1   g1041(.A1(new_n1199), .A2(new_n1132), .ZN(new_n1242));
  OR3_X1    g1042(.A1(new_n1242), .A2(new_n1002), .A3(new_n1122), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1060), .B1(G283), .B2(new_n797), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1244), .B1(new_n221), .B2(new_n815), .C1(new_n285), .C2(new_n823), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n819), .A2(new_n213), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n812), .A2(new_n202), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n407), .B1(new_n833), .B2(new_n799), .C1(new_n266), .C2(new_n804), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n315), .B1(G58), .B2(new_n1057), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT125), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G132), .A2(new_n800), .B1(new_n824), .B2(new_n1160), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1252), .B1(new_n1156), .B2(new_n804), .C1(new_n877), .C2(new_n796), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n808), .A2(new_n380), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n532), .A2(new_n815), .B1(new_n819), .B2(new_n805), .ZN(new_n1255));
  NOR4_X1   g1055(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n786), .B1(new_n1249), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n860), .A2(new_n378), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n775), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1111), .B2(new_n858), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1199), .B2(new_n772), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1243), .A2(new_n1261), .ZN(G381));
  NAND3_X1  g1062(.A1(new_n1022), .A2(new_n1046), .A3(new_n1104), .ZN(new_n1263));
  OR3_X1    g1063(.A1(new_n1263), .A2(G384), .A3(G381), .ZN(new_n1264));
  INV_X1    g1064(.A(G378), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1209), .A2(new_n1265), .A3(new_n1240), .ZN(new_n1266));
  OR3_X1    g1066(.A1(new_n1266), .A2(G396), .A3(G393), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1264), .A2(new_n1267), .ZN(G407));
  OAI211_X1 g1068(.A(G407), .B(G213), .C1(G343), .C2(new_n1266), .ZN(G409));
  XOR2_X1   g1069(.A(G393), .B(G396), .Z(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1022), .A2(new_n1104), .A3(new_n1046), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1104), .B1(new_n1022), .B2(new_n1046), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1271), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G387), .A2(G390), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1263), .A3(new_n1270), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1206), .A2(new_n1207), .A3(new_n1001), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1206), .A2(new_n1207), .A3(KEYINPUT126), .A4(new_n1001), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1265), .A3(new_n1240), .A4(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(G213), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(G343), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1265), .B1(new_n1209), .B2(new_n1240), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1278), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G375), .A2(G378), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1282), .A2(new_n1240), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G378), .B1(new_n1280), .B2(new_n1279), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1285), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(KEYINPUT127), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1242), .A2(KEYINPUT60), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1115), .A2(new_n1121), .A3(KEYINPUT60), .A4(new_n1107), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1135), .A2(new_n1297), .A3(new_n728), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1261), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(G384), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1290), .A2(new_n1293), .A3(new_n1300), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1295), .A2(new_n1303), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1285), .A2(G2897), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1300), .B(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1289), .A2(new_n1294), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT61), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1277), .B1(new_n1305), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1295), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1313));
  OR2_X1    g1113(.A1(new_n1300), .A2(new_n1306), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1300), .A2(new_n1306), .ZN(new_n1315));
  AOI22_X1  g1115(.A1(new_n1314), .A2(new_n1315), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1304), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1312), .A2(new_n1313), .A3(new_n1318), .A4(new_n1309), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1311), .A2(new_n1319), .ZN(G405));
  NAND2_X1  g1120(.A1(new_n1290), .A2(new_n1266), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(new_n1300), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(new_n1313), .ZN(G402));
endmodule


