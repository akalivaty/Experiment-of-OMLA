//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G97), .C2(G257), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G1), .B2(G20), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT1), .Z(new_n217));
  INV_X1    g0017(.A(G1), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR3_X1   g0019(.A1(new_n218), .A2(new_n219), .A3(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT0), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n201), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n219), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n221), .A2(new_n222), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n223), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT64), .Z(new_n232));
  NOR2_X1   g0032(.A1(new_n217), .A2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT66), .Z(new_n235));
  XOR2_X1   g0035(.A(G226), .B(G232), .Z(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  INV_X1    g0040(.A(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT67), .B(G250), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n239), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(KEYINPUT85), .ZN(new_n253));
  AND2_X1   g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(new_n227), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(G244), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT4), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G283), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n258), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(G250), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n257), .B1(new_n266), .B2(KEYINPUT4), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n255), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT68), .B1(new_n254), .B2(new_n227), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n270), .A2(new_n271), .A3(G1), .A4(G13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n274), .A2(KEYINPUT5), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(KEYINPUT5), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G257), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n269), .B2(new_n272), .ZN(new_n283));
  INV_X1    g0083(.A(new_n279), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND3_X1   g0085(.A1(new_n268), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G200), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n253), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n289), .A2(new_n219), .A3(G1), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n218), .A2(G33), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n293), .A2(KEYINPUT70), .A3(new_n227), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT70), .B1(new_n293), .B2(new_n227), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n291), .B(new_n292), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G97), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n290), .A2(new_n297), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n299), .B(KEYINPUT84), .Z(new_n300));
  INV_X1    g0100(.A(KEYINPUT7), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n256), .A2(new_n301), .A3(G20), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n259), .A2(new_n260), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT7), .B1(new_n303), .B2(new_n219), .ZN(new_n304));
  OAI21_X1  g0104(.A(G107), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G107), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(KEYINPUT6), .A3(G97), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n297), .A2(new_n306), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G97), .A2(G107), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n307), .B1(new_n310), .B2(KEYINPUT6), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G20), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G20), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G77), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n305), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n293), .A2(new_n227), .ZN(new_n316));
  AOI211_X1 g0116(.A(new_n298), .B(new_n300), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n286), .A2(G190), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n268), .A2(new_n281), .A3(new_n285), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(KEYINPUT85), .A3(G200), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n288), .A2(new_n317), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n289), .A2(G1), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n219), .A2(G107), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n296), .A2(new_n306), .B1(KEYINPUT25), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(G20), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G116), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n323), .B(KEYINPUT23), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT22), .ZN(new_n330));
  OR2_X1    g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  AOI21_X1  g0132(.A(G20), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n333), .B2(G87), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n219), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(KEYINPUT22), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n328), .B(new_n329), .C1(new_n334), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT24), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n335), .B(KEYINPUT22), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT24), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(new_n328), .A4(new_n329), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n325), .B1(new_n342), .B2(new_n316), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n256), .A2(G250), .A3(new_n257), .ZN(new_n344));
  INV_X1    g0144(.A(G294), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n256), .A2(G1698), .ZN(new_n346));
  OAI221_X1 g0146(.A(new_n344), .B1(new_n326), .B2(new_n345), .C1(new_n346), .C2(new_n241), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n255), .B1(new_n280), .B2(G264), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n285), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G200), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(G190), .A3(new_n285), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n324), .A2(KEYINPUT25), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n343), .A2(new_n350), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n315), .A2(new_n316), .ZN(new_n354));
  INV_X1    g0154(.A(new_n300), .ZN(new_n355));
  INV_X1    g0155(.A(new_n298), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G169), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n319), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n268), .A2(new_n360), .A3(new_n281), .A4(new_n285), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n357), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n321), .A2(new_n353), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  AOI21_X1  g0166(.A(G1), .B1(new_n274), .B2(new_n276), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n273), .A2(G274), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G97), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n256), .A2(new_n257), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n211), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n255), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n367), .B1(new_n269), .B2(new_n272), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G238), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n366), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT77), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(new_n366), .A3(new_n376), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI211_X1 g0181(.A(new_n379), .B(new_n366), .C1(new_n374), .C2(new_n376), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n365), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n294), .A2(new_n295), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n219), .A2(G33), .ZN(new_n386));
  INV_X1    g0186(.A(G77), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n386), .A2(new_n387), .B1(new_n219), .B2(G68), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n388), .B(KEYINPUT78), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n313), .A2(G50), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n391), .A2(KEYINPUT11), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n322), .A2(G20), .A3(new_n212), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n393), .B(KEYINPUT12), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(KEYINPUT11), .ZN(new_n395));
  INV_X1    g0195(.A(new_n316), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n218), .A2(G20), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(G68), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n392), .A2(new_n394), .A3(new_n395), .A4(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n287), .B1(new_n378), .B2(new_n380), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n384), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n380), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n402), .A2(KEYINPUT77), .A3(new_n377), .ZN(new_n403));
  OAI21_X1  g0203(.A(G179), .B1(new_n403), .B2(new_n382), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT14), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(G169), .C1(new_n402), .C2(new_n377), .ZN(new_n406));
  OAI21_X1  g0206(.A(G169), .B1(new_n402), .B2(new_n377), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT14), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n401), .B1(new_n399), .B2(new_n409), .ZN(new_n410));
  XOR2_X1   g0210(.A(KEYINPUT8), .B(G58), .Z(new_n411));
  XOR2_X1   g0211(.A(KEYINPUT15), .B(G87), .Z(new_n412));
  AOI22_X1  g0212(.A1(new_n313), .A2(new_n411), .B1(new_n412), .B2(new_n327), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n219), .B2(new_n387), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n316), .B1(new_n387), .B2(new_n290), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n396), .A2(G77), .A3(new_n397), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT69), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n346), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n256), .A2(KEYINPUT69), .A3(G1698), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n213), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n256), .A2(new_n306), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n256), .A2(G232), .A3(new_n257), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n255), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n375), .A2(G244), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n427), .A2(KEYINPUT76), .A3(new_n428), .A4(new_n368), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n430));
  INV_X1    g0230(.A(new_n255), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n428), .B(new_n368), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT76), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n418), .B1(new_n435), .B2(new_n287), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n365), .B1(new_n429), .B2(new_n434), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n417), .B1(new_n435), .B2(G169), .ZN(new_n439));
  AOI21_X1  g0239(.A(G179), .B1(new_n429), .B2(new_n434), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n410), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n397), .A2(G50), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT73), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n445));
  OAI22_X1  g0245(.A1(new_n444), .A2(new_n445), .B1(G50), .B2(new_n291), .ZN(new_n446));
  XOR2_X1   g0246(.A(new_n446), .B(KEYINPUT74), .Z(new_n447));
  NAND2_X1  g0247(.A1(new_n203), .A2(G20), .ZN(new_n448));
  INV_X1    g0248(.A(G150), .ZN(new_n449));
  INV_X1    g0249(.A(new_n313), .ZN(new_n450));
  NAND3_X1  g0250(.A1(KEYINPUT71), .A2(KEYINPUT72), .A3(G58), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(KEYINPUT8), .C1(KEYINPUT71), .C2(G58), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT8), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(KEYINPUT72), .A3(G58), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OAI221_X1 g0256(.A(new_n448), .B1(new_n449), .B2(new_n450), .C1(new_n456), .C2(new_n386), .ZN(new_n457));
  INV_X1    g0257(.A(new_n385), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n447), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT9), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n303), .A2(G1698), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G222), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n420), .A2(new_n421), .ZN(new_n465));
  INV_X1    g0265(.A(G223), .ZN(new_n466));
  OAI221_X1 g0266(.A(new_n464), .B1(new_n387), .B2(new_n256), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n369), .B1(new_n467), .B2(new_n255), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n375), .A2(G226), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G200), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT9), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n460), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n468), .A2(G190), .A3(new_n469), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n462), .A2(new_n471), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT10), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n470), .A2(new_n358), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n470), .A2(G179), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n478), .A2(KEYINPUT75), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(KEYINPUT75), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n460), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(G68), .B1(new_n302), .B2(new_n304), .ZN(new_n483));
  AND2_X1   g0283(.A1(KEYINPUT71), .A2(G58), .ZN(new_n484));
  NOR2_X1   g0284(.A1(KEYINPUT71), .A2(G58), .ZN(new_n485));
  OAI21_X1  g0285(.A(G68), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n219), .B1(new_n486), .B2(new_n224), .ZN(new_n487));
  INV_X1    g0287(.A(G159), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n450), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT79), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT79), .ZN(new_n491));
  INV_X1    g0291(.A(new_n489), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT71), .B(G58), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n201), .B1(new_n493), .B2(G68), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n491), .B(new_n492), .C1(new_n494), .C2(new_n219), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n490), .A2(new_n495), .A3(KEYINPUT80), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT80), .B1(new_n490), .B2(new_n495), .ZN(new_n497));
  OAI211_X1 g0297(.A(KEYINPUT16), .B(new_n483), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n490), .A2(new_n483), .A3(new_n495), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT16), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n396), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n455), .A2(new_n397), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n503), .A2(new_n445), .B1(new_n291), .B2(new_n455), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT81), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n375), .A2(G232), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n368), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n466), .A2(new_n257), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n256), .B(new_n509), .C1(G226), .C2(new_n257), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G87), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n431), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT82), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(new_n365), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n511), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n255), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n517), .A2(new_n365), .A3(new_n368), .A4(new_n507), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT82), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n368), .A3(new_n507), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n287), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n502), .A2(new_n506), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT17), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n505), .B1(new_n498), .B2(new_n501), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(KEYINPUT17), .A3(new_n522), .ZN(new_n527));
  INV_X1    g0327(.A(new_n526), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n513), .A2(G179), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n520), .A2(G169), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT18), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT18), .ZN(new_n533));
  INV_X1    g0333(.A(new_n531), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n526), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n525), .B(new_n527), .C1(new_n532), .C2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  OR2_X1    g0337(.A1(new_n537), .A2(KEYINPUT83), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(KEYINPUT83), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n442), .B(new_n482), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n343), .A2(new_n352), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n349), .A2(new_n358), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n348), .A2(new_n360), .A3(new_n285), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT88), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n463), .A2(new_n545), .A3(G257), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT88), .B1(new_n372), .B2(new_n241), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n303), .A2(G303), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n256), .A2(G264), .A3(G1698), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n546), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n255), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n280), .A2(G270), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n285), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n322), .A2(G20), .A3(new_n207), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n291), .A2(G116), .A3(new_n396), .A4(new_n292), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n264), .B(new_n219), .C1(G33), .C2(new_n297), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(new_n316), .C1(new_n219), .C2(G116), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT20), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n554), .B(new_n555), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n553), .A2(G169), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n553), .A2(new_n360), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n561), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n553), .A2(KEYINPUT21), .A3(G169), .A4(new_n561), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n544), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n561), .B1(new_n553), .B2(G200), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n365), .B2(new_n553), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT19), .B1(new_n327), .B2(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(G68), .B2(new_n333), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n371), .A2(new_n219), .ZN(new_n574));
  NOR4_X1   g0374(.A1(KEYINPUT87), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT87), .ZN(new_n576));
  NOR2_X1   g0376(.A1(G87), .A2(G97), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n306), .ZN(new_n578));
  OAI211_X1 g0378(.A(KEYINPUT19), .B(new_n574), .C1(new_n575), .C2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n396), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n291), .A2(new_n412), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G87), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n296), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n277), .A2(G250), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n277), .A2(new_n282), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n273), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT86), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n261), .B2(new_n257), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n256), .A2(KEYINPUT86), .A3(G244), .A4(G1698), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n256), .A2(G238), .A3(new_n257), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G116), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n588), .B1(new_n594), .B2(new_n255), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n582), .B(new_n585), .C1(new_n595), .C2(new_n287), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n255), .ZN(new_n597));
  INV_X1    g0397(.A(new_n588), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n365), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n595), .A2(G169), .ZN(new_n602));
  INV_X1    g0402(.A(new_n412), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n296), .A2(new_n603), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n580), .A2(new_n604), .A3(new_n581), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n599), .A2(G179), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n571), .A2(new_n601), .A3(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n364), .A2(new_n540), .A3(new_n569), .A4(new_n610), .ZN(G372));
  AND3_X1   g0411(.A1(new_n357), .A2(new_n359), .A3(new_n361), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n319), .A2(KEYINPUT85), .A3(G200), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT85), .B1(new_n319), .B2(G200), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n613), .A2(new_n614), .A3(new_n357), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n615), .B2(new_n318), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT90), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n607), .A2(new_n602), .A3(new_n605), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n600), .B1(new_n596), .B2(KEYINPUT89), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n580), .A2(new_n584), .A3(new_n581), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT89), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n621), .C1(new_n287), .C2(new_n595), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n618), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n616), .A2(new_n617), .A3(new_n353), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n596), .A2(KEYINPUT89), .ZN(new_n625));
  INV_X1    g0425(.A(new_n600), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n609), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT90), .B1(new_n363), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n568), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n624), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n623), .A2(new_n634), .A3(new_n612), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n612), .A2(new_n601), .A3(new_n609), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n635), .A2(new_n609), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n540), .A2(new_n639), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n532), .A2(new_n535), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n409), .A2(new_n399), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n441), .B2(new_n401), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n525), .A2(new_n527), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n476), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n481), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT91), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT91), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n650), .B(new_n481), .C1(new_n646), .C2(new_n647), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n640), .A2(new_n652), .ZN(G369));
  NOR2_X1   g0453(.A1(new_n289), .A2(G20), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n218), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n561), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n630), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT92), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n630), .A2(new_n571), .A3(new_n661), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G330), .ZN(new_n666));
  INV_X1    g0466(.A(new_n660), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n544), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n353), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n343), .B2(new_n352), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n631), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n668), .A2(new_n671), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n630), .A2(new_n660), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT93), .B1(new_n676), .B2(new_n668), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT93), .ZN(new_n678));
  INV_X1    g0478(.A(new_n668), .ZN(new_n679));
  AOI211_X1 g0479(.A(new_n678), .B(new_n679), .C1(new_n675), .C2(new_n671), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n673), .A2(new_n681), .ZN(G399));
  OR3_X1    g0482(.A1(new_n575), .A2(new_n578), .A3(G116), .ZN(new_n683));
  INV_X1    g0483(.A(new_n220), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n683), .A2(new_n218), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT94), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  INV_X1    g0489(.A(new_n685), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n688), .B(new_n689), .C1(new_n225), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n627), .A2(new_n612), .A3(new_n609), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n618), .B1(new_n694), .B2(KEYINPUT26), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n616), .A2(new_n353), .A3(new_n623), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n693), .B(new_n695), .C1(new_n696), .C2(new_n569), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT29), .B1(new_n698), .B2(new_n660), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n660), .B1(new_n633), .B2(new_n638), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n699), .B1(KEYINPUT29), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n550), .A2(new_n255), .B1(new_n284), .B2(new_n283), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(G179), .A3(new_n552), .A4(new_n595), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n286), .A2(new_n348), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT95), .ZN(new_n708));
  OR3_X1    g0508(.A1(new_n705), .A2(new_n706), .A3(new_n703), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n595), .A2(G179), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n553), .A2(new_n710), .A3(new_n349), .A4(new_n319), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT95), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n712), .B(new_n703), .C1(new_n705), .C2(new_n706), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n708), .A2(new_n709), .A3(new_n711), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n660), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n569), .A2(new_n364), .A3(new_n610), .A4(new_n667), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n709), .A2(new_n711), .A3(new_n707), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n702), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n692), .B1(new_n724), .B2(G1), .ZN(G364));
  NOR2_X1   g0525(.A1(new_n287), .A2(G179), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n219), .A2(G190), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G179), .A2(G200), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI22_X1  g0532(.A1(G283), .A2(new_n729), .B1(new_n732), .B2(G329), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n360), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n727), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G311), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n219), .A2(new_n365), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n360), .A2(new_n287), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n738), .B1(G326), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n739), .A2(new_n734), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G322), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n219), .B1(new_n730), .B2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G294), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n739), .A2(new_n726), .ZN(new_n750));
  INV_X1    g0550(.A(G303), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n303), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n740), .A2(new_n727), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT33), .B(G317), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n743), .A2(new_n746), .A3(new_n749), .A4(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n750), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G87), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n729), .A2(G107), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n759), .A2(new_n760), .A3(new_n256), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT100), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n731), .A2(new_n488), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT32), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n747), .A2(new_n297), .ZN(new_n765));
  INV_X1    g0565(.A(new_n493), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n766), .A2(new_n744), .B1(new_n753), .B2(new_n212), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n765), .B(new_n767), .C1(G77), .C2(new_n736), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n762), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n741), .A2(new_n202), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n757), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n227), .B1(G20), .B2(new_n358), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n218), .B1(new_n654), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n685), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT96), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n256), .A2(new_n220), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT97), .Z(new_n779));
  XOR2_X1   g0579(.A(G355), .B(KEYINPUT98), .Z(new_n780));
  AOI22_X1  g0580(.A1(new_n779), .A2(new_n780), .B1(new_n207), .B2(new_n684), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT99), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n684), .A2(new_n256), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n248), .A2(G45), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G45), .B2(new_n225), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n782), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n772), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n777), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n790), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n773), .B(new_n792), .C1(new_n665), .C2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n776), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n666), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n665), .A2(G330), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(G396));
  NOR3_X1   g0598(.A1(new_n439), .A2(new_n440), .A3(new_n660), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n436), .A2(new_n437), .B1(new_n418), .B2(new_n667), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(new_n441), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n639), .A2(new_n801), .A3(new_n667), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(KEYINPUT102), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT102), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n700), .A2(new_n804), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n801), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n701), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(new_n723), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n795), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n772), .A2(new_n788), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n387), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G143), .A2(new_n745), .B1(new_n754), .B2(G150), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n815), .B2(new_n741), .C1(new_n488), .C2(new_n735), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT34), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n729), .A2(G68), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n817), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n256), .B1(new_n731), .B2(new_n821), .C1(new_n202), .C2(new_n750), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n493), .B2(new_n748), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G294), .A2(new_n745), .B1(new_n729), .B2(G87), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n825), .B1(new_n306), .B2(new_n750), .C1(new_n207), .C2(new_n735), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT101), .B(G283), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n303), .B1(new_n741), .B2(new_n751), .C1(new_n753), .C2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n826), .A2(new_n765), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n831), .B2(new_n731), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n824), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n777), .B1(new_n833), .B2(new_n772), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n813), .B(new_n834), .C1(new_n801), .C2(new_n789), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n811), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  OAI21_X1  g0637(.A(new_n483), .B1(new_n496), .B2(new_n497), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n385), .B1(new_n838), .B2(new_n500), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n504), .B1(new_n839), .B2(new_n498), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n658), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n536), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n523), .B1(new_n840), .B2(new_n534), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n841), .B1(new_n844), .B2(KEYINPUT104), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT104), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(new_n523), .C1(new_n840), .C2(new_n534), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n843), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n526), .A2(new_n534), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n658), .B(KEYINPUT105), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n528), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n850), .A2(new_n852), .A3(new_n843), .A4(new_n523), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n842), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n838), .A2(new_n500), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n458), .A3(new_n498), .ZN(new_n859));
  INV_X1    g0659(.A(new_n504), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n534), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n523), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT104), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n841), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n847), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n854), .B1(new_n865), .B2(KEYINPUT37), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n842), .A2(KEYINPUT38), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n857), .A2(new_n870), .ZN(new_n871));
  OR3_X1    g0671(.A1(new_n384), .A2(new_n399), .A3(new_n400), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n399), .A2(new_n660), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n643), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n399), .B(new_n660), .C1(new_n401), .C2(new_n409), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(KEYINPUT106), .A2(KEYINPUT31), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n715), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n714), .B(new_n660), .C1(KEYINPUT106), .C2(KEYINPUT31), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n718), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n877), .A2(new_n882), .A3(new_n807), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT40), .B1(new_n871), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n852), .ZN(new_n885));
  INV_X1    g0685(.A(new_n851), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n523), .B1(new_n526), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n887), .B2(new_n849), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n536), .A2(new_n885), .B1(new_n888), .B2(new_n853), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n866), .A2(new_n868), .B1(KEYINPUT38), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT107), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n852), .B1(new_n641), .B2(new_n645), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n888), .A2(new_n853), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n856), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT107), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n894), .B(new_n895), .C1(new_n866), .C2(new_n868), .ZN(new_n896));
  AND4_X1   g0696(.A1(KEYINPUT40), .A2(new_n876), .A3(new_n881), .A4(new_n801), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n891), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT108), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT108), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n891), .A2(new_n896), .A3(new_n897), .A4(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n884), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n540), .A2(new_n881), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n870), .A2(new_n906), .A3(new_n894), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n855), .A2(new_n856), .B1(new_n867), .B2(new_n869), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n907), .B1(new_n908), .B2(new_n906), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n643), .A2(new_n660), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n642), .A2(new_n886), .ZN(new_n912));
  INV_X1    g0712(.A(new_n799), .ZN(new_n913));
  AND4_X1   g0713(.A1(new_n804), .A2(new_n639), .A3(new_n667), .A4(new_n801), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n804), .B1(new_n700), .B2(new_n801), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(new_n871), .A3(new_n876), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n911), .A2(new_n912), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n540), .A2(new_n702), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n652), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  XNOR2_X1  g0721(.A(new_n905), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n218), .B2(new_n654), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n311), .B(KEYINPUT103), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n207), .B1(new_n924), .B2(KEYINPUT35), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n925), .B(new_n228), .C1(KEYINPUT35), .C2(new_n924), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT36), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n226), .A2(G77), .A3(new_n486), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(G50), .B2(new_n212), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(G1), .A3(new_n289), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n923), .A2(new_n927), .A3(new_n930), .ZN(G367));
  NOR2_X1   g0731(.A1(new_n747), .A2(new_n212), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n493), .A2(new_n758), .B1(new_n736), .B2(G50), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n933), .B1(new_n815), .B2(new_n731), .C1(new_n488), .C2(new_n753), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n932), .B(new_n934), .C1(G143), .C2(new_n742), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n256), .B1(new_n728), .B2(new_n387), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT113), .Z(new_n937));
  OAI211_X1 g0737(.A(new_n935), .B(new_n937), .C1(new_n449), .C2(new_n744), .ZN(new_n938));
  AOI22_X1  g0738(.A1(G294), .A2(new_n754), .B1(new_n732), .B2(G317), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n831), .B2(new_n741), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n758), .A2(KEYINPUT46), .A3(G116), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT46), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n750), .B2(new_n207), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n941), .B(new_n943), .C1(new_n306), .C2(new_n747), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n303), .B1(new_n744), .B2(new_n751), .C1(new_n828), .C2(new_n735), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n940), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n297), .B2(new_n728), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n938), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n777), .B1(new_n949), .B2(new_n772), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n791), .B1(new_n220), .B2(new_n603), .C1(new_n244), .C2(new_n784), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n620), .A2(new_n667), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n618), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n628), .B2(new_n952), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n950), .B(new_n951), .C1(new_n793), .C2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT114), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n616), .B1(new_n317), .B2(new_n667), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n612), .A2(new_n660), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n677), .A2(new_n680), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT44), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n960), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n959), .B1(new_n677), .B2(new_n680), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT45), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n673), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n960), .B(KEYINPUT44), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT45), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n963), .B(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n673), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n672), .A2(new_n630), .A3(new_n660), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT112), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT112), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(new_n674), .C2(new_n675), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(new_n666), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n965), .A2(new_n724), .A3(new_n970), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n724), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n685), .B(KEYINPUT41), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n775), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n673), .A2(new_n959), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT42), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n971), .A2(new_n983), .A3(new_n959), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT111), .ZN(new_n985));
  INV_X1    g0785(.A(new_n959), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT42), .B1(new_n676), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(KEYINPUT111), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n362), .B1(new_n957), .B2(new_n631), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n667), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n985), .A2(new_n987), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n981), .A2(new_n982), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n981), .B1(new_n991), .B2(new_n982), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n954), .B(KEYINPUT109), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n992), .A2(new_n993), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n992), .B2(new_n993), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n956), .B1(new_n980), .B2(new_n1000), .ZN(G387));
  NAND2_X1  g0801(.A1(new_n976), .A2(new_n724), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n975), .B1(new_n702), .B2(new_n723), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(new_n685), .A3(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G311), .A2(new_n754), .B1(new_n745), .B2(G317), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n751), .B2(new_n735), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G322), .B2(new_n742), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT48), .Z(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n345), .B2(new_n750), .C1(new_n747), .C2(new_n828), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n732), .A2(G326), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n256), .B1(new_n729), .B2(G116), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n603), .A2(new_n747), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n758), .A2(G77), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n256), .C1(new_n297), .C2(new_n728), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1016), .B(new_n1018), .C1(G150), .C2(new_n732), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n741), .A2(new_n488), .B1(new_n735), .B2(new_n212), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n455), .B2(new_n754), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1019), .B(new_n1021), .C1(new_n202), .C2(new_n744), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n772), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n784), .B1(new_n239), .B2(G45), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n683), .B2(new_n779), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n411), .A2(new_n202), .ZN(new_n1027));
  AOI21_X1  g0827(.A(G45), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(KEYINPUT50), .B2(new_n1027), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n683), .B(new_n1029), .C1(G68), .C2(G77), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1026), .A2(new_n1030), .B1(G107), .B2(new_n220), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n777), .B1(new_n1031), .B2(new_n791), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1024), .B(new_n1032), .C1(new_n674), .C2(new_n793), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1004), .B(new_n1033), .C1(new_n774), .C2(new_n975), .ZN(G393));
  NAND2_X1  g0834(.A1(new_n965), .A2(new_n970), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n1002), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1036), .A2(new_n685), .A3(new_n977), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT118), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(KEYINPUT118), .A3(new_n685), .A4(new_n977), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n965), .A2(new_n775), .A3(new_n970), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n758), .A2(new_n827), .B1(new_n732), .B2(G322), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1043), .A2(KEYINPUT115), .B1(G107), .B2(new_n729), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n303), .C1(KEYINPUT115), .C2(new_n1043), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT116), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n736), .A2(G294), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G317), .A2(new_n742), .B1(new_n745), .B2(G311), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT52), .Z(new_n1049));
  AOI22_X1  g0849(.A1(new_n754), .A2(G303), .B1(new_n748), .B2(G116), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT117), .Z(new_n1052));
  AOI22_X1  g0852(.A1(G68), .A2(new_n758), .B1(new_n736), .B2(new_n411), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n732), .A2(G143), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n202), .C2(new_n753), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n303), .B(new_n1055), .C1(G77), .C2(new_n748), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n741), .A2(new_n449), .B1(new_n744), .B2(new_n488), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT51), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(new_n583), .C2(new_n728), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1052), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n777), .B1(new_n1060), .B2(new_n772), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n791), .B1(new_n297), .B2(new_n220), .C1(new_n251), .C2(new_n784), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n986), .A2(new_n790), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1041), .A2(new_n1042), .A3(new_n1064), .ZN(G390));
  NAND2_X1  g0865(.A1(new_n441), .A2(new_n800), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n697), .A2(new_n1066), .A3(new_n667), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n913), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n910), .B1(new_n1068), .B2(new_n876), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1069), .A2(new_n891), .A3(new_n896), .ZN(new_n1070));
  INV_X1    g0870(.A(G330), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n807), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n721), .A3(new_n876), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n910), .B1(new_n916), .B2(new_n876), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1070), .B(new_n1074), .C1(new_n1075), .C2(new_n909), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1069), .A2(new_n891), .A3(new_n896), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n910), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n799), .B1(new_n803), .B2(new_n805), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n877), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n890), .A2(KEYINPUT39), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n871), .B2(KEYINPUT39), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1077), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n882), .A2(new_n807), .A3(new_n1071), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1084), .A2(new_n876), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1076), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n482), .B1(new_n538), .B2(new_n539), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n442), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1087), .A2(G330), .A3(new_n1088), .A4(new_n881), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n919), .A2(new_n652), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n876), .B1(new_n1072), .B2(new_n721), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n916), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1068), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1073), .B(new_n1093), .C1(new_n876), .C2(new_n1084), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1090), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n690), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n744), .A2(new_n821), .ZN(new_n1098));
  INV_X1    g0898(.A(G128), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n256), .B1(new_n753), .B2(new_n815), .C1(new_n1099), .C2(new_n741), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(G159), .C2(new_n748), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT54), .B(G143), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n202), .A2(new_n728), .B1(new_n735), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n758), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT53), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n750), .B2(new_n449), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1103), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1101), .B(new_n1107), .C1(new_n1108), .C2(new_n731), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n753), .A2(new_n306), .B1(new_n731), .B2(new_n345), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G283), .B2(new_n742), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n387), .B2(new_n747), .C1(new_n297), .C2(new_n735), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n745), .A2(G116), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n759), .A2(new_n1113), .A3(new_n819), .A4(new_n303), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1109), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n777), .B1(new_n1115), .B2(new_n772), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n909), .B2(new_n789), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n456), .B2(new_n812), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1086), .B2(new_n775), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1097), .A2(new_n1119), .ZN(G378));
  XNOR2_X1  g0920(.A(new_n482), .B(KEYINPUT55), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n461), .A2(new_n658), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT56), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1121), .B(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n788), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1099), .A2(new_n744), .B1(new_n750), .B2(new_n1102), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT120), .Z(new_n1127));
  OAI22_X1  g0927(.A1(new_n753), .A2(new_n821), .B1(new_n735), .B2(new_n815), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G150), .B2(new_n748), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1127), .B(new_n1129), .C1(new_n1108), .C2(new_n741), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT59), .Z(new_n1131));
  AOI21_X1  g0931(.A(G41), .B1(new_n732), .B2(G124), .ZN(new_n1132));
  AOI21_X1  g0932(.A(G33), .B1(new_n729), .B2(G159), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n202), .B1(new_n259), .B2(G41), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G116), .A2(new_n742), .B1(new_n754), .B2(G97), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n732), .A2(G283), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n729), .A2(new_n493), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1136), .A2(new_n303), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G107), .A2(new_n745), .B1(new_n736), .B2(new_n412), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1017), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1139), .A2(new_n1141), .A3(G41), .A4(new_n932), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1135), .B1(new_n1142), .B2(KEYINPUT58), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT119), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1143), .A2(new_n1144), .B1(KEYINPUT58), .B2(new_n1142), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1134), .B(new_n1145), .C1(new_n1144), .C2(new_n1143), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(new_n772), .B1(new_n202), .B2(new_n812), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1125), .A2(new_n776), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n899), .A2(new_n901), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n884), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1150), .A2(G330), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1124), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n902), .A2(G330), .A3(new_n1124), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(KEYINPUT121), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n918), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1154), .A2(KEYINPUT121), .A3(new_n918), .A4(new_n1155), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1149), .B1(new_n1160), .B2(new_n775), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1086), .A2(new_n1095), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1090), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT57), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n902), .A2(G330), .A3(new_n1124), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1124), .B1(new_n902), .B2(G330), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n1157), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n918), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1169));
  OAI211_X1 g0969(.A(KEYINPUT57), .B(new_n1164), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n685), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1161), .B1(new_n1165), .B2(new_n1171), .ZN(G375));
  AOI22_X1  g0972(.A1(G294), .A2(new_n742), .B1(new_n745), .B2(G283), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n306), .B2(new_n735), .C1(new_n207), .C2(new_n753), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1016), .B(new_n1174), .C1(G77), .C2(new_n729), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n750), .A2(new_n297), .B1(new_n731), .B2(new_n751), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT122), .Z(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n303), .A3(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n741), .A2(new_n821), .B1(new_n753), .B2(new_n1102), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G137), .B2(new_n745), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT123), .Z(new_n1181));
  OAI21_X1  g0981(.A(new_n1138), .B1(new_n202), .B2(new_n747), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n303), .B(new_n1182), .C1(G150), .C2(new_n736), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n750), .A2(new_n488), .B1(new_n731), .B2(new_n1099), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT124), .Z(new_n1185));
  NAND3_X1  g0985(.A1(new_n1181), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1178), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n777), .B1(new_n1187), .B2(new_n772), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n876), .B2(new_n789), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n212), .B2(new_n812), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1191), .B2(new_n775), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1090), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n979), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1194), .B2(new_n1095), .ZN(G381));
  INV_X1    g0995(.A(G378), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n1161), .C1(new_n1165), .C2(new_n1171), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1064), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1000), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n978), .A2(new_n979), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n775), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1203), .A3(new_n956), .A4(new_n1042), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1204), .A2(G396), .A3(G393), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(G384), .A2(G381), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1198), .A2(new_n1205), .A3(new_n1206), .ZN(G407));
  OAI211_X1 g1007(.A(G407), .B(G213), .C1(G343), .C2(new_n1197), .ZN(G409));
  INV_X1    g1008(.A(KEYINPUT60), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1193), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1163), .A2(new_n1191), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1090), .A2(new_n1092), .A3(KEYINPUT60), .A4(new_n1094), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n685), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1192), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n836), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT125), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G384), .A2(new_n1192), .A3(new_n1213), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT125), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1214), .A2(new_n1218), .A3(new_n836), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n659), .A2(G213), .A3(G2897), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1221), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1216), .A2(new_n1217), .A3(new_n1219), .A4(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1090), .B1(new_n1086), .B2(new_n1191), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n979), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n775), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n1196), .A3(new_n1148), .A4(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n659), .A2(G213), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n685), .B(new_n1170), .C1(new_n1227), .C2(KEYINPUT57), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1196), .B1(new_n1233), .B2(new_n1161), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1225), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G375), .A2(G378), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1220), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1236), .A2(new_n1231), .A3(new_n1230), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT63), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1232), .A2(new_n1234), .A3(new_n1220), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1241), .A2(KEYINPUT63), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(G393), .B(G396), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G390), .A2(G387), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1245), .A2(new_n1246), .A3(new_n1204), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n1245), .B2(new_n1204), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1244), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1245), .A2(new_n1204), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1244), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1249), .A2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1240), .A2(new_n1242), .A3(new_n1243), .A4(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1248), .A2(new_n1244), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1245), .A2(new_n1246), .A3(new_n1204), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1251), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1258), .B2(new_n1244), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1243), .B1(new_n1241), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT62), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1259), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1255), .A2(new_n1263), .ZN(G405));
  OAI21_X1  g1064(.A(KEYINPUT127), .B1(new_n1198), .B2(new_n1234), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT127), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1236), .A2(new_n1266), .A3(new_n1197), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1265), .A2(new_n1220), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1220), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1254), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1198), .A2(new_n1234), .A3(KEYINPUT127), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1266), .B1(new_n1236), .B2(new_n1197), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1237), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1265), .A2(new_n1220), .A3(new_n1267), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1259), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1270), .A2(new_n1275), .ZN(G402));
endmodule


