

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768;

  XOR2_X1 U371 ( .A(G113), .B(G116), .Z(n351) );
  XNOR2_X2 U372 ( .A(n528), .B(KEYINPUT19), .ZN(n573) );
  NOR2_X2 U373 ( .A1(n361), .A2(n359), .ZN(n618) );
  AND2_X1 U374 ( .A1(n386), .A2(n384), .ZN(n383) );
  AND2_X1 U375 ( .A1(n377), .A2(n375), .ZN(n374) );
  AND2_X1 U376 ( .A1(n368), .A2(n366), .ZN(n365) );
  NAND2_X1 U377 ( .A1(n619), .A2(n695), .ZN(n626) );
  NAND2_X1 U378 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U379 ( .A(n360), .B(n404), .ZN(n359) );
  XNOR2_X1 U380 ( .A(n596), .B(n576), .ZN(n602) );
  XNOR2_X1 U381 ( .A(n581), .B(n580), .ZN(n733) );
  OR2_X1 U382 ( .A1(n627), .A2(n567), .ZN(n479) );
  BUF_X1 U383 ( .A(G143), .Z(n638) );
  NAND2_X1 U384 ( .A1(n383), .A2(n380), .ZN(n388) );
  NAND2_X1 U385 ( .A1(n374), .A2(n371), .ZN(n379) );
  NAND2_X1 U386 ( .A1(n365), .A2(n363), .ZN(n370) );
  NAND2_X1 U387 ( .A1(n382), .A2(n381), .ZN(n380) );
  NAND2_X1 U388 ( .A1(n373), .A2(n364), .ZN(n363) );
  NAND2_X1 U389 ( .A1(n373), .A2(n372), .ZN(n371) );
  NAND2_X1 U390 ( .A1(n390), .A2(G217), .ZN(n673) );
  NAND2_X1 U391 ( .A1(n354), .A2(n352), .ZN(n361) );
  AND2_X1 U392 ( .A1(n357), .A2(n355), .ZN(n354) );
  AND2_X1 U393 ( .A1(n395), .A2(KEYINPUT44), .ZN(n616) );
  OR2_X1 U394 ( .A1(n713), .A2(n750), .ZN(n533) );
  OR2_X1 U395 ( .A1(n556), .A2(n751), .ZN(n512) );
  XNOR2_X1 U396 ( .A(n398), .B(KEYINPUT32), .ZN(n650) );
  NOR2_X1 U397 ( .A1(n609), .A2(n592), .ZN(n593) );
  AND2_X1 U398 ( .A1(n367), .A2(n680), .ZN(n366) );
  AND2_X1 U399 ( .A1(n376), .A2(n680), .ZN(n375) );
  INV_X1 U400 ( .A(n631), .ZN(n364) );
  OR2_X1 U401 ( .A1(n631), .A2(G210), .ZN(n367) );
  AND2_X1 U402 ( .A1(n385), .A2(n680), .ZN(n384) );
  XNOR2_X1 U403 ( .A(n479), .B(n478), .ZN(n527) );
  OR2_X1 U404 ( .A1(n679), .A2(G472), .ZN(n376) );
  INV_X1 U405 ( .A(n679), .ZN(n372) );
  INV_X1 U406 ( .A(n636), .ZN(n381) );
  XOR2_X1 U407 ( .A(KEYINPUT122), .B(n671), .Z(n672) );
  OR2_X1 U408 ( .A1(n636), .A2(G475), .ZN(n385) );
  NAND2_X1 U409 ( .A1(n353), .A2(KEYINPUT86), .ZN(n352) );
  INV_X1 U410 ( .A(n606), .ZN(n353) );
  NOR2_X1 U411 ( .A1(n356), .A2(n616), .ZN(n355) );
  NOR2_X1 U412 ( .A1(n605), .A2(n607), .ZN(n356) );
  NAND2_X1 U413 ( .A1(n606), .A2(n358), .ZN(n357) );
  AND2_X1 U414 ( .A1(n605), .A2(n607), .ZN(n358) );
  NAND2_X1 U415 ( .A1(n362), .A2(n405), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n617), .B(n406), .ZN(n362) );
  NAND2_X1 U417 ( .A1(n390), .A2(G478), .ZN(n663) );
  NAND2_X1 U418 ( .A1(n390), .A2(G469), .ZN(n669) );
  NAND2_X1 U419 ( .A1(n676), .A2(n369), .ZN(n368) );
  AND2_X1 U420 ( .A1(n631), .A2(G210), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n370), .B(n633), .ZN(G51) );
  INV_X1 U422 ( .A(n389), .ZN(n373) );
  NAND2_X1 U423 ( .A1(n389), .A2(n378), .ZN(n377) );
  AND2_X1 U424 ( .A1(n679), .A2(G472), .ZN(n378) );
  XNOR2_X1 U425 ( .A(n379), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U426 ( .A(n391), .ZN(n382) );
  NAND2_X1 U427 ( .A1(n391), .A2(n387), .ZN(n386) );
  AND2_X1 U428 ( .A1(n636), .A2(G475), .ZN(n387) );
  XNOR2_X1 U429 ( .A(n388), .B(n637), .ZN(G60) );
  NAND2_X1 U430 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U431 ( .A1(n626), .A2(n625), .ZN(n389) );
  NAND2_X1 U432 ( .A1(n626), .A2(n625), .ZN(n390) );
  NAND2_X1 U433 ( .A1(n626), .A2(n625), .ZN(n391) );
  NAND2_X1 U434 ( .A1(n626), .A2(n625), .ZN(n676) );
  NAND2_X2 U435 ( .A1(n740), .A2(n624), .ZN(n625) );
  NAND2_X1 U436 ( .A1(n656), .A2(n650), .ZN(n395) );
  INV_X1 U437 ( .A(n594), .ZN(n579) );
  INV_X1 U438 ( .A(n395), .ZN(n405) );
  XNOR2_X1 U439 ( .A(n590), .B(n400), .ZN(n613) );
  INV_X1 U440 ( .A(KEYINPUT89), .ZN(n400) );
  XNOR2_X1 U441 ( .A(n589), .B(n397), .ZN(n399) );
  INV_X1 U442 ( .A(KEYINPUT22), .ZN(n397) );
  XNOR2_X1 U443 ( .A(n540), .B(KEYINPUT1), .ZN(n577) );
  NOR2_X1 U444 ( .A1(G953), .A2(G237), .ZN(n486) );
  INV_X1 U445 ( .A(KEYINPUT72), .ZN(n404) );
  NAND2_X1 U446 ( .A1(n579), .A2(n578), .ZN(n581) );
  INV_X1 U447 ( .A(n614), .ZN(n578) );
  NOR2_X1 U448 ( .A1(n716), .A2(n610), .ZN(n427) );
  XNOR2_X1 U449 ( .A(KEYINPUT3), .B(G119), .ZN(n420) );
  XNOR2_X1 U450 ( .A(G128), .B(G119), .ZN(n428) );
  AND2_X1 U451 ( .A1(n519), .A2(n600), .ZN(n530) );
  NOR2_X1 U452 ( .A1(n535), .A2(n610), .ZN(n518) );
  NAND2_X1 U453 ( .A1(n399), .A2(n396), .ZN(n609) );
  NAND2_X1 U454 ( .A1(n392), .A2(n399), .ZN(n398) );
  NAND2_X1 U455 ( .A1(n613), .A2(n394), .ZN(n615) );
  XOR2_X1 U456 ( .A(n615), .B(KEYINPUT76), .Z(n392) );
  XOR2_X1 U457 ( .A(n688), .B(n474), .Z(n393) );
  AND2_X1 U458 ( .A1(n614), .A2(n698), .ZN(n394) );
  INV_X1 U459 ( .A(n590), .ZN(n396) );
  XNOR2_X2 U460 ( .A(n401), .B(KEYINPUT35), .ZN(n659) );
  NAND2_X1 U461 ( .A1(n402), .A2(n407), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n403), .B(KEYINPUT34), .ZN(n402) );
  NOR2_X2 U463 ( .A1(n602), .A2(n733), .ZN(n403) );
  INV_X1 U464 ( .A(KEYINPUT69), .ZN(n406) );
  INV_X1 U465 ( .A(n582), .ZN(n407) );
  BUF_X1 U466 ( .A(n527), .Z(n547) );
  AND2_X1 U467 ( .A1(n453), .A2(n452), .ZN(n408) );
  XOR2_X1 U468 ( .A(n521), .B(KEYINPUT64), .Z(n409) );
  INV_X1 U469 ( .A(KEYINPUT87), .ZN(n583) );
  XNOR2_X1 U470 ( .A(n584), .B(n583), .ZN(n606) );
  XNOR2_X1 U471 ( .A(n522), .B(n409), .ZN(n553) );
  BUF_X1 U472 ( .A(n627), .Z(n630) );
  INV_X1 U473 ( .A(KEYINPUT60), .ZN(n637) );
  XNOR2_X1 U474 ( .A(G902), .B(KEYINPUT15), .ZN(n621) );
  INV_X1 U475 ( .A(n621), .ZN(n567) );
  INV_X1 U476 ( .A(G902), .ZN(n510) );
  INV_X1 U477 ( .A(G237), .ZN(n410) );
  NAND2_X1 U478 ( .A1(n510), .A2(n410), .ZN(n476) );
  NAND2_X1 U479 ( .A1(n476), .A2(G214), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n411), .B(KEYINPUT91), .ZN(n716) );
  XNOR2_X2 U481 ( .A(KEYINPUT78), .B(G143), .ZN(n413) );
  INV_X1 U482 ( .A(G128), .ZN(n412) );
  XNOR2_X2 U483 ( .A(n413), .B(n412), .ZN(n505) );
  INV_X1 U484 ( .A(KEYINPUT65), .ZN(n414) );
  XNOR2_X1 U485 ( .A(n414), .B(KEYINPUT4), .ZN(n415) );
  XNOR2_X2 U486 ( .A(n505), .B(n415), .ZN(n755) );
  XNOR2_X1 U487 ( .A(KEYINPUT68), .B(G101), .ZN(n416) );
  XNOR2_X2 U488 ( .A(n755), .B(n416), .ZN(n458) );
  XOR2_X1 U489 ( .A(G146), .B(G137), .Z(n418) );
  NAND2_X1 U490 ( .A1(n486), .A2(G210), .ZN(n417) );
  XNOR2_X1 U491 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U492 ( .A(n419), .B(KEYINPUT5), .Z(n423) );
  XNOR2_X1 U493 ( .A(n351), .B(n420), .ZN(n468) );
  INV_X1 U494 ( .A(G134), .ZN(n421) );
  XNOR2_X1 U495 ( .A(n421), .B(G131), .ZN(n460) );
  XNOR2_X1 U496 ( .A(n468), .B(n460), .ZN(n422) );
  XNOR2_X1 U497 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U498 ( .A(n458), .B(n424), .ZN(n678) );
  NAND2_X1 U499 ( .A1(n678), .A2(n510), .ZN(n426) );
  INV_X1 U500 ( .A(G472), .ZN(n425) );
  XNOR2_X2 U501 ( .A(n426), .B(n425), .ZN(n610) );
  XNOR2_X1 U502 ( .A(KEYINPUT30), .B(n427), .ZN(n454) );
  XOR2_X1 U503 ( .A(KEYINPUT24), .B(G110), .Z(n429) );
  XNOR2_X1 U504 ( .A(n429), .B(n428), .ZN(n432) );
  INV_X2 U505 ( .A(G953), .ZN(n761) );
  NAND2_X1 U506 ( .A1(G234), .A2(n761), .ZN(n430) );
  XOR2_X1 U507 ( .A(KEYINPUT8), .B(n430), .Z(n506) );
  NAND2_X1 U508 ( .A1(G221), .A2(n506), .ZN(n431) );
  XNOR2_X1 U509 ( .A(n432), .B(n431), .ZN(n438) );
  XNOR2_X1 U510 ( .A(G146), .B(G125), .ZN(n470) );
  INV_X1 U511 ( .A(KEYINPUT10), .ZN(n433) );
  XNOR2_X1 U512 ( .A(n433), .B(G140), .ZN(n434) );
  XNOR2_X1 U513 ( .A(n470), .B(n434), .ZN(n756) );
  XNOR2_X1 U514 ( .A(KEYINPUT70), .B(G137), .ZN(n459) );
  INV_X1 U515 ( .A(KEYINPUT23), .ZN(n435) );
  XNOR2_X1 U516 ( .A(n459), .B(n435), .ZN(n436) );
  XNOR2_X1 U517 ( .A(n756), .B(n436), .ZN(n437) );
  XNOR2_X1 U518 ( .A(n438), .B(n437), .ZN(n671) );
  NAND2_X1 U519 ( .A1(n671), .A2(n510), .ZN(n443) );
  NAND2_X1 U520 ( .A1(n621), .A2(G234), .ZN(n439) );
  XNOR2_X1 U521 ( .A(n439), .B(KEYINPUT20), .ZN(n444) );
  NAND2_X1 U522 ( .A1(G217), .A2(n444), .ZN(n441) );
  XOR2_X1 U523 ( .A(KEYINPUT75), .B(KEYINPUT25), .Z(n440) );
  XNOR2_X1 U524 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U525 ( .A(n443), .B(n442), .ZN(n698) );
  NAND2_X1 U526 ( .A1(n444), .A2(G221), .ZN(n446) );
  INV_X1 U527 ( .A(KEYINPUT21), .ZN(n445) );
  XNOR2_X1 U528 ( .A(n446), .B(n445), .ZN(n585) );
  INV_X1 U529 ( .A(n585), .ZN(n697) );
  OR2_X1 U530 ( .A1(n698), .A2(n697), .ZN(n701) );
  INV_X1 U531 ( .A(n701), .ZN(n453) );
  NAND2_X1 U532 ( .A1(G234), .A2(G237), .ZN(n447) );
  XNOR2_X1 U533 ( .A(n447), .B(KEYINPUT14), .ZN(n729) );
  NAND2_X1 U534 ( .A1(G953), .A2(G902), .ZN(n568) );
  NOR2_X1 U535 ( .A1(G900), .A2(n568), .ZN(n448) );
  NAND2_X1 U536 ( .A1(n729), .A2(n448), .ZN(n449) );
  XNOR2_X1 U537 ( .A(n449), .B(KEYINPUT105), .ZN(n451) );
  AND2_X1 U538 ( .A1(G952), .A2(n761), .ZN(n569) );
  AND2_X1 U539 ( .A1(n729), .A2(n569), .ZN(n450) );
  NOR2_X1 U540 ( .A1(n451), .A2(n450), .ZN(n516) );
  INV_X1 U541 ( .A(n516), .ZN(n452) );
  NAND2_X1 U542 ( .A1(n454), .A2(n408), .ZN(n545) );
  XNOR2_X1 U543 ( .A(G107), .B(G104), .ZN(n456) );
  XNOR2_X1 U544 ( .A(KEYINPUT74), .B(G110), .ZN(n455) );
  XNOR2_X1 U545 ( .A(n456), .B(n455), .ZN(n686) );
  XNOR2_X1 U546 ( .A(n686), .B(KEYINPUT71), .ZN(n457) );
  XNOR2_X2 U547 ( .A(n458), .B(n457), .ZN(n475) );
  XNOR2_X1 U548 ( .A(n460), .B(n459), .ZN(n757) );
  XNOR2_X1 U549 ( .A(G146), .B(G140), .ZN(n462) );
  NAND2_X1 U550 ( .A1(n761), .A2(G227), .ZN(n461) );
  XNOR2_X1 U551 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U552 ( .A(n757), .B(n463), .ZN(n464) );
  XNOR2_X1 U553 ( .A(n475), .B(n464), .ZN(n665) );
  OR2_X2 U554 ( .A1(n665), .A2(G902), .ZN(n466) );
  INV_X1 U555 ( .A(G469), .ZN(n465) );
  XNOR2_X2 U556 ( .A(n466), .B(n465), .ZN(n540) );
  NOR2_X1 U557 ( .A1(n545), .A2(n540), .ZN(n481) );
  XNOR2_X1 U558 ( .A(KEYINPUT16), .B(G122), .ZN(n467) );
  XNOR2_X1 U559 ( .A(n468), .B(n467), .ZN(n688) );
  XNOR2_X1 U560 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n469) );
  XNOR2_X1 U561 ( .A(n470), .B(n469), .ZN(n473) );
  NAND2_X1 U562 ( .A1(n761), .A2(G224), .ZN(n471) );
  XNOR2_X1 U563 ( .A(n471), .B(KEYINPUT90), .ZN(n472) );
  XNOR2_X1 U564 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U565 ( .A(n475), .B(n393), .ZN(n627) );
  NAND2_X1 U566 ( .A1(n476), .A2(G210), .ZN(n477) );
  XNOR2_X1 U567 ( .A(n477), .B(KEYINPUT79), .ZN(n478) );
  INV_X1 U568 ( .A(n547), .ZN(n560) );
  INV_X1 U569 ( .A(KEYINPUT38), .ZN(n480) );
  XNOR2_X1 U570 ( .A(n560), .B(n480), .ZN(n717) );
  INV_X1 U571 ( .A(n717), .ZN(n714) );
  NAND2_X1 U572 ( .A1(n481), .A2(n714), .ZN(n485) );
  XNOR2_X1 U573 ( .A(KEYINPUT85), .B(KEYINPUT39), .ZN(n483) );
  INV_X1 U574 ( .A(KEYINPUT73), .ZN(n482) );
  XNOR2_X1 U575 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U576 ( .A(n485), .B(n484), .ZN(n556) );
  NAND2_X1 U577 ( .A1(G214), .A2(n486), .ZN(n487) );
  XNOR2_X1 U578 ( .A(n756), .B(n487), .ZN(n494) );
  XNOR2_X1 U579 ( .A(n638), .B(G131), .ZN(n488) );
  XNOR2_X1 U580 ( .A(n488), .B(G104), .ZN(n492) );
  XOR2_X1 U581 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n490) );
  XNOR2_X1 U582 ( .A(G113), .B(G122), .ZN(n489) );
  XNOR2_X1 U583 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U584 ( .A(n492), .B(n491), .Z(n493) );
  XNOR2_X1 U585 ( .A(n494), .B(n493), .ZN(n635) );
  NOR2_X1 U586 ( .A1(G902), .A2(n635), .ZN(n496) );
  XNOR2_X1 U587 ( .A(KEYINPUT94), .B(KEYINPUT13), .ZN(n495) );
  XNOR2_X1 U588 ( .A(n496), .B(n495), .ZN(n498) );
  INV_X1 U589 ( .A(G475), .ZN(n497) );
  XNOR2_X1 U590 ( .A(n498), .B(n497), .ZN(n543) );
  XOR2_X1 U591 ( .A(G122), .B(G107), .Z(n500) );
  XNOR2_X1 U592 ( .A(G116), .B(G134), .ZN(n499) );
  XNOR2_X1 U593 ( .A(n500), .B(n499), .ZN(n504) );
  XOR2_X1 U594 ( .A(KEYINPUT96), .B(KEYINPUT9), .Z(n502) );
  XNOR2_X1 U595 ( .A(KEYINPUT7), .B(KEYINPUT95), .ZN(n501) );
  XNOR2_X1 U596 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U597 ( .A(n504), .B(n503), .Z(n509) );
  NAND2_X1 U598 ( .A1(G217), .A2(n506), .ZN(n507) );
  XNOR2_X1 U599 ( .A(n505), .B(n507), .ZN(n508) );
  XNOR2_X1 U600 ( .A(n509), .B(n508), .ZN(n661) );
  NAND2_X1 U601 ( .A1(n661), .A2(n510), .ZN(n511) );
  XNOR2_X1 U602 ( .A(n511), .B(G478), .ZN(n523) );
  OR2_X1 U603 ( .A1(n543), .A2(n523), .ZN(n751) );
  XNOR2_X1 U604 ( .A(n512), .B(KEYINPUT40), .ZN(n642) );
  INV_X1 U605 ( .A(n523), .ZN(n542) );
  AND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n719) );
  INV_X1 U607 ( .A(n716), .ZN(n526) );
  NAND2_X1 U608 ( .A1(n719), .A2(n526), .ZN(n513) );
  OR2_X1 U609 ( .A1(n717), .A2(n513), .ZN(n515) );
  XNOR2_X1 U610 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n514) );
  XNOR2_X1 U611 ( .A(n515), .B(n514), .ZN(n711) );
  INV_X1 U612 ( .A(n698), .ZN(n591) );
  NOR2_X1 U613 ( .A1(n516), .A2(n591), .ZN(n517) );
  NAND2_X1 U614 ( .A1(n517), .A2(n585), .ZN(n535) );
  XNOR2_X1 U615 ( .A(n518), .B(KEYINPUT28), .ZN(n519) );
  INV_X1 U616 ( .A(n540), .ZN(n600) );
  NAND2_X1 U617 ( .A1(n711), .A2(n530), .ZN(n520) );
  XNOR2_X1 U618 ( .A(n520), .B(KEYINPUT42), .ZN(n641) );
  NAND2_X1 U619 ( .A1(n642), .A2(n641), .ZN(n522) );
  XNOR2_X1 U620 ( .A(KEYINPUT84), .B(KEYINPUT46), .ZN(n521) );
  NAND2_X1 U621 ( .A1(n543), .A2(n523), .ZN(n524) );
  XNOR2_X1 U622 ( .A(n524), .B(KEYINPUT97), .ZN(n651) );
  INV_X1 U623 ( .A(n751), .ZN(n653) );
  NOR2_X1 U624 ( .A1(n651), .A2(n653), .ZN(n525) );
  XNOR2_X1 U625 ( .A(n525), .B(KEYINPUT98), .ZN(n713) );
  NAND2_X1 U626 ( .A1(n527), .A2(n526), .ZN(n528) );
  BUF_X1 U627 ( .A(n573), .Z(n529) );
  NAND2_X1 U628 ( .A1(n530), .A2(n529), .ZN(n532) );
  INV_X1 U629 ( .A(KEYINPUT77), .ZN(n531) );
  XNOR2_X1 U630 ( .A(n532), .B(n531), .ZN(n750) );
  XNOR2_X1 U631 ( .A(n533), .B(KEYINPUT47), .ZN(n551) );
  XNOR2_X1 U632 ( .A(KEYINPUT99), .B(KEYINPUT6), .ZN(n534) );
  XNOR2_X1 U633 ( .A(n610), .B(n534), .ZN(n614) );
  NOR2_X1 U634 ( .A1(n535), .A2(n614), .ZN(n536) );
  NAND2_X1 U635 ( .A1(n653), .A2(n536), .ZN(n537) );
  NOR2_X1 U636 ( .A1(n537), .A2(n716), .ZN(n558) );
  NAND2_X1 U637 ( .A1(n558), .A2(n547), .ZN(n539) );
  XNOR2_X1 U638 ( .A(KEYINPUT107), .B(KEYINPUT36), .ZN(n538) );
  XNOR2_X1 U639 ( .A(n539), .B(n538), .ZN(n541) );
  INV_X1 U640 ( .A(n577), .ZN(n590) );
  NAND2_X1 U641 ( .A1(n541), .A2(n613), .ZN(n754) );
  OR2_X1 U642 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U643 ( .A(n544), .B(KEYINPUT104), .ZN(n582) );
  NOR2_X1 U644 ( .A1(n545), .A2(n582), .ZN(n546) );
  AND2_X1 U645 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U646 ( .A1(n548), .A2(n600), .ZN(n639) );
  XNOR2_X1 U647 ( .A(n639), .B(KEYINPUT80), .ZN(n549) );
  NAND2_X1 U648 ( .A1(n754), .A2(n549), .ZN(n550) );
  NOR2_X1 U649 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U650 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U651 ( .A(KEYINPUT83), .B(KEYINPUT48), .ZN(n554) );
  XNOR2_X1 U652 ( .A(n555), .B(n554), .ZN(n563) );
  INV_X1 U653 ( .A(n651), .ZN(n745) );
  OR2_X1 U654 ( .A1(n556), .A2(n745), .ZN(n557) );
  XNOR2_X1 U655 ( .A(n557), .B(KEYINPUT108), .ZN(n768) );
  NAND2_X1 U656 ( .A1(n558), .A2(n396), .ZN(n559) );
  XNOR2_X1 U657 ( .A(n559), .B(KEYINPUT43), .ZN(n561) );
  NAND2_X1 U658 ( .A1(n561), .A2(n560), .ZN(n640) );
  AND2_X1 U659 ( .A1(n768), .A2(n640), .ZN(n562) );
  XOR2_X1 U660 ( .A(KEYINPUT82), .B(n564), .Z(n760) );
  INV_X1 U661 ( .A(n564), .ZN(n565) );
  NAND2_X1 U662 ( .A1(n565), .A2(KEYINPUT2), .ZN(n566) );
  AND2_X1 U663 ( .A1(n760), .A2(n566), .ZN(n696) );
  AND2_X1 U664 ( .A1(n567), .A2(n696), .ZN(n619) );
  NOR2_X1 U665 ( .A1(G898), .A2(n568), .ZN(n570) );
  OR2_X1 U666 ( .A1(n570), .A2(n569), .ZN(n571) );
  AND2_X1 U667 ( .A1(n729), .A2(n571), .ZN(n572) );
  XNOR2_X1 U668 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n574) );
  XNOR2_X2 U669 ( .A(n575), .B(n574), .ZN(n596) );
  INV_X1 U670 ( .A(KEYINPUT92), .ZN(n576) );
  OR2_X2 U671 ( .A1(n577), .A2(n701), .ZN(n594) );
  XNOR2_X1 U672 ( .A(KEYINPUT103), .B(KEYINPUT33), .ZN(n580) );
  NAND2_X1 U673 ( .A1(n659), .A2(KEYINPUT44), .ZN(n584) );
  NAND2_X1 U674 ( .A1(n719), .A2(n585), .ZN(n587) );
  INV_X1 U675 ( .A(KEYINPUT100), .ZN(n586) );
  XNOR2_X1 U676 ( .A(n587), .B(n586), .ZN(n588) );
  NAND2_X1 U677 ( .A1(n596), .A2(n588), .ZN(n589) );
  NAND2_X1 U678 ( .A1(n614), .A2(n591), .ZN(n592) );
  XOR2_X1 U679 ( .A(KEYINPUT101), .B(n593), .Z(n658) );
  NOR2_X1 U680 ( .A1(n594), .A2(n610), .ZN(n595) );
  XNOR2_X1 U681 ( .A(n595), .B(KEYINPUT93), .ZN(n709) );
  INV_X1 U682 ( .A(n596), .ZN(n597) );
  NOR2_X1 U683 ( .A1(n709), .A2(n597), .ZN(n598) );
  XOR2_X1 U684 ( .A(KEYINPUT31), .B(n598), .Z(n654) );
  INV_X1 U685 ( .A(n610), .ZN(n705) );
  NOR2_X1 U686 ( .A1(n705), .A2(n701), .ZN(n599) );
  NAND2_X1 U687 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U688 ( .A1(n602), .A2(n601), .ZN(n646) );
  NOR2_X1 U689 ( .A1(n654), .A2(n646), .ZN(n603) );
  NOR2_X1 U690 ( .A1(n603), .A2(n713), .ZN(n604) );
  NOR2_X1 U691 ( .A1(n658), .A2(n604), .ZN(n605) );
  INV_X1 U692 ( .A(KEYINPUT86), .ZN(n607) );
  INV_X1 U693 ( .A(KEYINPUT102), .ZN(n608) );
  XNOR2_X1 U694 ( .A(n609), .B(n608), .ZN(n612) );
  AND2_X1 U695 ( .A1(n610), .A2(n698), .ZN(n611) );
  NAND2_X1 U696 ( .A1(n612), .A2(n611), .ZN(n656) );
  NOR2_X1 U697 ( .A1(n659), .A2(KEYINPUT44), .ZN(n617) );
  XNOR2_X1 U698 ( .A(n618), .B(KEYINPUT45), .ZN(n620) );
  INV_X1 U699 ( .A(n620), .ZN(n695) );
  OR2_X2 U700 ( .A1(n620), .A2(n564), .ZN(n740) );
  XOR2_X1 U701 ( .A(KEYINPUT81), .B(n621), .Z(n623) );
  INV_X1 U702 ( .A(KEYINPUT2), .ZN(n622) );
  NOR2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U704 ( .A(KEYINPUT88), .B(KEYINPUT54), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n628), .B(KEYINPUT55), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n630), .B(n629), .ZN(n631) );
  INV_X1 U707 ( .A(G952), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n632), .A2(G953), .ZN(n680) );
  INV_X1 U709 ( .A(KEYINPUT56), .ZN(n633) );
  XNOR2_X1 U710 ( .A(KEYINPUT66), .B(KEYINPUT59), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(G45) );
  XNOR2_X1 U713 ( .A(n640), .B(G140), .ZN(G42) );
  XNOR2_X1 U714 ( .A(n641), .B(G137), .ZN(G39) );
  XNOR2_X1 U715 ( .A(n642), .B(G131), .ZN(G33) );
  NAND2_X1 U716 ( .A1(n646), .A2(n653), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n643), .B(G104), .ZN(G6) );
  XOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n645) );
  XNOR2_X1 U719 ( .A(G107), .B(KEYINPUT111), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n645), .B(n644), .ZN(n648) );
  NAND2_X1 U721 ( .A1(n646), .A2(n651), .ZN(n647) );
  XOR2_X1 U722 ( .A(n648), .B(n647), .Z(G9) );
  XOR2_X1 U723 ( .A(G119), .B(KEYINPUT127), .Z(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(G21) );
  NAND2_X1 U725 ( .A1(n654), .A2(n651), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n652), .B(G116), .ZN(G18) );
  NAND2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n655), .B(G113), .ZN(G15) );
  XNOR2_X1 U729 ( .A(n656), .B(G110), .ZN(G12) );
  XOR2_X1 U730 ( .A(G101), .B(KEYINPUT110), .Z(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(G3) );
  BUF_X1 U732 ( .A(n659), .Z(n660) );
  XOR2_X1 U733 ( .A(n660), .B(G122), .Z(G24) );
  XNOR2_X1 U734 ( .A(n661), .B(KEYINPUT121), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(n664) );
  INV_X1 U736 ( .A(n680), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n664), .A2(n674), .ZN(G63) );
  XOR2_X1 U738 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n666) );
  XNOR2_X1 U739 ( .A(n666), .B(KEYINPUT58), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n665), .B(n667), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U742 ( .A1(n670), .A2(n674), .ZN(G54) );
  XNOR2_X1 U743 ( .A(n673), .B(n672), .ZN(n675) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(G66) );
  XOR2_X1 U745 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n677) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U747 ( .A1(n761), .A2(n695), .ZN(n684) );
  NAND2_X1 U748 ( .A1(G953), .A2(G224), .ZN(n681) );
  XNOR2_X1 U749 ( .A(KEYINPUT61), .B(n681), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n682), .A2(G898), .ZN(n683) );
  NAND2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n694) );
  XOR2_X1 U752 ( .A(G101), .B(KEYINPUT124), .Z(n685) );
  XNOR2_X1 U753 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U754 ( .A(n688), .B(n687), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n761), .A2(G898), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n692) );
  XNOR2_X1 U757 ( .A(KEYINPUT123), .B(KEYINPUT125), .ZN(n691) );
  XNOR2_X1 U758 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n694), .B(n693), .ZN(G69) );
  AND2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n739) );
  XOR2_X1 U761 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n700) );
  NAND2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U763 ( .A(n700), .B(n699), .ZN(n707) );
  NAND2_X1 U764 ( .A1(n396), .A2(n701), .ZN(n702) );
  XNOR2_X1 U765 ( .A(n702), .B(KEYINPUT115), .ZN(n703) );
  XNOR2_X1 U766 ( .A(KEYINPUT50), .B(n703), .ZN(n704) );
  NOR2_X1 U767 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U769 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U770 ( .A(KEYINPUT51), .B(n710), .ZN(n712) );
  INV_X1 U771 ( .A(n711), .ZN(n734) );
  NOR2_X1 U772 ( .A1(n712), .A2(n734), .ZN(n727) );
  NOR2_X1 U773 ( .A1(n713), .A2(n716), .ZN(n715) );
  NAND2_X1 U774 ( .A1(n715), .A2(n714), .ZN(n722) );
  NAND2_X1 U775 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U776 ( .A(n718), .B(KEYINPUT116), .ZN(n720) );
  NAND2_X1 U777 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U778 ( .A1(n722), .A2(n721), .ZN(n724) );
  INV_X1 U779 ( .A(n733), .ZN(n723) );
  NAND2_X1 U780 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U781 ( .A(n725), .B(KEYINPUT117), .ZN(n726) );
  NOR2_X1 U782 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U783 ( .A(n728), .B(KEYINPUT52), .ZN(n731) );
  NAND2_X1 U784 ( .A1(n729), .A2(G952), .ZN(n730) );
  NOR2_X1 U785 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U786 ( .A(KEYINPUT118), .B(n732), .Z(n737) );
  NOR2_X1 U787 ( .A1(n733), .A2(n734), .ZN(n735) );
  NOR2_X1 U788 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U789 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U790 ( .A1(n739), .A2(n738), .ZN(n742) );
  NAND2_X1 U791 ( .A1(n740), .A2(KEYINPUT2), .ZN(n741) );
  NAND2_X1 U792 ( .A1(n742), .A2(n741), .ZN(n744) );
  XNOR2_X1 U793 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n743) );
  XNOR2_X1 U794 ( .A(n744), .B(n743), .ZN(G75) );
  NOR2_X1 U795 ( .A1(n750), .A2(n745), .ZN(n749) );
  XOR2_X1 U796 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n747) );
  XNOR2_X1 U797 ( .A(G128), .B(KEYINPUT29), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X1 U799 ( .A(n749), .B(n748), .ZN(G30) );
  NOR2_X1 U800 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U801 ( .A(G146), .B(n752), .Z(G48) );
  XOR2_X1 U802 ( .A(G125), .B(KEYINPUT37), .Z(n753) );
  XNOR2_X1 U803 ( .A(n754), .B(n753), .ZN(G27) );
  XNOR2_X1 U804 ( .A(n757), .B(n756), .ZN(n758) );
  XNOR2_X1 U805 ( .A(n758), .B(KEYINPUT126), .ZN(n759) );
  XOR2_X1 U806 ( .A(n755), .B(n759), .Z(n763) );
  XNOR2_X1 U807 ( .A(n760), .B(n763), .ZN(n762) );
  NAND2_X1 U808 ( .A1(n762), .A2(n761), .ZN(n767) );
  XOR2_X1 U809 ( .A(G227), .B(n763), .Z(n764) );
  NAND2_X1 U810 ( .A1(n764), .A2(G900), .ZN(n765) );
  NAND2_X1 U811 ( .A1(n765), .A2(G953), .ZN(n766) );
  NAND2_X1 U812 ( .A1(n767), .A2(n766), .ZN(G72) );
  XNOR2_X1 U813 ( .A(G134), .B(n768), .ZN(G36) );
endmodule

