

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739;

  OR2_X1 U374 ( .A1(n695), .A2(G902), .ZN(n355) );
  INV_X1 U375 ( .A(n389), .ZN(n354) );
  XNOR2_X1 U376 ( .A(n406), .B(n405), .ZN(n513) );
  XNOR2_X1 U377 ( .A(n720), .B(G146), .ZN(n388) );
  XNOR2_X1 U378 ( .A(n446), .B(G128), .ZN(n419) );
  XNOR2_X2 U379 ( .A(n355), .B(n354), .ZN(n561) );
  NOR2_X2 U380 ( .A1(n484), .A2(n497), .ZN(n412) );
  INV_X1 U381 ( .A(G953), .ZN(n724) );
  XOR2_X1 U382 ( .A(G475), .B(n459), .Z(n356) );
  NOR2_X2 U383 ( .A1(n547), .A2(n546), .ZN(n578) );
  NOR2_X2 U384 ( .A1(n643), .A2(KEYINPUT2), .ZN(n645) );
  OR2_X2 U385 ( .A1(n547), .A2(n518), .ZN(n519) );
  OR2_X2 U386 ( .A1(n705), .A2(G902), .ZN(n406) );
  XOR2_X2 U387 ( .A(G137), .B(G140), .Z(n396) );
  BUF_X1 U388 ( .A(n561), .Z(n357) );
  XNOR2_X2 U389 ( .A(n475), .B(n474), .ZN(n735) );
  XNOR2_X1 U390 ( .A(n404), .B(KEYINPUT25), .ZN(n405) );
  XNOR2_X1 U391 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U392 ( .A(n522), .B(n521), .ZN(n562) );
  NAND2_X1 U393 ( .A1(n694), .A2(G472), .ZN(n600) );
  AND2_X1 U394 ( .A1(n601), .A2(G953), .ZN(n708) );
  XNOR2_X1 U395 ( .A(G119), .B(G113), .ZN(n370) );
  XNOR2_X1 U396 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U397 ( .A(n419), .B(n366), .ZN(n471) );
  INV_X1 U398 ( .A(G134), .ZN(n366) );
  XNOR2_X1 U399 ( .A(n386), .B(n385), .ZN(n387) );
  AND2_X1 U400 ( .A1(n723), .A2(n641), .ZN(n642) );
  INV_X1 U401 ( .A(n665), .ZN(n491) );
  XNOR2_X1 U402 ( .A(n402), .B(n363), .ZN(n705) );
  XNOR2_X1 U403 ( .A(n362), .B(n397), .ZN(n398) );
  NOR2_X1 U404 ( .A1(n582), .A2(n581), .ZN(n583) );
  AND2_X2 U405 ( .A1(n562), .A2(n364), .ZN(n632) );
  XNOR2_X1 U406 ( .A(n600), .B(n365), .ZN(n602) );
  XOR2_X1 U407 ( .A(n382), .B(n422), .Z(n358) );
  XOR2_X1 U408 ( .A(KEYINPUT70), .B(KEYINPUT48), .Z(n359) );
  NAND2_X1 U409 ( .A1(n586), .A2(n360), .ZN(n723) );
  AND2_X1 U410 ( .A1(n669), .A2(n357), .ZN(n530) );
  AND2_X1 U411 ( .A1(n585), .A2(n640), .ZN(n360) );
  OR2_X1 U412 ( .A1(n555), .A2(n537), .ZN(n361) );
  XOR2_X1 U413 ( .A(n396), .B(n395), .Z(n362) );
  AND2_X1 U414 ( .A1(n467), .A2(G221), .ZN(n363) );
  AND2_X1 U415 ( .A1(n357), .A2(n523), .ZN(n364) );
  XOR2_X1 U416 ( .A(n599), .B(KEYINPUT113), .Z(n365) );
  NOR2_X1 U417 ( .A1(n540), .A2(n539), .ZN(n541) );
  INV_X1 U418 ( .A(KEYINPUT4), .ZN(n367) );
  INV_X1 U419 ( .A(KEYINPUT46), .ZN(n573) );
  XNOR2_X1 U420 ( .A(n388), .B(n379), .ZN(n598) );
  XNOR2_X1 U421 ( .A(G122), .B(G104), .ZN(n448) );
  XNOR2_X1 U422 ( .A(n719), .B(n358), .ZN(n386) );
  XNOR2_X1 U423 ( .A(KEYINPUT105), .B(n530), .ZN(n531) );
  XNOR2_X1 U424 ( .A(n471), .B(n369), .ZN(n720) );
  INV_X1 U425 ( .A(KEYINPUT34), .ZN(n444) );
  XNOR2_X1 U426 ( .A(n577), .B(n359), .ZN(n586) );
  NOR2_X1 U427 ( .A1(n555), .A2(n652), .ZN(n557) );
  BUF_X1 U428 ( .A(n694), .Z(n704) );
  INV_X1 U429 ( .A(KEYINPUT35), .ZN(n474) );
  INV_X2 U430 ( .A(G143), .ZN(n446) );
  XNOR2_X1 U431 ( .A(G131), .B(KEYINPUT69), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n370), .B(KEYINPUT3), .ZN(n373) );
  INV_X1 U433 ( .A(KEYINPUT81), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n371), .B(G101), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n416) );
  XOR2_X1 U436 ( .A(KEYINPUT73), .B(KEYINPUT5), .Z(n375) );
  XNOR2_X1 U437 ( .A(G116), .B(G137), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n377) );
  NOR2_X1 U439 ( .A1(G953), .A2(G237), .ZN(n450) );
  NAND2_X1 U440 ( .A1(n450), .A2(G210), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n416), .B(n378), .ZN(n379) );
  NOR2_X1 U443 ( .A1(n598), .A2(G902), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n380), .B(G472), .ZN(n518) );
  INV_X1 U445 ( .A(n518), .ZN(n532) );
  XNOR2_X1 U446 ( .A(n532), .B(KEYINPUT6), .ZN(n484) );
  XOR2_X1 U447 ( .A(KEYINPUT85), .B(n396), .Z(n719) );
  NAND2_X1 U448 ( .A1(G227), .A2(n724), .ZN(n382) );
  INV_X1 U449 ( .A(KEYINPUT71), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n381), .B(G110), .ZN(n422) );
  XOR2_X1 U451 ( .A(KEYINPUT86), .B(G101), .Z(n384) );
  XNOR2_X1 U452 ( .A(G104), .B(G107), .ZN(n383) );
  XNOR2_X1 U453 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n695) );
  INV_X1 U455 ( .A(G469), .ZN(n389) );
  XNOR2_X2 U456 ( .A(n561), .B(KEYINPUT1), .ZN(n480) );
  XOR2_X1 U457 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n392) );
  XNOR2_X1 U458 ( .A(G128), .B(KEYINPUT87), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U460 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n393) );
  XNOR2_X1 U461 ( .A(G146), .B(G125), .ZN(n418) );
  XNOR2_X1 U462 ( .A(n393), .B(n418), .ZN(n721) );
  XNOR2_X1 U463 ( .A(n394), .B(n721), .ZN(n399) );
  XOR2_X1 U464 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n395) );
  XNOR2_X1 U465 ( .A(G119), .B(G110), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n402) );
  NAND2_X1 U467 ( .A1(n724), .A2(G234), .ZN(n401) );
  XNOR2_X1 U468 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n467) );
  XNOR2_X1 U470 ( .A(G902), .B(KEYINPUT15), .ZN(n512) );
  NAND2_X1 U471 ( .A1(n512), .A2(G234), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n403), .B(KEYINPUT20), .ZN(n407) );
  NAND2_X1 U473 ( .A1(n407), .A2(G217), .ZN(n404) );
  AND2_X1 U474 ( .A1(n407), .A2(G221), .ZN(n409) );
  INV_X1 U475 ( .A(KEYINPUT21), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n477) );
  NOR2_X1 U477 ( .A1(n513), .A2(n477), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n410), .B(KEYINPUT66), .ZN(n669) );
  NAND2_X1 U479 ( .A1(n480), .A2(n669), .ZN(n497) );
  XNOR2_X1 U480 ( .A(KEYINPUT102), .B(KEYINPUT33), .ZN(n411) );
  XNOR2_X1 U481 ( .A(n412), .B(n411), .ZN(n651) );
  XNOR2_X1 U482 ( .A(n448), .B(KEYINPUT16), .ZN(n414) );
  INV_X1 U483 ( .A(G116), .ZN(n413) );
  XNOR2_X1 U484 ( .A(n413), .B(G107), .ZN(n462) );
  XNOR2_X1 U485 ( .A(n414), .B(n462), .ZN(n415) );
  XNOR2_X1 U486 ( .A(n416), .B(n415), .ZN(n709) );
  XNOR2_X1 U487 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n417) );
  XNOR2_X1 U488 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n420), .B(n419), .ZN(n425) );
  NAND2_X1 U490 ( .A1(n724), .A2(G224), .ZN(n421) );
  XNOR2_X1 U491 ( .A(n421), .B(KEYINPUT4), .ZN(n423) );
  XNOR2_X1 U492 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U493 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n709), .B(n426), .ZN(n618) );
  INV_X1 U495 ( .A(n512), .ZN(n590) );
  OR2_X2 U496 ( .A1(n618), .A2(n590), .ZN(n431) );
  INV_X1 U497 ( .A(G902), .ZN(n428) );
  INV_X1 U498 ( .A(G237), .ZN(n427) );
  NAND2_X1 U499 ( .A1(n428), .A2(n427), .ZN(n432) );
  NAND2_X1 U500 ( .A1(n432), .A2(G210), .ZN(n429) );
  XNOR2_X1 U501 ( .A(n429), .B(KEYINPUT82), .ZN(n430) );
  XNOR2_X2 U502 ( .A(n431), .B(n430), .ZN(n554) );
  NAND2_X1 U503 ( .A1(n432), .A2(G214), .ZN(n653) );
  INV_X1 U504 ( .A(n653), .ZN(n563) );
  OR2_X2 U505 ( .A1(n554), .A2(n563), .ZN(n433) );
  XNOR2_X2 U506 ( .A(n433), .B(KEYINPUT19), .ZN(n523) );
  NAND2_X1 U507 ( .A1(G234), .A2(G237), .ZN(n434) );
  XNOR2_X1 U508 ( .A(n434), .B(KEYINPUT14), .ZN(n439) );
  NAND2_X1 U509 ( .A1(G902), .A2(n439), .ZN(n435) );
  XNOR2_X1 U510 ( .A(KEYINPUT83), .B(n435), .ZN(n436) );
  NAND2_X1 U511 ( .A1(n436), .A2(G953), .ZN(n514) );
  NOR2_X1 U512 ( .A1(G898), .A2(n514), .ZN(n438) );
  INV_X1 U513 ( .A(KEYINPUT84), .ZN(n437) );
  XNOR2_X1 U514 ( .A(n438), .B(n437), .ZN(n441) );
  NAND2_X1 U515 ( .A1(n439), .A2(G952), .ZN(n684) );
  NOR2_X1 U516 ( .A1(n684), .A2(G953), .ZN(n517) );
  INV_X1 U517 ( .A(n517), .ZN(n440) );
  NAND2_X1 U518 ( .A1(n441), .A2(n440), .ZN(n442) );
  NAND2_X1 U519 ( .A1(n523), .A2(n442), .ZN(n443) );
  XNOR2_X2 U520 ( .A(n443), .B(KEYINPUT0), .ZN(n498) );
  NOR2_X1 U521 ( .A1(n651), .A2(n498), .ZN(n445) );
  XNOR2_X1 U522 ( .A(n445), .B(n444), .ZN(n473) );
  XNOR2_X1 U523 ( .A(n446), .B(G113), .ZN(n447) );
  XNOR2_X1 U524 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U525 ( .A(n721), .B(n449), .ZN(n458) );
  XOR2_X1 U526 ( .A(KEYINPUT11), .B(KEYINPUT93), .Z(n452) );
  NAND2_X1 U527 ( .A1(n450), .A2(G214), .ZN(n451) );
  XNOR2_X1 U528 ( .A(n452), .B(n451), .ZN(n456) );
  XOR2_X1 U529 ( .A(KEYINPUT12), .B(KEYINPUT92), .Z(n454) );
  XNOR2_X1 U530 ( .A(G131), .B(G140), .ZN(n453) );
  XNOR2_X1 U531 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U532 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U533 ( .A(n458), .B(n457), .ZN(n611) );
  NOR2_X1 U534 ( .A1(G902), .A2(n611), .ZN(n459) );
  INV_X1 U535 ( .A(KEYINPUT13), .ZN(n460) );
  XNOR2_X1 U536 ( .A(n356), .B(n460), .ZN(n504) );
  XNOR2_X1 U537 ( .A(G122), .B(KEYINPUT9), .ZN(n461) );
  XNOR2_X1 U538 ( .A(n462), .B(n461), .ZN(n466) );
  XOR2_X1 U539 ( .A(KEYINPUT7), .B(KEYINPUT96), .Z(n464) );
  XNOR2_X1 U540 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n463) );
  XNOR2_X1 U541 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U542 ( .A(n466), .B(n465), .Z(n469) );
  NAND2_X1 U543 ( .A1(G217), .A2(n467), .ZN(n468) );
  XNOR2_X1 U544 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U545 ( .A(n471), .B(n470), .ZN(n701) );
  NOR2_X1 U546 ( .A1(n701), .A2(G902), .ZN(n472) );
  XNOR2_X1 U547 ( .A(G478), .B(n472), .ZN(n503) );
  INV_X1 U548 ( .A(n503), .ZN(n476) );
  NAND2_X1 U549 ( .A1(n504), .A2(n476), .ZN(n537) );
  NOR2_X2 U550 ( .A1(n473), .A2(n537), .ZN(n475) );
  NOR2_X1 U551 ( .A1(n504), .A2(n476), .ZN(n566) );
  INV_X1 U552 ( .A(n477), .ZN(n664) );
  NAND2_X1 U553 ( .A1(n566), .A2(n664), .ZN(n478) );
  OR2_X2 U554 ( .A1(n498), .A2(n478), .ZN(n479) );
  XNOR2_X1 U555 ( .A(n479), .B(KEYINPUT22), .ZN(n485) );
  NOR2_X1 U556 ( .A1(n485), .A2(n480), .ZN(n481) );
  XNOR2_X1 U557 ( .A(n481), .B(KEYINPUT101), .ZN(n483) );
  INV_X1 U558 ( .A(n532), .ZN(n668) );
  INV_X1 U559 ( .A(n513), .ZN(n665) );
  NAND2_X1 U560 ( .A1(n668), .A2(n491), .ZN(n482) );
  NOR2_X1 U561 ( .A1(n483), .A2(n482), .ZN(n605) );
  NOR2_X1 U562 ( .A1(n735), .A2(n605), .ZN(n489) );
  INV_X1 U563 ( .A(n484), .ZN(n542) );
  NOR2_X1 U564 ( .A1(n485), .A2(n542), .ZN(n493) );
  INV_X1 U565 ( .A(n480), .ZN(n579) );
  NOR2_X1 U566 ( .A1(n579), .A2(n665), .ZN(n486) );
  NAND2_X1 U567 ( .A1(n493), .A2(n486), .ZN(n488) );
  XNOR2_X1 U568 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n487) );
  XNOR2_X1 U569 ( .A(n488), .B(n487), .ZN(n608) );
  NAND2_X1 U570 ( .A1(n489), .A2(n608), .ZN(n490) );
  XNOR2_X1 U571 ( .A(n490), .B(KEYINPUT44), .ZN(n510) );
  NOR2_X1 U572 ( .A1(n480), .A2(n491), .ZN(n492) );
  NAND2_X1 U573 ( .A1(n493), .A2(n492), .ZN(n494) );
  XOR2_X1 U574 ( .A(KEYINPUT99), .B(n494), .Z(n607) );
  NAND2_X1 U575 ( .A1(n530), .A2(n668), .ZN(n495) );
  NOR2_X1 U576 ( .A1(n495), .A2(n498), .ZN(n496) );
  XOR2_X1 U577 ( .A(KEYINPUT90), .B(n496), .Z(n624) );
  NOR2_X1 U578 ( .A1(n668), .A2(n497), .ZN(n675) );
  INV_X1 U579 ( .A(n498), .ZN(n499) );
  NAND2_X1 U580 ( .A1(n675), .A2(n499), .ZN(n501) );
  XNOR2_X1 U581 ( .A(KEYINPUT91), .B(KEYINPUT31), .ZN(n500) );
  XNOR2_X1 U582 ( .A(n501), .B(n500), .ZN(n637) );
  NAND2_X1 U583 ( .A1(n624), .A2(n637), .ZN(n506) );
  NAND2_X1 U584 ( .A1(n504), .A2(n503), .ZN(n502) );
  XNOR2_X2 U585 ( .A(KEYINPUT97), .B(n502), .ZN(n631) );
  NOR2_X1 U586 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U587 ( .A(n505), .B(KEYINPUT98), .ZN(n628) );
  NOR2_X1 U588 ( .A1(n631), .A2(n628), .ZN(n658) );
  XOR2_X1 U589 ( .A(KEYINPUT76), .B(n658), .Z(n526) );
  NAND2_X1 U590 ( .A1(n506), .A2(n526), .ZN(n507) );
  NAND2_X1 U591 ( .A1(n607), .A2(n507), .ZN(n508) );
  XNOR2_X1 U592 ( .A(n508), .B(KEYINPUT100), .ZN(n509) );
  NOR2_X1 U593 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U594 ( .A(n511), .B(KEYINPUT45), .ZN(n595) );
  OR2_X1 U595 ( .A1(n595), .A2(n512), .ZN(n587) );
  NAND2_X1 U596 ( .A1(n513), .A2(n664), .ZN(n544) );
  NOR2_X1 U597 ( .A1(G900), .A2(n514), .ZN(n515) );
  XOR2_X1 U598 ( .A(KEYINPUT103), .B(n515), .Z(n516) );
  NOR2_X1 U599 ( .A1(n517), .A2(n516), .ZN(n547) );
  OR2_X2 U600 ( .A1(n544), .A2(n519), .ZN(n520) );
  XNOR2_X1 U601 ( .A(n520), .B(KEYINPUT106), .ZN(n522) );
  INV_X1 U602 ( .A(KEYINPUT28), .ZN(n521) );
  INV_X1 U603 ( .A(KEYINPUT47), .ZN(n525) );
  NOR2_X1 U604 ( .A1(n632), .A2(n525), .ZN(n524) );
  XNOR2_X1 U605 ( .A(n524), .B(KEYINPUT75), .ZN(n529) );
  AND2_X1 U606 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U607 ( .A1(n632), .A2(n527), .ZN(n528) );
  NAND2_X1 U608 ( .A1(n529), .A2(n528), .ZN(n540) );
  NAND2_X1 U609 ( .A1(n658), .A2(KEYINPUT47), .ZN(n538) );
  INV_X1 U610 ( .A(n531), .ZN(n536) );
  NAND2_X1 U611 ( .A1(n532), .A2(n653), .ZN(n533) );
  XNOR2_X1 U612 ( .A(KEYINPUT30), .B(n533), .ZN(n534) );
  NOR2_X1 U613 ( .A1(n547), .A2(n534), .ZN(n535) );
  NAND2_X1 U614 ( .A1(n536), .A2(n535), .ZN(n555) );
  OR2_X1 U615 ( .A1(n554), .A2(n361), .ZN(n610) );
  NAND2_X1 U616 ( .A1(n538), .A2(n610), .ZN(n539) );
  XNOR2_X1 U617 ( .A(n541), .B(KEYINPUT72), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n631), .A2(n542), .ZN(n543) );
  NOR2_X1 U619 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U620 ( .A1(n545), .A2(n653), .ZN(n546) );
  INV_X1 U621 ( .A(n554), .ZN(n581) );
  NAND2_X1 U622 ( .A1(n578), .A2(n581), .ZN(n549) );
  XOR2_X1 U623 ( .A(KEYINPUT36), .B(KEYINPUT80), .Z(n548) );
  XNOR2_X1 U624 ( .A(n549), .B(n548), .ZN(n550) );
  NAND2_X1 U625 ( .A1(n550), .A2(n480), .ZN(n551) );
  XNOR2_X1 U626 ( .A(n551), .B(KEYINPUT112), .ZN(n738) );
  AND2_X1 U627 ( .A1(n552), .A2(n738), .ZN(n576) );
  INV_X1 U628 ( .A(KEYINPUT38), .ZN(n553) );
  XNOR2_X1 U629 ( .A(n554), .B(n553), .ZN(n652) );
  XNOR2_X1 U630 ( .A(KEYINPUT79), .B(KEYINPUT39), .ZN(n556) );
  XNOR2_X1 U631 ( .A(n557), .B(n556), .ZN(n584) );
  NAND2_X1 U632 ( .A1(n584), .A2(n631), .ZN(n560) );
  XOR2_X1 U633 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n558) );
  XNOR2_X1 U634 ( .A(n558), .B(KEYINPUT107), .ZN(n559) );
  XNOR2_X1 U635 ( .A(n560), .B(n559), .ZN(n734) );
  AND2_X1 U636 ( .A1(n562), .A2(n357), .ZN(n569) );
  OR2_X1 U637 ( .A1(n652), .A2(n563), .ZN(n565) );
  INV_X1 U638 ( .A(KEYINPUT109), .ZN(n564) );
  XNOR2_X1 U639 ( .A(n565), .B(n564), .ZN(n657) );
  INV_X1 U640 ( .A(n566), .ZN(n655) );
  OR2_X1 U641 ( .A1(n657), .A2(n655), .ZN(n568) );
  XNOR2_X1 U642 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n567) );
  XNOR2_X1 U643 ( .A(n568), .B(n567), .ZN(n677) );
  NAND2_X1 U644 ( .A1(n569), .A2(n677), .ZN(n572) );
  INV_X1 U645 ( .A(KEYINPUT111), .ZN(n570) );
  XNOR2_X1 U646 ( .A(n570), .B(KEYINPUT42), .ZN(n571) );
  XNOR2_X1 U647 ( .A(n572), .B(n571), .ZN(n609) );
  NAND2_X1 U648 ( .A1(n734), .A2(n609), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U651 ( .A(KEYINPUT43), .B(n580), .Z(n582) );
  XNOR2_X1 U652 ( .A(n583), .B(KEYINPUT104), .ZN(n737) );
  INV_X1 U653 ( .A(n737), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n584), .A2(n628), .ZN(n640) );
  NOR2_X1 U655 ( .A1(n587), .A2(n723), .ZN(n594) );
  NAND2_X1 U656 ( .A1(n590), .A2(KEYINPUT2), .ZN(n588) );
  AND2_X1 U657 ( .A1(n588), .A2(KEYINPUT65), .ZN(n592) );
  INV_X1 U658 ( .A(KEYINPUT2), .ZN(n641) );
  NOR2_X1 U659 ( .A1(n641), .A2(KEYINPUT65), .ZN(n589) );
  AND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n591) );
  OR2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  OR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n597) );
  INV_X1 U663 ( .A(n595), .ZN(n643) );
  NOR2_X1 U664 ( .A1(n723), .A2(n641), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n643), .A2(n596), .ZN(n649) );
  AND2_X2 U666 ( .A1(n597), .A2(n649), .ZN(n694) );
  XNOR2_X1 U667 ( .A(n598), .B(KEYINPUT62), .ZN(n599) );
  INV_X1 U668 ( .A(G952), .ZN(n601) );
  NOR2_X2 U669 ( .A1(n602), .A2(n708), .ZN(n604) );
  INV_X1 U670 ( .A(KEYINPUT63), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n604), .B(n603), .ZN(G57) );
  XOR2_X1 U672 ( .A(n605), .B(G110), .Z(G12) );
  XNOR2_X1 U673 ( .A(G101), .B(KEYINPUT114), .ZN(n606) );
  XNOR2_X1 U674 ( .A(n607), .B(n606), .ZN(G3) );
  XNOR2_X1 U675 ( .A(n608), .B(G119), .ZN(G21) );
  XNOR2_X1 U676 ( .A(n609), .B(G137), .ZN(G39) );
  XNOR2_X1 U677 ( .A(n610), .B(G143), .ZN(G45) );
  NAND2_X1 U678 ( .A1(n694), .A2(G475), .ZN(n613) );
  XOR2_X1 U679 ( .A(KEYINPUT59), .B(n611), .Z(n612) );
  XNOR2_X1 U680 ( .A(n613), .B(n612), .ZN(n614) );
  NOR2_X2 U681 ( .A1(n614), .A2(n708), .ZN(n616) );
  XNOR2_X1 U682 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n615) );
  XNOR2_X1 U683 ( .A(n616), .B(n615), .ZN(G60) );
  NAND2_X1 U684 ( .A1(n694), .A2(G210), .ZN(n620) );
  XOR2_X1 U685 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n617) );
  XNOR2_X1 U686 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U687 ( .A(n620), .B(n619), .ZN(n621) );
  NOR2_X2 U688 ( .A1(n621), .A2(n708), .ZN(n622) );
  XNOR2_X1 U689 ( .A(n622), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U690 ( .A(n631), .ZN(n634) );
  NOR2_X1 U691 ( .A1(n624), .A2(n634), .ZN(n623) );
  XOR2_X1 U692 ( .A(G104), .B(n623), .Z(G6) );
  XNOR2_X1 U693 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n626) );
  INV_X1 U694 ( .A(n628), .ZN(n638) );
  NOR2_X1 U695 ( .A1(n638), .A2(n624), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U697 ( .A(G107), .B(n627), .ZN(G9) );
  XOR2_X1 U698 ( .A(G128), .B(KEYINPUT29), .Z(n630) );
  NAND2_X1 U699 ( .A1(n632), .A2(n628), .ZN(n629) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(G30) );
  NAND2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n633), .B(G146), .ZN(G48) );
  NOR2_X1 U703 ( .A1(n634), .A2(n637), .ZN(n636) );
  XNOR2_X1 U704 ( .A(G113), .B(KEYINPUT115), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(G15) );
  NOR2_X1 U706 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U707 ( .A(G116), .B(n639), .Z(G18) );
  XNOR2_X1 U708 ( .A(G134), .B(n640), .ZN(G36) );
  XNOR2_X1 U709 ( .A(n642), .B(KEYINPUT78), .ZN(n647) );
  INV_X1 U710 ( .A(KEYINPUT77), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X1 U712 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U713 ( .A(n648), .B(KEYINPUT74), .ZN(n650) );
  AND2_X2 U714 ( .A1(n650), .A2(n649), .ZN(n691) );
  BUF_X1 U715 ( .A(n651), .Z(n686) );
  INV_X1 U716 ( .A(n652), .ZN(n654) );
  NOR2_X1 U717 ( .A1(n654), .A2(n653), .ZN(n656) );
  NOR2_X1 U718 ( .A1(n656), .A2(n655), .ZN(n661) );
  NOR2_X1 U719 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U720 ( .A(n659), .B(KEYINPUT118), .ZN(n660) );
  NOR2_X1 U721 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U722 ( .A(KEYINPUT119), .B(n662), .Z(n663) );
  NOR2_X1 U723 ( .A1(n686), .A2(n663), .ZN(n681) );
  NOR2_X1 U724 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U725 ( .A(n666), .B(KEYINPUT49), .ZN(n667) );
  NAND2_X1 U726 ( .A1(n668), .A2(n667), .ZN(n672) );
  NOR2_X1 U727 ( .A1(n480), .A2(n669), .ZN(n670) );
  XNOR2_X1 U728 ( .A(n670), .B(KEYINPUT50), .ZN(n671) );
  NOR2_X1 U729 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U730 ( .A(n673), .B(KEYINPUT116), .ZN(n674) );
  NOR2_X1 U731 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U732 ( .A(KEYINPUT51), .B(n676), .Z(n678) );
  INV_X1 U733 ( .A(n677), .ZN(n685) );
  NOR2_X1 U734 ( .A1(n678), .A2(n685), .ZN(n679) );
  XOR2_X1 U735 ( .A(n679), .B(KEYINPUT117), .Z(n680) );
  NOR2_X1 U736 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U737 ( .A(n682), .B(KEYINPUT52), .ZN(n683) );
  NOR2_X1 U738 ( .A1(n684), .A2(n683), .ZN(n688) );
  NOR2_X1 U739 ( .A1(n686), .A2(n685), .ZN(n687) );
  OR2_X1 U740 ( .A1(n688), .A2(n687), .ZN(n689) );
  OR2_X1 U741 ( .A1(G953), .A2(n689), .ZN(n690) );
  NOR2_X2 U742 ( .A1(n691), .A2(n690), .ZN(n693) );
  XNOR2_X1 U743 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n692) );
  XNOR2_X1 U744 ( .A(n693), .B(n692), .ZN(G75) );
  NAND2_X1 U745 ( .A1(n704), .A2(G469), .ZN(n699) );
  XNOR2_X1 U746 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n697) );
  XNOR2_X1 U747 ( .A(n695), .B(KEYINPUT57), .ZN(n696) );
  XNOR2_X1 U748 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U749 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U750 ( .A1(n708), .A2(n700), .ZN(G54) );
  NAND2_X1 U751 ( .A1(n704), .A2(G478), .ZN(n702) );
  XNOR2_X1 U752 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U753 ( .A1(n708), .A2(n703), .ZN(G63) );
  NAND2_X1 U754 ( .A1(n704), .A2(G217), .ZN(n706) );
  XNOR2_X1 U755 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U756 ( .A1(n708), .A2(n707), .ZN(G66) );
  XOR2_X1 U757 ( .A(G110), .B(n709), .Z(n711) );
  NOR2_X1 U758 ( .A1(G898), .A2(n724), .ZN(n710) );
  NOR2_X1 U759 ( .A1(n711), .A2(n710), .ZN(n718) );
  NAND2_X1 U760 ( .A1(n643), .A2(n724), .ZN(n716) );
  XOR2_X1 U761 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n713) );
  NAND2_X1 U762 ( .A1(G224), .A2(G953), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U764 ( .A1(n714), .A2(G898), .ZN(n715) );
  NAND2_X1 U765 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U766 ( .A(n718), .B(n717), .ZN(G69) );
  XOR2_X1 U767 ( .A(n720), .B(n719), .Z(n722) );
  XNOR2_X1 U768 ( .A(n722), .B(n721), .ZN(n726) );
  XNOR2_X1 U769 ( .A(n723), .B(n726), .ZN(n725) );
  NAND2_X1 U770 ( .A1(n725), .A2(n724), .ZN(n732) );
  XNOR2_X1 U771 ( .A(KEYINPUT124), .B(n726), .ZN(n727) );
  XNOR2_X1 U772 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U773 ( .A1(G900), .A2(n728), .ZN(n729) );
  NAND2_X1 U774 ( .A1(G953), .A2(n729), .ZN(n730) );
  XOR2_X1 U775 ( .A(KEYINPUT125), .B(n730), .Z(n731) );
  NAND2_X1 U776 ( .A1(n732), .A2(n731), .ZN(G72) );
  XOR2_X1 U777 ( .A(G131), .B(KEYINPUT127), .Z(n733) );
  XNOR2_X1 U778 ( .A(n734), .B(n733), .ZN(G33) );
  XOR2_X1 U779 ( .A(n735), .B(G122), .Z(n736) );
  XNOR2_X1 U780 ( .A(KEYINPUT126), .B(n736), .ZN(G24) );
  XOR2_X1 U781 ( .A(G140), .B(n737), .Z(G42) );
  XOR2_X1 U782 ( .A(G125), .B(n738), .Z(n739) );
  XNOR2_X1 U783 ( .A(KEYINPUT37), .B(n739), .ZN(G27) );
endmodule

