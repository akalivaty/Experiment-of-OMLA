//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1246, new_n1247, new_n1248, new_n1249;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  XOR2_X1   g007(.A(KEYINPUT66), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G137), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n462), .A2(G2104), .ZN(new_n468));
  OAI22_X1  g043(.A1(new_n461), .A2(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT68), .B(G2105), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n469), .A2(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n459), .A2(new_n460), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n470), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(G2105), .ZN(new_n477));
  AOI22_X1  g052(.A1(G124), .A2(new_n476), .B1(new_n477), .B2(G136), .ZN(new_n478));
  OAI221_X1 g053(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n470), .C2(G112), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g056(.A(G114), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(G126), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n459), .B2(new_n460), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G138), .B1(new_n459), .B2(new_n460), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT4), .B1(new_n488), .B2(new_n466), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n490));
  INV_X1    g065(.A(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n494), .A2(new_n470), .A3(new_n495), .A4(G138), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n487), .B1(new_n489), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(G50), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(new_n502), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(G651), .A2(new_n504), .B1(new_n508), .B2(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n499), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n511), .A2(KEYINPUT70), .A3(new_n512), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(G51), .A3(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n500), .A2(new_n501), .B1(new_n511), .B2(new_n512), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n522), .A3(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  NAND2_X1  g101(.A1(G77), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G64), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n506), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n529), .A2(G651), .B1(G90), .B2(new_n523), .ZN(new_n530));
  INV_X1    g105(.A(new_n512), .ZN(new_n531));
  NOR2_X1   g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n519), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n533), .A2(G543), .A3(new_n521), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n530), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n500), .B2(new_n501), .ZN(new_n540));
  AND2_X1   g115(.A1(G68), .A2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(G651), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n523), .A2(G81), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT71), .B(G43), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n533), .A2(new_n521), .A3(G543), .A4(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n533), .A2(new_n521), .A3(G53), .A4(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n554), .B2(KEYINPUT73), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n520), .A2(G53), .A3(new_n521), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n523), .A2(G91), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n500), .B2(new_n501), .ZN(new_n561));
  AND2_X1   g136(.A1(G78), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n520), .A2(new_n566), .A3(G53), .A4(new_n521), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n558), .A2(new_n565), .A3(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(new_n508), .A2(new_n513), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n571), .B1(new_n510), .B2(new_n503), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT74), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n574));
  NAND2_X1  g149(.A1(G166), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(G303));
  NAND2_X1  g151(.A1(new_n523), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n578));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n578), .C1(new_n534), .C2(new_n579), .ZN(G288));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n500), .B2(new_n501), .ZN(new_n582));
  AND2_X1   g157(.A1(G73), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n513), .A2(G48), .A3(G543), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n523), .A2(G86), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n506), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G85), .B2(new_n523), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n535), .A2(G47), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G301), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n502), .A2(new_n513), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n506), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n600), .A2(new_n601), .B1(new_n604), .B2(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n534), .A2(KEYINPUT75), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n520), .A2(new_n607), .A3(new_n521), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(new_n608), .A3(G54), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n605), .A2(new_n609), .A3(KEYINPUT76), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n596), .B1(new_n614), .B2(new_n595), .ZN(G284));
  AOI21_X1  g190(.A(new_n596), .B1(new_n614), .B2(new_n595), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(G299), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n614), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g201(.A1(new_n475), .A2(new_n468), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  AOI22_X1  g207(.A1(G123), .A2(new_n476), .B1(new_n477), .B2(G135), .ZN(new_n633));
  OAI221_X1 g208(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n470), .C2(G111), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND3_X1  g211(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT77), .ZN(new_n651));
  INV_X1    g226(.A(G14), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n648), .B2(new_n649), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  OR3_X1    g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  INV_X1    g237(.A(new_n656), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n657), .B(KEYINPUT17), .Z(new_n664));
  OAI211_X1 g239(.A(new_n661), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n656), .A3(new_n657), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n660), .A3(new_n663), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n630), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT79), .B(G2096), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  MUX2_X1   g262(.A(new_n687), .B(new_n686), .S(new_n679), .Z(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT80), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n690), .B(new_n691), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n698), .A2(new_n695), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n676), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(new_n696), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n695), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n701), .A2(new_n675), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G229));
  AOI22_X1  g280(.A1(G129), .A2(new_n476), .B1(new_n477), .B2(G141), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n707));
  NAND3_X1  g282(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n706), .B(new_n709), .C1(new_n710), .C2(new_n468), .ZN(new_n711));
  MUX2_X1   g286(.A(G32), .B(new_n711), .S(G29), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT27), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1996), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G27), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G164), .B2(new_n715), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT95), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G2078), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(G2078), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G5), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G171), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT94), .ZN(new_n725));
  INV_X1    g300(.A(G1961), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n722), .A2(G21), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G168), .B2(new_n722), .ZN(new_n729));
  INV_X1    g304(.A(G1966), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n722), .A2(G19), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n547), .B2(new_n722), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G1341), .Z(new_n734));
  NAND2_X1  g309(.A1(G160), .A2(G29), .ZN(new_n735));
  INV_X1    g310(.A(G34), .ZN(new_n736));
  AOI21_X1  g311(.A(G29), .B1(new_n736), .B2(KEYINPUT24), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(KEYINPUT24), .B2(new_n736), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n735), .A2(G2084), .A3(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT31), .B(G11), .Z(new_n740));
  INV_X1    g315(.A(G28), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT93), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n635), .B2(new_n715), .ZN(new_n746));
  AOI21_X1  g321(.A(G2084), .B1(new_n735), .B2(new_n738), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n739), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n715), .A2(G33), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  NAND2_X1  g326(.A1(G115), .A2(G2104), .ZN(new_n752));
  INV_X1    g327(.A(G127), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n475), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n470), .B1(new_n754), .B2(KEYINPUT90), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(KEYINPUT90), .B2(new_n754), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n477), .A2(G139), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n751), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n749), .B1(new_n758), .B2(G29), .ZN(new_n759));
  INV_X1    g334(.A(G2072), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n731), .A2(new_n734), .A3(new_n748), .A4(new_n761), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n720), .A2(new_n721), .A3(new_n727), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G29), .A2(G35), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G162), .B2(G29), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT29), .Z(new_n766));
  INV_X1    g341(.A(G2090), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n759), .A2(new_n760), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT91), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n715), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT88), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  AOI22_X1  g350(.A1(G128), .A2(new_n476), .B1(new_n477), .B2(G140), .ZN(new_n776));
  OAI221_X1 g351(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n470), .C2(G116), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AND3_X1   g353(.A1(new_n778), .A2(KEYINPUT87), .A3(G29), .ZN(new_n779));
  AOI21_X1  g354(.A(KEYINPUT87), .B1(new_n778), .B2(G29), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT89), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2067), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n722), .A2(G4), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n614), .B2(new_n722), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G1348), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(G1348), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n783), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n722), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n618), .B2(new_n722), .ZN(new_n793));
  INV_X1    g368(.A(G1956), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n763), .A2(new_n772), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G16), .A2(G23), .ZN(new_n797));
  NAND2_X1  g372(.A1(G288), .A2(KEYINPUT82), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G288), .A2(KEYINPUT82), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n797), .B1(new_n801), .B2(G16), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT33), .B(G1976), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G166), .A2(new_n722), .ZN(new_n805));
  INV_X1    g380(.A(G22), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(G16), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT83), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT83), .ZN(new_n809));
  INV_X1    g384(.A(new_n807), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n809), .B(new_n810), .C1(G166), .C2(new_n722), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G1971), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n722), .A2(G6), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G305), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT32), .B(G1981), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n808), .A2(new_n811), .A3(G1971), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n814), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n804), .A2(new_n820), .A3(KEYINPUT84), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT84), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n814), .A2(new_n818), .A3(new_n819), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n802), .A2(new_n803), .ZN(new_n824));
  INV_X1    g399(.A(new_n803), .ZN(new_n825));
  AOI211_X1 g400(.A(new_n797), .B(new_n825), .C1(new_n801), .C2(G16), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n822), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT34), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n821), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n821), .B2(new_n828), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n715), .A2(G25), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n477), .A2(G131), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT81), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n476), .A2(G119), .ZN(new_n836));
  OAI221_X1 g411(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n833), .B1(new_n840), .B2(new_n715), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT35), .B(G1991), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n841), .B(new_n843), .ZN(new_n844));
  MUX2_X1   g419(.A(G24), .B(G290), .S(G16), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G1986), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT85), .B1(new_n832), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT84), .B1(new_n804), .B2(new_n820), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n823), .A2(new_n827), .A3(new_n822), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT34), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT85), .ZN(new_n852));
  INV_X1    g427(.A(new_n847), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n831), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT86), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT36), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n832), .A2(KEYINPUT85), .A3(new_n847), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n858), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n831), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n796), .B1(new_n859), .B2(new_n864), .ZN(G311));
  INV_X1    g440(.A(new_n796), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n863), .B1(new_n862), .B2(new_n831), .ZN(new_n867));
  AOI211_X1 g442(.A(new_n830), .B(new_n858), .C1(new_n860), .C2(new_n861), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(G150));
  INV_X1    g444(.A(G67), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n500), .B2(new_n501), .ZN(new_n871));
  AND2_X1   g446(.A1(G80), .A2(G543), .ZN(new_n872));
  OAI21_X1  g447(.A(G651), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n523), .A2(G93), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n533), .A2(new_n521), .A3(G55), .A4(G543), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(G860), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT98), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n614), .A2(G559), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT38), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n546), .A2(new_n876), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n546), .A2(new_n876), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n881), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT39), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT97), .Z(new_n887));
  INV_X1    g462(.A(G860), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n885), .B2(KEYINPUT39), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n879), .B1(new_n887), .B2(new_n889), .ZN(G145));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n778), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n758), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n839), .B(new_n628), .Z(new_n894));
  AND2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n487), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n488), .A2(new_n466), .A3(KEYINPUT4), .ZN(new_n897));
  INV_X1    g472(.A(G138), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(new_n492), .B2(new_n493), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n495), .B1(new_n899), .B2(new_n470), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n896), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n711), .B(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n477), .A2(G142), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT101), .ZN(new_n904));
  INV_X1    g479(.A(G118), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  OAI21_X1  g481(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n466), .A2(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n476), .B2(G130), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n476), .A2(new_n910), .A3(G130), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n904), .B(new_n909), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n902), .B(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n893), .A2(new_n894), .ZN(new_n916));
  OR3_X1    g491(.A1(new_n895), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n915), .B1(new_n895), .B2(new_n916), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(G160), .B(KEYINPUT99), .Z(new_n920));
  XNOR2_X1  g495(.A(G162), .B(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n921), .B(new_n635), .Z(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  INV_X1    g499(.A(new_n922), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n917), .A2(new_n925), .A3(new_n918), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g503(.A1(new_n623), .A2(new_n884), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n614), .B(new_n621), .C1(new_n882), .C2(new_n883), .ZN(new_n930));
  NAND3_X1  g505(.A1(G299), .A2(new_n609), .A3(new_n605), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n555), .A2(new_n557), .B1(new_n567), .B2(new_n568), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n610), .A2(new_n932), .A3(new_n565), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT41), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n929), .A2(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(KEYINPUT104), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n931), .A2(new_n933), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n929), .A2(new_n930), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n943), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n940), .B1(new_n945), .B2(new_n937), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(G290), .B(G166), .ZN(new_n948));
  INV_X1    g523(.A(new_n800), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n949), .A2(G305), .A3(new_n798), .ZN(new_n950));
  AOI21_X1  g525(.A(G305), .B1(new_n949), .B2(new_n798), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n801), .A2(G305), .ZN(new_n953));
  XNOR2_X1  g528(.A(G290), .B(new_n572), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n587), .B(new_n586), .C1(new_n799), .C2(new_n800), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(KEYINPUT104), .B2(new_n939), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n947), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n944), .A2(new_n959), .A3(new_n946), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(G868), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n876), .A2(new_n595), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(G295));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n967), .A3(new_n965), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n595), .B1(new_n961), .B2(new_n962), .ZN(new_n969));
  INV_X1    g544(.A(new_n965), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT105), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(G331));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n931), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n518), .A2(new_n522), .A3(KEYINPUT106), .A4(new_n524), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n882), .B2(new_n883), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n543), .A2(new_n542), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n874), .A2(new_n873), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n545), .A4(new_n875), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n546), .A2(new_n876), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n981), .A3(new_n975), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n983));
  AOI22_X1  g558(.A1(G286), .A2(new_n983), .B1(new_n530), .B2(new_n536), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n977), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n977), .B2(new_n982), .ZN(new_n986));
  OAI22_X1  g561(.A1(new_n974), .A2(new_n934), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n986), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n977), .A2(new_n982), .A3(new_n984), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n942), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n990), .A3(new_n957), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT107), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n987), .A2(new_n990), .A3(new_n993), .A4(new_n957), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n992), .A2(new_n924), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n934), .A2(KEYINPUT109), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n936), .B1(new_n934), .B2(KEYINPUT109), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n996), .A2(new_n997), .B1(new_n985), .B2(new_n986), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n957), .B1(new_n998), .B2(new_n990), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n973), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n987), .A2(new_n990), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n958), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n992), .A2(new_n1003), .A3(new_n924), .A4(new_n994), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT44), .B1(new_n1004), .B2(KEYINPUT43), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT110), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n992), .A2(new_n924), .A3(new_n994), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT43), .B1(new_n1007), .B2(new_n999), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n994), .A2(new_n924), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(new_n973), .A3(new_n992), .A4(new_n1003), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1008), .A2(new_n1009), .A3(KEYINPUT44), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1004), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n995), .A2(new_n973), .A3(new_n1000), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1013), .A2(new_n1021), .ZN(G397));
  INV_X1    g597(.A(G125), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n492), .B2(new_n493), .ZN(new_n1024));
  INV_X1    g599(.A(new_n472), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n466), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n468), .A2(new_n467), .ZN(new_n1027));
  INV_X1    g602(.A(G137), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n492), .B2(new_n493), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1027), .B1(new_n1029), .B2(new_n470), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1030), .A3(G40), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1026), .A2(new_n1030), .A3(KEYINPUT111), .A4(G40), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(G164), .B2(G1384), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n840), .A2(new_n842), .ZN(new_n1039));
  INV_X1    g614(.A(G1996), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n711), .B(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n778), .A2(G2067), .ZN(new_n1042));
  INV_X1    g617(.A(G2067), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n776), .A2(new_n1043), .A3(new_n777), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n839), .A2(new_n843), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1039), .A2(new_n1041), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G290), .A2(G1986), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1035), .B(new_n1037), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G290), .A2(G1986), .ZN(new_n1052));
  OR3_X1    g627(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1038), .A2(new_n1047), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT126), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G286), .A2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1384), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n901), .A2(KEYINPUT45), .A3(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1060), .A2(new_n1037), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n730), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT111), .B1(G160), .B2(G40), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1034), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2084), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n901), .A2(new_n1068), .A3(new_n1059), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1062), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1058), .B1(new_n1071), .B2(G8), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT45), .B1(new_n901), .B2(new_n1059), .ZN(new_n1073));
  NOR3_X1   g648(.A1(G164), .A2(new_n1036), .A3(G1384), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1966), .B1(new_n1075), .B2(new_n1065), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1069), .A2(new_n1067), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(G2084), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT125), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT125), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1062), .A2(new_n1070), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(G168), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1072), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1056), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1085), .A2(KEYINPUT62), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n801), .A2(G1976), .ZN(new_n1088));
  INV_X1    g663(.A(G1976), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(G288), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n489), .A2(new_n496), .ZN(new_n1091));
  AOI21_X1  g666(.A(G1384), .B1(new_n1091), .B2(new_n896), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1033), .A2(new_n1092), .A3(new_n1034), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1093), .A2(KEYINPUT114), .A3(G8), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT114), .B1(new_n1093), .B2(G8), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1088), .B(new_n1090), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT115), .B(G86), .Z(new_n1097));
  NAND2_X1  g672(.A1(new_n523), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(new_n584), .A3(new_n585), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(G1981), .ZN(new_n1100));
  INV_X1    g675(.A(G1981), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n587), .A2(new_n584), .A3(new_n1101), .A4(new_n585), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT116), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(KEYINPUT49), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT49), .ZN(new_n1105));
  AOI211_X1 g680(.A(KEYINPUT116), .B(new_n1105), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1094), .A2(new_n1095), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1096), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1093), .A2(G8), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1093), .A2(KEYINPUT114), .A3(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1109), .B1(new_n1114), .B2(new_n1088), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1068), .B1(new_n901), .B2(new_n1059), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1035), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1067), .A2(KEYINPUT118), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n767), .A3(new_n1069), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1061), .A2(new_n813), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(G8), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n573), .A2(G8), .A3(new_n575), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT55), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1122), .B1(G2090), .B2(new_n1077), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT113), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1122), .B(KEYINPUT113), .C1(G2090), .C2(new_n1077), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(G8), .A3(new_n1127), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1061), .B2(G2078), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1077), .A2(new_n726), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1135), .A2(G2078), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1136), .B(new_n1137), .C1(new_n1061), .C2(new_n1138), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1139), .A2(G171), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1116), .A2(new_n1129), .A3(new_n1134), .A4(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1055), .B1(new_n1087), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1141), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1086), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1062), .A2(new_n1070), .A3(new_n1080), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1080), .B1(new_n1062), .B2(new_n1070), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1083), .B1(new_n1148), .B2(G168), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1144), .B(new_n1145), .C1(new_n1149), .C2(new_n1072), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1143), .A2(new_n1150), .A3(KEYINPUT126), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1145), .B1(new_n1149), .B2(new_n1072), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT62), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1142), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(G8), .B(G168), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT119), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1071), .A2(new_n1157), .A3(G8), .A4(G168), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1159), .A2(new_n1116), .A3(new_n1129), .A4(new_n1134), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1161), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1132), .A2(G8), .A3(new_n1133), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1128), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1163), .A2(new_n1165), .A3(new_n1134), .A4(new_n1116), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1134), .A2(new_n1115), .A3(new_n1108), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1102), .B(KEYINPUT117), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1107), .ZN(new_n1170));
  OR2_X1    g745(.A1(G288), .A2(G1976), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1168), .B1(new_n1114), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n612), .B2(new_n613), .ZN(new_n1175));
  INV_X1    g750(.A(G1348), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1093), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1077), .A2(new_n1176), .B1(new_n1177), .B2(new_n1043), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n612), .A2(new_n1174), .A3(new_n613), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1175), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1077), .A2(new_n1176), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1177), .A2(new_n1043), .ZN(new_n1182));
  AND4_X1   g757(.A1(KEYINPUT60), .A2(new_n1181), .A3(new_n1182), .A4(new_n614), .ZN(new_n1183));
  XNOR2_X1  g758(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(G1341), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1093), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(new_n1061), .B2(G1996), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT59), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1187), .A2(new_n1188), .A3(new_n547), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1188), .B1(new_n1187), .B2(new_n547), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1180), .A2(new_n1183), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT57), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n559), .A2(new_n563), .A3(KEYINPUT121), .ZN(new_n1193));
  AOI21_X1  g768(.A(KEYINPUT121), .B1(new_n559), .B2(new_n563), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n932), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT120), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n932), .A2(KEYINPUT120), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1200), .B1(new_n1192), .B2(new_n618), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1120), .A2(new_n1069), .ZN(new_n1202));
  AOI21_X1  g777(.A(G1956), .B1(new_n1202), .B2(new_n1119), .ZN(new_n1203));
  XOR2_X1   g778(.A(KEYINPUT56), .B(G2072), .Z(new_n1204));
  NOR2_X1   g779(.A1(new_n1061), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1201), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1119), .A2(new_n1069), .A3(new_n1120), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1205), .B1(new_n1207), .B2(new_n794), .ZN(new_n1208));
  AOI22_X1  g783(.A1(new_n1198), .A2(new_n1199), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1191), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1201), .B1(new_n1208), .B2(KEYINPUT122), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT122), .ZN(new_n1215));
  NOR3_X1   g790(.A1(new_n1203), .A2(new_n1215), .A3(new_n1205), .ZN(new_n1216));
  OAI211_X1 g791(.A(KEYINPUT61), .B(new_n1210), .C1(new_n1214), .C2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n614), .ZN(new_n1218));
  OAI22_X1  g793(.A1(new_n1214), .A2(new_n1216), .B1(new_n1218), .B2(new_n1178), .ZN(new_n1219));
  AOI22_X1  g794(.A1(new_n1213), .A2(new_n1217), .B1(new_n1210), .B2(new_n1219), .ZN(new_n1220));
  AND3_X1   g795(.A1(new_n1116), .A2(new_n1129), .A3(new_n1134), .ZN(new_n1221));
  XNOR2_X1  g796(.A(G301), .B(KEYINPUT54), .ZN(new_n1222));
  AND2_X1   g797(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n1031), .A2(new_n1138), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1222), .B1(new_n1075), .B2(new_n1224), .ZN(new_n1225));
  AOI22_X1  g800(.A1(new_n1139), .A2(new_n1222), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1152), .A2(new_n1221), .A3(new_n1226), .ZN(new_n1227));
  OAI211_X1 g802(.A(new_n1167), .B(new_n1173), .C1(new_n1220), .C2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1054), .B1(new_n1154), .B2(new_n1228), .ZN(new_n1229));
  AND2_X1   g804(.A1(new_n1038), .A2(new_n1052), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1230), .A2(KEYINPUT48), .ZN(new_n1231));
  AND2_X1   g806(.A1(new_n1230), .A2(KEYINPUT48), .ZN(new_n1232));
  AOI211_X1 g807(.A(new_n1231), .B(new_n1232), .C1(new_n1038), .C2(new_n1047), .ZN(new_n1233));
  INV_X1    g808(.A(new_n1045), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n1038), .B1(new_n1234), .B2(new_n711), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1236));
  AND2_X1   g811(.A1(new_n1236), .A2(KEYINPUT46), .ZN(new_n1237));
  NOR2_X1   g812(.A1(new_n1236), .A2(KEYINPUT46), .ZN(new_n1238));
  OAI21_X1  g813(.A(new_n1235), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  XOR2_X1   g814(.A(new_n1239), .B(KEYINPUT47), .Z(new_n1240));
  NAND2_X1  g815(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1241));
  OAI21_X1  g816(.A(new_n1044), .B1(new_n1241), .B2(new_n1039), .ZN(new_n1242));
  AOI211_X1 g817(.A(new_n1233), .B(new_n1240), .C1(new_n1038), .C2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1229), .A2(new_n1243), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g819(.A(G319), .B1(new_n672), .B2(new_n673), .ZN(new_n1246));
  OR2_X1    g820(.A1(new_n1246), .A2(KEYINPUT127), .ZN(new_n1247));
  NAND2_X1  g821(.A1(new_n1246), .A2(KEYINPUT127), .ZN(new_n1248));
  AOI22_X1  g822(.A1(new_n651), .A2(new_n653), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND4_X1  g823(.A1(new_n1019), .A2(new_n704), .A3(new_n927), .A4(new_n1249), .ZN(G225));
  INV_X1    g824(.A(G225), .ZN(G308));
endmodule


