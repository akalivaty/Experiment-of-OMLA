

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715;

  AND2_X1 U365 ( .A1(n489), .A2(n488), .ZN(n346) );
  XNOR2_X1 U366 ( .A(n426), .B(KEYINPUT4), .ZN(n460) );
  XNOR2_X1 U367 ( .A(n346), .B(n490), .ZN(n643) );
  INV_X1 U368 ( .A(G953), .ZN(n702) );
  INV_X1 U369 ( .A(n579), .ZN(n557) );
  NOR2_X2 U370 ( .A1(n686), .A2(n592), .ZN(n595) );
  NAND2_X2 U371 ( .A1(n515), .A2(n514), .ZN(n355) );
  XOR2_X2 U372 ( .A(G472), .B(n471), .Z(n649) );
  XNOR2_X2 U373 ( .A(n434), .B(n349), .ZN(n517) );
  XNOR2_X2 U374 ( .A(n386), .B(n429), .ZN(n468) );
  XOR2_X2 U375 ( .A(n557), .B(KEYINPUT38), .Z(n635) );
  NOR2_X1 U376 ( .A1(n599), .A2(n686), .ZN(n601) );
  OR2_X1 U377 ( .A1(n629), .A2(n560), .ZN(n572) );
  XNOR2_X1 U378 ( .A(n672), .B(n352), .ZN(n673) );
  XNOR2_X1 U379 ( .A(n431), .B(n343), .ZN(n405) );
  XOR2_X1 U380 ( .A(n403), .B(n402), .Z(n343) );
  XNOR2_X2 U381 ( .A(n479), .B(n478), .ZN(n520) );
  NOR2_X2 U382 ( .A1(G902), .A2(n677), .ZN(n479) );
  XOR2_X1 U383 ( .A(G146), .B(G125), .Z(n421) );
  XNOR2_X1 U384 ( .A(n460), .B(n459), .ZN(n473) );
  XNOR2_X1 U385 ( .A(n421), .B(n397), .ZN(n700) );
  XNOR2_X1 U386 ( .A(n362), .B(n361), .ZN(n360) );
  XNOR2_X1 U387 ( .A(G101), .B(G146), .ZN(n362) );
  XNOR2_X1 U388 ( .A(G107), .B(G104), .ZN(n361) );
  XOR2_X1 U389 ( .A(KEYINPUT71), .B(G110), .Z(n474) );
  NAND2_X1 U390 ( .A1(n517), .A2(n634), .ZN(n552) );
  INV_X1 U391 ( .A(G469), .ZN(n478) );
  NOR2_X1 U392 ( .A1(G902), .A2(n596), .ZN(n471) );
  XNOR2_X1 U393 ( .A(n520), .B(KEYINPUT1), .ZN(n359) );
  XOR2_X1 U394 ( .A(KEYINPUT8), .B(n413), .Z(n450) );
  INV_X1 U395 ( .A(n700), .ZN(n368) );
  XNOR2_X1 U396 ( .A(n365), .B(n451), .ZN(n364) );
  XNOR2_X1 U397 ( .A(n452), .B(n449), .ZN(n365) );
  XNOR2_X1 U398 ( .A(KEYINPUT87), .B(KEYINPUT24), .ZN(n449) );
  AND2_X1 U399 ( .A1(n344), .A2(n351), .ZN(n374) );
  AND2_X1 U400 ( .A1(n372), .A2(n358), .ZN(n371) );
  OR2_X1 U401 ( .A1(n344), .A2(n351), .ZN(n372) );
  XNOR2_X1 U402 ( .A(n448), .B(n447), .ZN(n499) );
  INV_X1 U403 ( .A(KEYINPUT22), .ZN(n447) );
  NOR2_X1 U404 ( .A1(n446), .A2(n647), .ZN(n448) );
  XNOR2_X1 U405 ( .A(n385), .B(G107), .ZN(n430) );
  INV_X1 U406 ( .A(G116), .ZN(n385) );
  XNOR2_X1 U407 ( .A(G131), .B(G143), .ZN(n398) );
  XNOR2_X1 U408 ( .A(G116), .B(G113), .ZN(n461) );
  XOR2_X1 U409 ( .A(G137), .B(G146), .Z(n462) );
  XNOR2_X1 U410 ( .A(n430), .B(KEYINPUT16), .ZN(n384) );
  XNOR2_X1 U411 ( .A(n401), .B(G122), .ZN(n431) );
  XNOR2_X1 U412 ( .A(G113), .B(G104), .ZN(n401) );
  XNOR2_X1 U413 ( .A(G119), .B(G101), .ZN(n429) );
  XNOR2_X1 U414 ( .A(n428), .B(KEYINPUT67), .ZN(n386) );
  XNOR2_X1 U415 ( .A(KEYINPUT3), .B(KEYINPUT82), .ZN(n428) );
  XOR2_X1 U416 ( .A(KEYINPUT88), .B(G110), .Z(n452) );
  INV_X1 U417 ( .A(n421), .ZN(n422) );
  XNOR2_X1 U418 ( .A(KEYINPUT83), .B(KEYINPUT72), .ZN(n420) );
  AND2_X1 U419 ( .A1(n389), .A2(n348), .ZN(n388) );
  INV_X1 U420 ( .A(n638), .ZN(n393) );
  NAND2_X1 U421 ( .A1(n387), .A2(n345), .ZN(n390) );
  AND2_X1 U422 ( .A1(n633), .A2(n583), .ZN(n584) );
  XNOR2_X1 U423 ( .A(n383), .B(n381), .ZN(n693) );
  XNOR2_X1 U424 ( .A(n431), .B(n382), .ZN(n381) );
  XNOR2_X1 U425 ( .A(n468), .B(n384), .ZN(n383) );
  INV_X1 U426 ( .A(n474), .ZN(n382) );
  XNOR2_X1 U427 ( .A(n699), .B(n477), .ZN(n677) );
  XNOR2_X1 U428 ( .A(n360), .B(n474), .ZN(n476) );
  INV_X1 U429 ( .A(KEYINPUT39), .ZN(n543) );
  NOR2_X1 U430 ( .A1(n555), .A2(n542), .ZN(n544) );
  NOR2_X1 U431 ( .A1(n643), .A2(n502), .ZN(n492) );
  XNOR2_X1 U432 ( .A(n366), .B(n364), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n453), .B(n368), .ZN(n367) );
  NAND2_X1 U434 ( .A1(n450), .A2(G221), .ZN(n366) );
  XOR2_X1 U435 ( .A(KEYINPUT81), .B(n394), .Z(n686) );
  XNOR2_X1 U436 ( .A(n535), .B(n534), .ZN(n710) );
  INV_X1 U437 ( .A(KEYINPUT42), .ZN(n534) );
  NAND2_X1 U438 ( .A1(n373), .A2(n371), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n380), .B(KEYINPUT32), .ZN(n714) );
  NOR2_X1 U440 ( .A1(n561), .A2(n562), .ZN(n620) );
  INV_X1 U441 ( .A(KEYINPUT101), .ZN(n378) );
  NAND2_X1 U442 ( .A1(n482), .A2(n480), .ZN(n379) );
  AND2_X1 U443 ( .A1(n619), .A2(n376), .ZN(n344) );
  NOR2_X1 U444 ( .A1(n442), .A2(KEYINPUT0), .ZN(n345) );
  XOR2_X1 U445 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n347) );
  AND2_X1 U446 ( .A1(n393), .A2(n392), .ZN(n348) );
  AND2_X1 U447 ( .A1(n435), .A2(G210), .ZN(n349) );
  INV_X1 U448 ( .A(n358), .ZN(n553) );
  BUF_X1 U449 ( .A(n359), .Z(n358) );
  NOR2_X1 U450 ( .A1(n539), .A2(n647), .ZN(n350) );
  INV_X1 U451 ( .A(n486), .ZN(n527) );
  XOR2_X1 U452 ( .A(KEYINPUT36), .B(KEYINPUT78), .Z(n351) );
  XNOR2_X1 U453 ( .A(n379), .B(n378), .ZN(n712) );
  XNOR2_X1 U454 ( .A(n473), .B(n472), .ZN(n699) );
  XNOR2_X1 U455 ( .A(n367), .B(n363), .ZN(n683) );
  XNOR2_X1 U456 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n352) );
  NOR2_X2 U457 ( .A1(n686), .A2(n675), .ZN(n676) );
  NAND2_X1 U458 ( .A1(n388), .A2(n390), .ZN(n446) );
  NOR2_X2 U459 ( .A1(n690), .A2(n701), .ZN(n354) );
  XNOR2_X2 U460 ( .A(n355), .B(n516), .ZN(n690) );
  NAND2_X1 U461 ( .A1(n482), .A2(n481), .ZN(n380) );
  NOR2_X1 U462 ( .A1(n602), .A2(G902), .ZN(n419) );
  XNOR2_X1 U463 ( .A(n416), .B(n417), .ZN(n602) );
  NAND2_X1 U464 ( .A1(n585), .A2(n584), .ZN(n701) );
  XNOR2_X1 U465 ( .A(n353), .B(n547), .ZN(n574) );
  NAND2_X1 U466 ( .A1(n715), .A2(n710), .ZN(n353) );
  XNOR2_X2 U467 ( .A(n354), .B(KEYINPUT2), .ZN(n666) );
  NAND2_X1 U468 ( .A1(n496), .A2(n356), .ZN(n498) );
  INV_X1 U469 ( .A(n357), .ZN(n356) );
  NAND2_X1 U470 ( .A1(n357), .A2(n483), .ZN(n497) );
  XNOR2_X1 U471 ( .A(n357), .B(G122), .ZN(n709) );
  XNOR2_X2 U472 ( .A(n495), .B(KEYINPUT35), .ZN(n357) );
  NAND2_X1 U473 ( .A1(n645), .A2(n359), .ZN(n487) );
  AND2_X1 U474 ( .A1(n553), .A2(n528), .ZN(n480) );
  NOR2_X1 U475 ( .A1(n645), .A2(n358), .ZN(n646) );
  AND2_X1 U476 ( .A1(n549), .A2(n358), .ZN(n481) );
  NOR2_X1 U477 ( .A1(n576), .A2(n358), .ZN(n577) );
  NOR2_X1 U478 ( .A1(n501), .A2(n358), .ZN(n608) );
  NOR2_X4 U479 ( .A1(n666), .A2(n586), .ZN(n671) );
  XNOR2_X1 U480 ( .A(n369), .B(KEYINPUT66), .ZN(n548) );
  NAND2_X1 U481 ( .A1(n486), .A2(n350), .ZN(n369) );
  NOR2_X1 U482 ( .A1(n375), .A2(n370), .ZN(n629) );
  NAND2_X1 U483 ( .A1(n551), .A2(n374), .ZN(n373) );
  NOR2_X1 U484 ( .A1(n551), .A2(n351), .ZN(n375) );
  NAND2_X1 U485 ( .A1(n551), .A2(n619), .ZN(n576) );
  INV_X1 U486 ( .A(n552), .ZN(n376) );
  XNOR2_X1 U487 ( .A(n377), .B(n485), .ZN(n496) );
  NAND2_X1 U488 ( .A1(n712), .A2(n714), .ZN(n377) );
  NAND2_X1 U489 ( .A1(n561), .A2(KEYINPUT0), .ZN(n389) );
  XNOR2_X2 U490 ( .A(n552), .B(n436), .ZN(n561) );
  AND2_X1 U491 ( .A1(n389), .A2(n392), .ZN(n391) );
  INV_X1 U492 ( .A(n561), .ZN(n387) );
  NAND2_X1 U493 ( .A1(n391), .A2(n390), .ZN(n505) );
  NAND2_X1 U494 ( .A1(n442), .A2(KEYINPUT0), .ZN(n392) );
  NOR2_X1 U495 ( .A1(n605), .A2(n686), .ZN(n607) );
  XNOR2_X1 U496 ( .A(n484), .B(KEYINPUT77), .ZN(n485) );
  XNOR2_X1 U497 ( .A(G131), .B(G134), .ZN(n459) );
  XNOR2_X1 U498 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U499 ( .A(n468), .B(n467), .ZN(n469) );
  BUF_X1 U500 ( .A(n643), .Z(n662) );
  XNOR2_X1 U501 ( .A(n470), .B(n469), .ZN(n596) );
  INV_X1 U502 ( .A(KEYINPUT45), .ZN(n516) );
  XNOR2_X1 U503 ( .A(n674), .B(n673), .ZN(n675) );
  INV_X1 U504 ( .A(KEYINPUT63), .ZN(n600) );
  INV_X1 U505 ( .A(KEYINPUT121), .ZN(n606) );
  XNOR2_X1 U506 ( .A(n595), .B(n594), .ZN(G60) );
  NOR2_X1 U507 ( .A1(G952), .A2(n702), .ZN(n394) );
  XOR2_X1 U508 ( .A(KEYINPUT97), .B(KEYINPUT13), .Z(n396) );
  XNOR2_X1 U509 ( .A(KEYINPUT96), .B(G475), .ZN(n395) );
  XNOR2_X1 U510 ( .A(n396), .B(n395), .ZN(n409) );
  INV_X1 U511 ( .A(KEYINPUT10), .ZN(n397) );
  XOR2_X1 U512 ( .A(KEYINPUT94), .B(G140), .Z(n399) );
  XNOR2_X1 U513 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U514 ( .A(n700), .B(n400), .ZN(n407) );
  XOR2_X1 U515 ( .A(KEYINPUT93), .B(KEYINPUT11), .Z(n403) );
  XNOR2_X1 U516 ( .A(KEYINPUT95), .B(KEYINPUT12), .ZN(n402) );
  NOR2_X1 U517 ( .A1(G953), .A2(G237), .ZN(n464) );
  NAND2_X1 U518 ( .A1(G214), .A2(n464), .ZN(n404) );
  XNOR2_X1 U519 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U520 ( .A(n407), .B(n406), .ZN(n587) );
  NOR2_X1 U521 ( .A1(G902), .A2(n587), .ZN(n408) );
  XNOR2_X1 U522 ( .A(n409), .B(n408), .ZN(n508) );
  XOR2_X1 U523 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n412) );
  XNOR2_X2 U524 ( .A(G143), .B(G128), .ZN(n426) );
  INV_X1 U525 ( .A(n426), .ZN(n410) );
  XNOR2_X1 U526 ( .A(n410), .B(n430), .ZN(n411) );
  XNOR2_X1 U527 ( .A(n412), .B(n411), .ZN(n417) );
  XOR2_X1 U528 ( .A(G122), .B(G134), .Z(n415) );
  NAND2_X1 U529 ( .A1(G234), .A2(n702), .ZN(n413) );
  NAND2_X1 U530 ( .A1(G217), .A2(n450), .ZN(n414) );
  XNOR2_X1 U531 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U532 ( .A(KEYINPUT99), .B(G478), .ZN(n418) );
  XNOR2_X1 U533 ( .A(n419), .B(n418), .ZN(n510) );
  OR2_X1 U534 ( .A1(n508), .A2(n510), .ZN(n638) );
  XNOR2_X1 U535 ( .A(n347), .B(n420), .ZN(n423) );
  XNOR2_X1 U536 ( .A(n423), .B(n422), .ZN(n425) );
  NAND2_X1 U537 ( .A1(G224), .A2(n702), .ZN(n424) );
  XNOR2_X1 U538 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U539 ( .A(n427), .B(n460), .ZN(n432) );
  XNOR2_X1 U540 ( .A(n693), .B(n432), .ZN(n672) );
  XNOR2_X1 U541 ( .A(KEYINPUT15), .B(G902), .ZN(n586) );
  NAND2_X1 U542 ( .A1(n672), .A2(n586), .ZN(n434) );
  NOR2_X1 U543 ( .A1(G237), .A2(G902), .ZN(n433) );
  XOR2_X1 U544 ( .A(KEYINPUT70), .B(n433), .Z(n435) );
  NAND2_X1 U545 ( .A1(n435), .A2(G214), .ZN(n634) );
  XNOR2_X1 U546 ( .A(KEYINPUT19), .B(KEYINPUT65), .ZN(n436) );
  NAND2_X1 U547 ( .A1(G234), .A2(G237), .ZN(n437) );
  XNOR2_X1 U548 ( .A(n437), .B(KEYINPUT14), .ZN(n439) );
  NAND2_X1 U549 ( .A1(G952), .A2(n439), .ZN(n661) );
  NOR2_X1 U550 ( .A1(G953), .A2(n661), .ZN(n525) );
  NOR2_X1 U551 ( .A1(G898), .A2(n702), .ZN(n438) );
  XOR2_X1 U552 ( .A(KEYINPUT84), .B(n438), .Z(n694) );
  NAND2_X1 U553 ( .A1(G902), .A2(n439), .ZN(n521) );
  NOR2_X1 U554 ( .A1(n694), .A2(n521), .ZN(n440) );
  XOR2_X1 U555 ( .A(KEYINPUT85), .B(n440), .Z(n441) );
  NOR2_X1 U556 ( .A1(n525), .A2(n441), .ZN(n442) );
  NAND2_X1 U557 ( .A1(n586), .A2(G234), .ZN(n444) );
  XNOR2_X1 U558 ( .A(KEYINPUT20), .B(KEYINPUT90), .ZN(n443) );
  XNOR2_X1 U559 ( .A(n444), .B(n443), .ZN(n454) );
  NAND2_X1 U560 ( .A1(n454), .A2(G221), .ZN(n445) );
  XNOR2_X1 U561 ( .A(n445), .B(KEYINPUT21), .ZN(n647) );
  XOR2_X1 U562 ( .A(G137), .B(G140), .Z(n472) );
  XNOR2_X1 U563 ( .A(n472), .B(KEYINPUT23), .ZN(n453) );
  XNOR2_X1 U564 ( .A(G119), .B(G128), .ZN(n451) );
  NOR2_X1 U565 ( .A1(G902), .A2(n683), .ZN(n458) );
  NAND2_X1 U566 ( .A1(n454), .A2(G217), .ZN(n456) );
  XNOR2_X1 U567 ( .A(KEYINPUT89), .B(KEYINPUT25), .ZN(n455) );
  XNOR2_X1 U568 ( .A(n458), .B(n457), .ZN(n486) );
  NOR2_X2 U569 ( .A1(n499), .A2(n527), .ZN(n482) );
  XNOR2_X1 U570 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U571 ( .A(n473), .B(n463), .ZN(n470) );
  XOR2_X1 U572 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n466) );
  NAND2_X1 U573 ( .A1(n464), .A2(G210), .ZN(n465) );
  XNOR2_X1 U574 ( .A(n466), .B(n465), .ZN(n467) );
  INV_X1 U575 ( .A(n649), .ZN(n528) );
  NAND2_X1 U576 ( .A1(G227), .A2(n702), .ZN(n475) );
  XNOR2_X1 U577 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U578 ( .A(n649), .B(KEYINPUT6), .ZN(n549) );
  INV_X1 U579 ( .A(KEYINPUT44), .ZN(n483) );
  NAND2_X1 U580 ( .A1(n483), .A2(KEYINPUT76), .ZN(n484) );
  XNOR2_X1 U581 ( .A(n505), .B(KEYINPUT86), .ZN(n502) );
  NOR2_X1 U582 ( .A1(n647), .A2(n486), .ZN(n645) );
  XNOR2_X1 U583 ( .A(n487), .B(KEYINPUT69), .ZN(n504) );
  XNOR2_X1 U584 ( .A(n504), .B(KEYINPUT102), .ZN(n489) );
  INV_X1 U585 ( .A(n549), .ZN(n488) );
  XOR2_X1 U586 ( .A(KEYINPUT33), .B(KEYINPUT79), .Z(n490) );
  XNOR2_X1 U587 ( .A(KEYINPUT68), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U588 ( .A(n492), .B(n491), .ZN(n494) );
  NAND2_X1 U589 ( .A1(n510), .A2(n508), .ZN(n554) );
  INV_X1 U590 ( .A(n554), .ZN(n493) );
  NAND2_X1 U591 ( .A1(n494), .A2(n493), .ZN(n495) );
  NAND2_X1 U592 ( .A1(n498), .A2(n497), .ZN(n515) );
  NOR2_X1 U593 ( .A1(n486), .A2(n499), .ZN(n500) );
  NAND2_X1 U594 ( .A1(n500), .A2(n549), .ZN(n501) );
  INV_X1 U595 ( .A(n608), .ZN(n513) );
  NAND2_X1 U596 ( .A1(n520), .A2(n645), .ZN(n536) );
  NOR2_X1 U597 ( .A1(n536), .A2(n502), .ZN(n503) );
  NAND2_X1 U598 ( .A1(n503), .A2(n528), .ZN(n610) );
  NAND2_X1 U599 ( .A1(n649), .A2(n504), .ZN(n654) );
  NOR2_X1 U600 ( .A1(n505), .A2(n654), .ZN(n506) );
  XNOR2_X1 U601 ( .A(n506), .B(KEYINPUT31), .ZN(n507) );
  XNOR2_X1 U602 ( .A(n507), .B(KEYINPUT92), .ZN(n626) );
  NAND2_X1 U603 ( .A1(n610), .A2(n626), .ZN(n511) );
  XOR2_X1 U604 ( .A(KEYINPUT98), .B(n508), .Z(n509) );
  NOR2_X1 U605 ( .A1(n510), .A2(n509), .ZN(n619) );
  NAND2_X1 U606 ( .A1(n510), .A2(n509), .ZN(n625) );
  XOR2_X1 U607 ( .A(KEYINPUT100), .B(n625), .Z(n582) );
  NOR2_X1 U608 ( .A1(n619), .A2(n582), .ZN(n640) );
  INV_X1 U609 ( .A(n640), .ZN(n564) );
  NAND2_X1 U610 ( .A1(n511), .A2(n564), .ZN(n512) );
  AND2_X1 U611 ( .A1(n513), .A2(n512), .ZN(n514) );
  XOR2_X1 U612 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n547) );
  INV_X1 U613 ( .A(n517), .ZN(n579) );
  NAND2_X1 U614 ( .A1(n635), .A2(n634), .ZN(n639) );
  NOR2_X1 U615 ( .A1(n638), .A2(n639), .ZN(n519) );
  XNOR2_X1 U616 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U617 ( .A(n519), .B(n518), .ZN(n663) );
  XNOR2_X1 U618 ( .A(n520), .B(KEYINPUT106), .ZN(n533) );
  NOR2_X1 U619 ( .A1(G900), .A2(n521), .ZN(n522) );
  NAND2_X1 U620 ( .A1(G953), .A2(n522), .ZN(n523) );
  XNOR2_X1 U621 ( .A(KEYINPUT103), .B(n523), .ZN(n524) );
  NOR2_X1 U622 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U623 ( .A(KEYINPUT73), .B(n526), .Z(n539) );
  NOR2_X1 U624 ( .A1(n548), .A2(n528), .ZN(n531) );
  XNOR2_X1 U625 ( .A(KEYINPUT28), .B(KEYINPUT107), .ZN(n529) );
  XNOR2_X1 U626 ( .A(n529), .B(KEYINPUT108), .ZN(n530) );
  XOR2_X1 U627 ( .A(n531), .B(n530), .Z(n532) );
  NAND2_X1 U628 ( .A1(n533), .A2(n532), .ZN(n562) );
  NOR2_X1 U629 ( .A1(n663), .A2(n562), .ZN(n535) );
  XOR2_X1 U630 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n546) );
  XNOR2_X1 U631 ( .A(KEYINPUT105), .B(n536), .ZN(n541) );
  NAND2_X1 U632 ( .A1(n649), .A2(n634), .ZN(n537) );
  XNOR2_X1 U633 ( .A(KEYINPUT30), .B(n537), .ZN(n538) );
  NOR2_X1 U634 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U635 ( .A1(n541), .A2(n540), .ZN(n555) );
  INV_X1 U636 ( .A(n635), .ZN(n542) );
  XNOR2_X1 U637 ( .A(n544), .B(n543), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n581), .A2(n619), .ZN(n545) );
  XNOR2_X1 U639 ( .A(n546), .B(n545), .ZN(n715) );
  NOR2_X1 U640 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U641 ( .A(n550), .B(KEYINPUT104), .ZN(n551) );
  NAND2_X1 U642 ( .A1(n640), .A2(KEYINPUT47), .ZN(n558) );
  NOR2_X1 U643 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U644 ( .A1(n557), .A2(n556), .ZN(n618) );
  NAND2_X1 U645 ( .A1(n558), .A2(n618), .ZN(n559) );
  XNOR2_X1 U646 ( .A(n559), .B(KEYINPUT74), .ZN(n560) );
  XNOR2_X1 U647 ( .A(n620), .B(KEYINPUT75), .ZN(n563) );
  NAND2_X1 U648 ( .A1(n563), .A2(KEYINPUT47), .ZN(n570) );
  INV_X1 U649 ( .A(KEYINPUT75), .ZN(n566) );
  NAND2_X1 U650 ( .A1(n620), .A2(n564), .ZN(n565) );
  NAND2_X1 U651 ( .A1(n566), .A2(n565), .ZN(n568) );
  INV_X1 U652 ( .A(KEYINPUT47), .ZN(n567) );
  NAND2_X1 U653 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U654 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U655 ( .A1(n572), .A2(n571), .ZN(n573) );
  AND2_X1 U656 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U657 ( .A(n575), .B(KEYINPUT48), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n577), .A2(n634), .ZN(n578) );
  XNOR2_X1 U659 ( .A(n578), .B(KEYINPUT43), .ZN(n580) );
  NAND2_X1 U660 ( .A1(n580), .A2(n579), .ZN(n633) );
  AND2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n632) );
  INV_X1 U662 ( .A(n632), .ZN(n583) );
  NAND2_X1 U663 ( .A1(n671), .A2(G475), .ZN(n591) );
  XOR2_X1 U664 ( .A(KEYINPUT59), .B(KEYINPUT118), .Z(n589) );
  XNOR2_X1 U665 ( .A(n587), .B(KEYINPUT80), .ZN(n588) );
  XNOR2_X1 U666 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U667 ( .A(n591), .B(n590), .ZN(n592) );
  INV_X1 U668 ( .A(KEYINPUT119), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n593), .B(KEYINPUT60), .ZN(n594) );
  XNOR2_X1 U670 ( .A(n596), .B(KEYINPUT62), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n671), .A2(G472), .ZN(n597) );
  XNOR2_X1 U672 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n601), .B(n600), .ZN(G57) );
  XNOR2_X1 U674 ( .A(n602), .B(KEYINPUT120), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G478), .A2(n671), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n607), .B(n606), .ZN(G63) );
  XOR2_X1 U678 ( .A(G101), .B(n608), .Z(G3) );
  INV_X1 U679 ( .A(n619), .ZN(n622) );
  NOR2_X1 U680 ( .A1(n622), .A2(n610), .ZN(n609) );
  XOR2_X1 U681 ( .A(G104), .B(n609), .Z(G6) );
  NOR2_X1 U682 ( .A1(n610), .A2(n625), .ZN(n614) );
  XOR2_X1 U683 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n612) );
  XNOR2_X1 U684 ( .A(G107), .B(KEYINPUT111), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n614), .B(n613), .ZN(G9) );
  INV_X1 U687 ( .A(n620), .ZN(n615) );
  NOR2_X1 U688 ( .A1(n625), .A2(n615), .ZN(n617) );
  XNOR2_X1 U689 ( .A(G128), .B(KEYINPUT29), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n617), .B(n616), .ZN(G30) );
  XNOR2_X1 U691 ( .A(G143), .B(n618), .ZN(G45) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n621), .B(G146), .ZN(G48) );
  NOR2_X1 U694 ( .A1(n626), .A2(n622), .ZN(n624) );
  XNOR2_X1 U695 ( .A(G113), .B(KEYINPUT113), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n624), .B(n623), .ZN(G15) );
  NOR2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U698 ( .A(KEYINPUT114), .B(n627), .Z(n628) );
  XNOR2_X1 U699 ( .A(G116), .B(n628), .ZN(G18) );
  XOR2_X1 U700 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n631) );
  XNOR2_X1 U701 ( .A(G125), .B(n629), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n631), .B(n630), .ZN(G27) );
  XOR2_X1 U703 ( .A(G134), .B(n632), .Z(G36) );
  XNOR2_X1 U704 ( .A(G140), .B(n633), .ZN(G42) );
  NOR2_X1 U705 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U706 ( .A(n636), .B(KEYINPUT116), .ZN(n637) );
  NOR2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n644) );
  NOR2_X1 U710 ( .A1(n644), .A2(n662), .ZN(n658) );
  XOR2_X1 U711 ( .A(KEYINPUT50), .B(n646), .Z(n652) );
  NAND2_X1 U712 ( .A1(n486), .A2(n647), .ZN(n648) );
  XNOR2_X1 U713 ( .A(n648), .B(KEYINPUT49), .ZN(n650) );
  NOR2_X1 U714 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U715 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U716 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U717 ( .A(KEYINPUT51), .B(n655), .ZN(n656) );
  NOR2_X1 U718 ( .A1(n663), .A2(n656), .ZN(n657) );
  NOR2_X1 U719 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U720 ( .A(n659), .B(KEYINPUT52), .ZN(n660) );
  NOR2_X1 U721 ( .A1(n661), .A2(n660), .ZN(n665) );
  NOR2_X1 U722 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U723 ( .A1(n665), .A2(n664), .ZN(n668) );
  BUF_X1 U724 ( .A(n666), .Z(n667) );
  NAND2_X1 U725 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U726 ( .A1(n669), .A2(G953), .ZN(n670) );
  XNOR2_X1 U727 ( .A(n670), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U728 ( .A1(n671), .A2(G210), .ZN(n674) );
  XNOR2_X1 U729 ( .A(KEYINPUT56), .B(n676), .ZN(G51) );
  XOR2_X1 U730 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n679) );
  XNOR2_X1 U731 ( .A(n677), .B(KEYINPUT117), .ZN(n678) );
  XNOR2_X1 U732 ( .A(n679), .B(n678), .ZN(n681) );
  NAND2_X1 U733 ( .A1(n671), .A2(G469), .ZN(n680) );
  XOR2_X1 U734 ( .A(n681), .B(n680), .Z(n682) );
  NOR2_X1 U735 ( .A1(n686), .A2(n682), .ZN(G54) );
  NAND2_X1 U736 ( .A1(G217), .A2(n671), .ZN(n684) );
  XNOR2_X1 U737 ( .A(n683), .B(n684), .ZN(n685) );
  NOR2_X1 U738 ( .A1(n686), .A2(n685), .ZN(G66) );
  NAND2_X1 U739 ( .A1(G953), .A2(G224), .ZN(n687) );
  XNOR2_X1 U740 ( .A(KEYINPUT61), .B(n687), .ZN(n688) );
  NAND2_X1 U741 ( .A1(n688), .A2(G898), .ZN(n689) );
  XOR2_X1 U742 ( .A(KEYINPUT122), .B(n689), .Z(n692) );
  NOR2_X1 U743 ( .A1(G953), .A2(n690), .ZN(n691) );
  NOR2_X1 U744 ( .A1(n692), .A2(n691), .ZN(n698) );
  XOR2_X1 U745 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n696) );
  NAND2_X1 U746 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U747 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U748 ( .A(n698), .B(n697), .ZN(G69) );
  XNOR2_X1 U749 ( .A(n700), .B(n699), .ZN(n704) );
  XNOR2_X1 U750 ( .A(n701), .B(n704), .ZN(n703) );
  NAND2_X1 U751 ( .A1(n703), .A2(n702), .ZN(n708) );
  XNOR2_X1 U752 ( .A(G227), .B(n704), .ZN(n705) );
  NAND2_X1 U753 ( .A1(n705), .A2(G900), .ZN(n706) );
  NAND2_X1 U754 ( .A1(n706), .A2(G953), .ZN(n707) );
  NAND2_X1 U755 ( .A1(n708), .A2(n707), .ZN(G72) );
  XNOR2_X1 U756 ( .A(n709), .B(KEYINPUT125), .ZN(G24) );
  XNOR2_X1 U757 ( .A(G137), .B(n710), .ZN(n711) );
  XNOR2_X1 U758 ( .A(n711), .B(KEYINPUT126), .ZN(G39) );
  XNOR2_X1 U759 ( .A(G110), .B(KEYINPUT112), .ZN(n713) );
  XNOR2_X1 U760 ( .A(n713), .B(n712), .ZN(G12) );
  XNOR2_X1 U761 ( .A(G119), .B(n714), .ZN(G21) );
  XNOR2_X1 U762 ( .A(G131), .B(n715), .ZN(G33) );
endmodule

