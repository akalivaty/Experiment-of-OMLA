//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0004(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n205));
  INV_X1    g0005(.A(G116), .ZN(new_n206));
  INV_X1    g0006(.A(G270), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n208), .B(new_n214), .C1(G58), .C2(G232), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G1), .B2(G20), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT64), .B(KEYINPUT1), .Z(new_n217));
  XNOR2_X1  g0017(.A(new_n216), .B(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR3_X1   g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G1), .ZN(new_n223));
  NOR3_X1   g0023(.A1(new_n223), .A2(new_n220), .A3(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NOR3_X1   g0026(.A1(new_n218), .A2(new_n222), .A3(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  INV_X1    g0031(.A(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n207), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G107), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT74), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(KEYINPUT14), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G97), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  OR2_X1    g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n229), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI211_X1 g0055(.A(G226), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n258), .A2(new_n259), .A3(G226), .A4(new_n253), .ZN(new_n260));
  AOI221_X4 g0060(.A(new_n249), .B1(G1698), .B2(new_n252), .C1(new_n257), .C2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT69), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT65), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n221), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT65), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G33), .A3(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n223), .B1(G41), .B2(G45), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G238), .ZN(new_n274));
  OAI211_X1 g0074(.A(G232), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(new_n257), .B2(new_n260), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n248), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT69), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(new_n262), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n264), .A2(new_n274), .A3(new_n280), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT13), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT71), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n284), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n263), .B1(new_n277), .B2(new_n248), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n283), .B1(new_n289), .B2(new_n279), .ZN(new_n290));
  AOI211_X1 g0090(.A(KEYINPUT69), .B(new_n263), .C1(new_n277), .C2(new_n248), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT13), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n292), .A2(KEYINPUT70), .A3(new_n293), .A4(new_n274), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT70), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(new_n284), .B2(KEYINPUT13), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n287), .A2(new_n288), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n247), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n274), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n290), .A2(new_n300), .A3(new_n291), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT70), .B1(new_n301), .B2(new_n293), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n284), .A2(new_n295), .A3(KEYINPUT13), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n284), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n304));
  AOI21_X1  g0104(.A(KEYINPUT71), .B1(new_n284), .B2(KEYINPUT13), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n302), .A2(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G169), .A3(new_n246), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n278), .A2(new_n262), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n282), .B1(new_n308), .B2(KEYINPUT69), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n309), .A2(new_n293), .A3(new_n274), .A4(new_n280), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT72), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n285), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n301), .A2(KEYINPUT72), .A3(new_n293), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n314), .A2(G179), .B1(new_n245), .B2(KEYINPUT14), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n299), .A2(new_n307), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n221), .ZN(new_n318));
  NOR2_X1   g0118(.A1(G20), .A2(G33), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G50), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n220), .A2(G33), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n320), .A2(new_n321), .B1(new_n322), .B2(new_n202), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n220), .A2(G68), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n318), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT73), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n329));
  INV_X1    g0129(.A(G13), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n330), .A2(new_n220), .A3(G1), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT12), .A3(new_n210), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT12), .B1(new_n331), .B2(new_n210), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n318), .B1(new_n223), .B2(G20), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(G68), .B2(new_n334), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n328), .A2(new_n329), .A3(new_n332), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n316), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n258), .A2(G223), .A3(new_n253), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G87), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n258), .A2(G1698), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n338), .B(new_n339), .C1(new_n340), .C2(new_n232), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n282), .B1(new_n341), .B2(new_n262), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n273), .A2(G232), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT78), .B1(new_n344), .B2(G179), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n298), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT78), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n342), .A2(new_n347), .A3(new_n348), .A4(new_n343), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n345), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT8), .B(G58), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n331), .ZN(new_n353));
  INV_X1    g0153(.A(new_n334), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(new_n352), .ZN(new_n355));
  INV_X1    g0155(.A(new_n318), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G58), .A2(G68), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n357), .B(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G58), .B2(G68), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(G20), .B1(G159), .B2(new_n319), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n254), .A2(new_n255), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT7), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(new_n220), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n258), .A2(G20), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n364), .B(G68), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n356), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n258), .A2(new_n366), .A3(G20), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT76), .B1(new_n365), .B2(KEYINPUT7), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n373), .B(G68), .C1(new_n374), .C2(new_n371), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(KEYINPUT16), .A3(new_n361), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n355), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n350), .A2(new_n377), .ZN(new_n378));
  OR3_X1    g0178(.A1(new_n378), .A2(KEYINPUT79), .A3(KEYINPUT18), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT18), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n350), .B2(new_n377), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n350), .A2(new_n377), .A3(new_n380), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(KEYINPUT79), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n344), .A2(G200), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n342), .A2(G190), .A3(new_n343), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n377), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT17), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n386), .A2(KEYINPUT17), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n379), .A2(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n258), .A2(new_n253), .ZN(new_n391));
  INV_X1    g0191(.A(G222), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n390), .B1(new_n202), .B2(new_n258), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n262), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n273), .A2(G226), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n283), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n319), .A2(G150), .ZN(new_n397));
  OAI221_X1 g0197(.A(new_n397), .B1(new_n201), .B2(new_n220), .C1(new_n351), .C2(new_n322), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n318), .B1(new_n321), .B2(new_n331), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n321), .B2(new_n354), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT9), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n396), .A2(G200), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G190), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n402), .B1(new_n401), .B2(new_n400), .C1(new_n403), .C2(new_n396), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT10), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n396), .A2(new_n298), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n400), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT66), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(G179), .B2(new_n396), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n352), .A2(new_n319), .B1(G20), .B2(G77), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT15), .B(G87), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n410), .B1(new_n322), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(new_n318), .B1(new_n202), .B2(new_n331), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n334), .A2(G77), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n258), .A2(G232), .A3(new_n253), .ZN(new_n416));
  INV_X1    g0216(.A(G107), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n416), .B1(new_n417), .B2(new_n258), .C1(new_n340), .C2(new_n211), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n262), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n273), .A2(G244), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n283), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n415), .B1(G200), .B2(new_n421), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n421), .A2(new_n403), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AND4_X1   g0225(.A1(new_n389), .A2(new_n405), .A3(new_n409), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n421), .A2(new_n298), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n415), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT67), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT67), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(new_n430), .A3(new_n415), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n421), .A2(G179), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n336), .ZN(new_n434));
  INV_X1    g0234(.A(G200), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n434), .B1(new_n297), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n403), .B1(new_n312), .B2(new_n313), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AND4_X1   g0239(.A1(new_n337), .A2(new_n426), .A3(new_n433), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n331), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(G116), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n220), .C1(G33), .C2(new_n212), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT84), .ZN(new_n445));
  AOI221_X4 g0245(.A(new_n445), .B1(new_n206), .B2(G20), .C1(new_n317), .C2(new_n221), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n206), .A2(G20), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT84), .B1(new_n318), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n444), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT20), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(KEYINPUT20), .B(new_n444), .C1(new_n446), .C2(new_n448), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n442), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n441), .B(new_n356), .C1(G1), .C2(new_n265), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G116), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n298), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n362), .A2(G303), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n459), .C1(new_n391), .C2(new_n213), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n262), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT5), .B(G41), .ZN(new_n462));
  INV_X1    g0262(.A(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G1), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(G274), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n464), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n466), .A2(new_n271), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G270), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n461), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT21), .B1(new_n457), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n442), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n318), .A2(new_n447), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n445), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n318), .A2(KEYINPUT84), .A3(new_n447), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT20), .B1(new_n475), .B2(new_n444), .ZN(new_n476));
  INV_X1    g0276(.A(new_n452), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n471), .B(new_n456), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n478), .A2(KEYINPUT21), .A3(new_n469), .A4(G169), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n411), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n441), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT19), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n220), .B1(new_n248), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  INV_X1    g0286(.A(G87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n258), .A2(new_n220), .A3(G68), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT82), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n485), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n484), .B1(new_n322), .B2(new_n212), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n490), .A2(new_n491), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n483), .B1(new_n495), .B2(new_n318), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n455), .A2(G87), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(G244), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n499));
  OAI211_X1 g0299(.A(G238), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G116), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n262), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n464), .A2(G274), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n271), .B(G250), .C1(G1), .C2(new_n463), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(new_n403), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n502), .A2(new_n262), .B1(G274), .B2(new_n464), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n435), .B1(new_n508), .B2(new_n505), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n498), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT83), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n455), .A2(new_n482), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n496), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n496), .B2(new_n512), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n506), .A2(G169), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n348), .B2(new_n506), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n469), .A2(new_n348), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n478), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n220), .B(G87), .C1(new_n254), .C2(new_n255), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT22), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT22), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n258), .A2(new_n523), .A3(new_n220), .A4(G87), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n220), .A2(G33), .A3(G116), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT85), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n522), .A2(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n220), .A2(G107), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT23), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n529), .B2(new_n532), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n318), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n454), .A2(new_n417), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n331), .A2(new_n417), .ZN(new_n538));
  XOR2_X1   g0338(.A(new_n538), .B(KEYINPUT25), .Z(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n258), .A2(G257), .A3(G1698), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n258), .A2(G250), .A3(new_n253), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n262), .A2(new_n544), .B1(new_n467), .B2(G264), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n465), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n298), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n348), .A3(new_n465), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n540), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n481), .A2(new_n518), .A3(new_n520), .A4(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(G244), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n443), .A4(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n556), .A2(KEYINPUT80), .A3(new_n262), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT80), .B1(new_n556), .B2(new_n262), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n465), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n467), .B2(G257), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n559), .A2(KEYINPUT81), .A3(new_n348), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n553), .A2(new_n554), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n555), .A2(new_n443), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n262), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT80), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n556), .A2(KEYINPUT80), .A3(new_n262), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n567), .A2(new_n348), .A3(new_n561), .A4(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT81), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n441), .A2(G97), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n364), .B(G107), .C1(new_n365), .C2(new_n366), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT6), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n212), .A2(new_n417), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(new_n486), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n417), .A2(KEYINPUT6), .A3(G97), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G20), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n319), .A2(G77), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n573), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n572), .B1(new_n581), .B2(new_n318), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n454), .A2(new_n212), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n565), .A2(new_n561), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n582), .A2(new_n584), .B1(new_n585), .B2(new_n298), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n562), .A2(new_n571), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n522), .A2(new_n524), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n528), .A2(new_n527), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n532), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT24), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n536), .B1(new_n593), .B2(new_n318), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n546), .A2(G200), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n545), .A2(G190), .A3(new_n465), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n539), .ZN(new_n597));
  AOI211_X1 g0397(.A(new_n572), .B(new_n583), .C1(new_n581), .C2(new_n318), .ZN(new_n598));
  INV_X1    g0398(.A(new_n585), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G190), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n567), .A2(new_n561), .A3(new_n568), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n598), .B(new_n600), .C1(new_n601), .C2(new_n435), .ZN(new_n602));
  INV_X1    g0402(.A(new_n478), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n469), .A2(G200), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n603), .B(new_n604), .C1(new_n403), .C2(new_n469), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n587), .A2(new_n597), .A3(new_n602), .A4(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n550), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n440), .A2(new_n607), .ZN(G372));
  NAND2_X1  g0408(.A1(new_n337), .A2(new_n433), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n388), .A2(new_n387), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n609), .A2(new_n439), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n382), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n381), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n405), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n615), .A2(new_n409), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n587), .A2(new_n602), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT86), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n498), .A2(new_n509), .ZN(new_n619));
  INV_X1    g0419(.A(new_n507), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n496), .A2(new_n512), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n619), .A2(new_n620), .B1(new_n517), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n617), .A2(new_n618), .A3(new_n597), .A4(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n540), .A2(new_n547), .A3(new_n548), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n478), .A2(G169), .A3(new_n469), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT21), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n520), .A3(new_n479), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n587), .A2(new_n597), .A3(new_n602), .A4(new_n622), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT86), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n623), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n510), .ZN(new_n634));
  INV_X1    g0434(.A(new_n514), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n496), .A2(new_n511), .A3(new_n512), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n517), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT26), .B1(new_n638), .B2(new_n587), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n562), .A2(new_n571), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n586), .A4(new_n622), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n517), .A2(new_n621), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n633), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n440), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n616), .A2(new_n647), .ZN(G369));
  NOR2_X1   g0448(.A1(new_n330), .A2(G20), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n223), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n603), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n628), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(G330), .A3(new_n605), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n540), .A2(new_n655), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n597), .A2(new_n661), .ZN(new_n662));
  MUX2_X1   g0462(.A(new_n655), .B(new_n662), .S(new_n549), .Z(new_n663));
  NAND2_X1  g0463(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n662), .A2(new_n628), .A3(new_n549), .A4(new_n656), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n624), .A2(new_n656), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT87), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(KEYINPUT87), .A3(new_n666), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n664), .A2(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n224), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n488), .A2(G116), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n219), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  INV_X1    g0479(.A(new_n622), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT26), .B1(new_n680), .B2(new_n587), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n518), .A2(new_n640), .A3(new_n641), .A4(new_n586), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n681), .B(new_n682), .C1(new_n629), .C2(new_n631), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n643), .B(KEYINPUT91), .Z(new_n684));
  OAI21_X1  g0484(.A(new_n656), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT29), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n646), .A2(new_n656), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(KEYINPUT29), .ZN(new_n688));
  AND4_X1   g0488(.A1(new_n587), .A2(new_n597), .A3(new_n602), .A4(new_n605), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n629), .A3(new_n518), .A4(new_n656), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n550), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(KEYINPUT90), .A3(new_n689), .A4(new_n656), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT88), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n544), .A2(new_n262), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n467), .A2(G264), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n695), .B1(new_n698), .B2(new_n506), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n545), .A2(KEYINPUT88), .A3(new_n505), .A4(new_n508), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n519), .A2(new_n699), .A3(new_n700), .A4(new_n599), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT89), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(new_n701), .B2(new_n702), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n546), .A2(new_n469), .A3(new_n348), .A4(new_n506), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n601), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT31), .B1(new_n708), .B2(new_n656), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  INV_X1    g0510(.A(new_n705), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n710), .B(new_n655), .C1(new_n713), .C2(new_n707), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n692), .A2(new_n694), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n688), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n679), .B1(new_n718), .B2(G1), .ZN(G364));
  AOI21_X1  g0519(.A(new_n221), .B1(G20), .B2(new_n298), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n220), .A2(new_n348), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G190), .A2(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT94), .ZN(new_n725));
  INV_X1    g0525(.A(new_n722), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n726), .A2(new_n403), .A3(G200), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n725), .A2(G77), .B1(G58), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n403), .A2(new_n435), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n722), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n728), .B1(new_n321), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT95), .Z(new_n732));
  NOR2_X1   g0532(.A1(new_n220), .A2(G179), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n435), .A2(G190), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n722), .A2(new_n735), .ZN(new_n736));
  OAI221_X1 g0536(.A(new_n258), .B1(new_n734), .B2(new_n487), .C1(new_n210), .C2(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n403), .A2(G179), .A3(G200), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n220), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n737), .B1(G97), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n733), .A2(new_n735), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G107), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n733), .A2(new_n723), .ZN(new_n745));
  INV_X1    g0545(.A(G159), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n732), .A2(new_n741), .A3(new_n744), .A4(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n736), .ZN(new_n751));
  INV_X1    g0551(.A(G317), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(KEYINPUT33), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n752), .A2(KEYINPUT33), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n751), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n745), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G329), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n755), .B(new_n757), .C1(new_n758), .C2(new_n742), .ZN(new_n759));
  INV_X1    g0559(.A(new_n734), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(G303), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n362), .B1(new_n724), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G294), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n739), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(KEYINPUT97), .B(G326), .Z(new_n766));
  INV_X1    g0566(.A(new_n730), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n763), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  INV_X1    g0569(.A(new_n727), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n761), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n721), .B1(new_n750), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n658), .A2(new_n605), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n772), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n223), .B1(new_n649), .B2(G45), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n674), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n362), .A2(new_n224), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT92), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n240), .B2(G45), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G45), .B2(new_n219), .ZN(new_n786));
  INV_X1    g0586(.A(G355), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n258), .A2(new_n224), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n786), .B1(G116), .B2(new_n224), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n776), .A2(new_n720), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n781), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n777), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n773), .A2(new_n716), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(new_n659), .A3(new_n781), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(new_n795), .ZN(G396));
  INV_X1    g0596(.A(new_n415), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n433), .B1(new_n797), .B2(new_n656), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n656), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n429), .A2(new_n431), .A3(new_n432), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n424), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n646), .A2(new_n656), .A3(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT100), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n655), .B1(new_n633), .B2(new_n645), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n805), .A2(KEYINPUT100), .A3(new_n801), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n805), .B2(new_n801), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n709), .A2(new_n714), .ZN(new_n809));
  AOI21_X1  g0609(.A(KEYINPUT90), .B1(new_n607), .B2(new_n656), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n550), .A2(new_n606), .A3(new_n691), .A4(new_n655), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G330), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n808), .A2(new_n813), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n814), .A2(new_n781), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  INV_X1    g0617(.A(G150), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n730), .A2(new_n817), .B1(new_n736), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT99), .Z(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  INV_X1    g0621(.A(new_n725), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n770), .C1(new_n746), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n258), .B1(new_n745), .B2(new_n825), .C1(new_n321), .C2(new_n734), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G58), .B2(new_n740), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n824), .B(new_n827), .C1(new_n210), .C2(new_n742), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n727), .A2(G294), .B1(G283), .B2(new_n751), .ZN(new_n829));
  INV_X1    g0629(.A(G303), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n212), .B2(new_n739), .C1(new_n830), .C2(new_n730), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n258), .B(new_n831), .C1(G107), .C2(new_n760), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n742), .A2(new_n487), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G311), .B2(new_n756), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT98), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n832), .B(new_n835), .C1(new_n206), .C2(new_n822), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n721), .B1(new_n828), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n720), .A2(new_n774), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n202), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n839), .B(new_n780), .C1(new_n775), .C2(new_n801), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n816), .A2(new_n840), .ZN(G384));
  NAND2_X1  g0641(.A1(new_n336), .A2(new_n655), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n337), .A2(new_n439), .A3(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n336), .B(new_n655), .C1(new_n316), .C2(new_n438), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n378), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n377), .A2(new_n653), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n846), .A2(new_n847), .A3(new_n386), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n375), .A2(new_n361), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT103), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n850), .A2(new_n851), .A3(new_n369), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n375), .B(new_n361), .C1(KEYINPUT103), .C2(KEYINPUT16), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n852), .A2(new_n318), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n355), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n350), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n386), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n653), .B1(new_n854), .B2(new_n855), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n849), .B1(new_n859), .B2(new_n847), .ZN(new_n860));
  INV_X1    g0660(.A(new_n858), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n389), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n860), .B(KEYINPUT38), .C1(new_n389), .C2(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n801), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n715), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n845), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT40), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n848), .B1(new_n610), .B2(new_n613), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n377), .B1(new_n350), .B2(new_n653), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT37), .B1(new_n857), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n849), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n863), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n870), .B1(new_n865), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n845), .A2(new_n868), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n871), .A2(G330), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n440), .A2(new_n717), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT104), .Z(new_n882));
  AND2_X1   g0682(.A1(new_n845), .A2(new_n868), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n883), .A2(new_n877), .B1(new_n869), .B2(new_n870), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n440), .A3(new_n812), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n440), .A2(new_n688), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n616), .A2(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n433), .A2(new_n655), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n889), .B(new_n890), .ZN(new_n891));
  AND4_X1   g0691(.A1(KEYINPUT100), .A2(new_n646), .A3(new_n656), .A4(new_n801), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT100), .B1(new_n805), .B2(new_n801), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n866), .A3(new_n845), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n614), .A2(new_n653), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n316), .A2(new_n336), .A3(new_n656), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n865), .A2(new_n876), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(KEYINPUT39), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n864), .B2(new_n865), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n898), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n895), .A2(new_n896), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n888), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n886), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n223), .B2(new_n649), .ZN(new_n908));
  OAI211_X1 g0708(.A(G20), .B(new_n268), .C1(new_n578), .C2(KEYINPUT35), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n206), .B(new_n909), .C1(KEYINPUT35), .C2(new_n578), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT36), .Z(new_n911));
  INV_X1    g0711(.A(new_n219), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n359), .A2(G77), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT101), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n210), .A2(G50), .ZN(new_n915));
  OAI211_X1 g0715(.A(G1), .B(new_n330), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(new_n911), .A3(new_n916), .ZN(G367));
  AOI22_X1  g0717(.A1(new_n727), .A2(G303), .B1(G317), .B2(new_n756), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n764), .B2(new_n736), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(G283), .B2(new_n725), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n734), .A2(new_n206), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT46), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n742), .A2(new_n212), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n739), .A2(new_n417), .ZN(new_n924));
  NOR4_X1   g0724(.A1(new_n922), .A2(new_n258), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n920), .B(new_n925), .C1(new_n762), .C2(new_n730), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n258), .B1(new_n745), .B2(new_n817), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n739), .A2(new_n210), .B1(new_n736), .B2(new_n746), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n927), .B(new_n928), .C1(G77), .C2(new_n743), .ZN(new_n929));
  INV_X1    g0729(.A(G58), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n730), .A2(new_n821), .B1(new_n734), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n725), .B2(G50), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n929), .B(new_n932), .C1(new_n818), .C2(new_n770), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT109), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT47), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n781), .B1(new_n936), .B2(new_n720), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n790), .B1(new_n224), .B2(new_n411), .C1(new_n236), .C2(new_n784), .ZN(new_n938));
  INV_X1    g0738(.A(new_n776), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n498), .A2(new_n655), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n622), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n643), .B2(new_n940), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n937), .B(new_n938), .C1(new_n939), .C2(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n587), .B(new_n602), .C1(new_n598), .C2(new_n656), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n640), .A2(new_n586), .A3(new_n655), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n944), .A2(KEYINPUT105), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT105), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n669), .A2(new_n670), .A3(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT44), .Z(new_n950));
  AOI21_X1  g0750(.A(new_n948), .B1(new_n669), .B2(new_n670), .ZN(new_n951));
  XOR2_X1   g0751(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n950), .A2(new_n664), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n664), .B1(new_n950), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT107), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n813), .B(new_n686), .C1(new_n687), .C2(KEYINPUT29), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n628), .A2(new_n656), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n663), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(new_n659), .A3(new_n665), .ZN(new_n964));
  INV_X1    g0764(.A(new_n665), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n660), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n959), .B1(new_n960), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n718), .A2(KEYINPUT107), .A3(new_n967), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT108), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n971), .B1(new_n969), .B2(new_n970), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n958), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n718), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n674), .B(KEYINPUT41), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n779), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n978));
  INV_X1    g0778(.A(new_n948), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n965), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT42), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n624), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n655), .B1(new_n982), .B2(new_n587), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n978), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n979), .A2(new_n660), .A3(new_n663), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n943), .B1(new_n977), .B2(new_n988), .ZN(G387));
  NAND2_X1  g0789(.A1(new_n969), .A2(new_n970), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n990), .B(new_n674), .C1(new_n718), .C2(new_n967), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n756), .A2(new_n766), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G322), .A2(new_n767), .B1(new_n751), .B2(G311), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n752), .B2(new_n770), .C1(new_n822), .C2(new_n830), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT48), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n758), .B2(new_n739), .C1(new_n764), .C2(new_n734), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT49), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n258), .B(new_n992), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n997), .B2(new_n996), .C1(new_n206), .C2(new_n742), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n730), .A2(new_n746), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n724), .A2(new_n210), .B1(new_n745), .B2(new_n818), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G50), .C2(new_n727), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n760), .A2(G77), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n740), .A2(new_n482), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n362), .B(new_n923), .C1(new_n352), .C2(new_n751), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n721), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n233), .A2(new_n463), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT110), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n676), .B(KEYINPUT111), .Z(new_n1010));
  NOR2_X1   g0810(.A1(new_n351), .A2(G50), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(G68), .A2(G77), .ZN(new_n1014));
  AOI21_X1  g0814(.A(G45), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1010), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1008), .A2(KEYINPUT110), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1009), .A2(new_n783), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(G107), .B2(new_n224), .C1(new_n676), .C2(new_n788), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1007), .B1(new_n790), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n780), .C1(new_n663), .C2(new_n939), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n991), .B(new_n1021), .C1(new_n778), .C2(new_n968), .ZN(G393));
  AOI22_X1  g0822(.A1(new_n243), .A2(new_n783), .B1(G97), .B2(new_n673), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n781), .B1(new_n1023), .B2(new_n790), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT114), .Z(new_n1025));
  NOR2_X1   g0825(.A1(new_n979), .A2(new_n939), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n727), .A2(G311), .B1(new_n767), .B2(G317), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT52), .Z(new_n1028));
  OAI211_X1 g0828(.A(new_n744), .B(new_n362), .C1(new_n764), .C2(new_n724), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G116), .B2(new_n740), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n751), .A2(G303), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n734), .A2(new_n758), .B1(new_n745), .B2(new_n769), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT115), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n727), .A2(G159), .B1(new_n767), .B2(G150), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT51), .Z(new_n1036));
  NOR2_X1   g0836(.A1(new_n739), .A2(new_n202), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n736), .A2(new_n321), .B1(new_n745), .B2(new_n821), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(G68), .C2(new_n760), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n725), .A2(new_n352), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n1039), .A3(new_n258), .A4(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1034), .B1(new_n1041), .B2(new_n833), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1025), .B(new_n1026), .C1(new_n720), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT113), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n956), .B2(new_n957), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n957), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(KEYINPUT113), .A3(new_n955), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1043), .B1(new_n1048), .B2(new_n779), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n990), .B1(new_n956), .B2(new_n957), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n974), .A2(new_n674), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(G390));
  NOR2_X1   g0852(.A1(new_n900), .A2(new_n902), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n774), .ZN(new_n1054));
  XOR2_X1   g0854(.A(KEYINPUT54), .B(G143), .Z(new_n1055));
  AOI22_X1  g0855(.A1(new_n725), .A2(new_n1055), .B1(G159), .B2(new_n740), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n817), .B2(new_n736), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT119), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n734), .A2(new_n818), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT53), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n258), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n767), .A2(G128), .B1(new_n756), .B2(G125), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n825), .B2(new_n770), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(new_n1060), .C2(new_n1059), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1058), .B(new_n1064), .C1(new_n321), .C2(new_n742), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n362), .B1(new_n487), .B2(new_n734), .C1(new_n770), .C2(new_n206), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1037), .B(new_n1066), .C1(G68), .C2(new_n743), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n736), .A2(new_n417), .B1(new_n745), .B2(new_n764), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n725), .B2(G97), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(new_n758), .C2(new_n730), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n721), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n351), .B2(new_n838), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1054), .A2(new_n780), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n899), .A2(new_n897), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n801), .B(new_n656), .C1(new_n683), .C2(new_n684), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT116), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n1076), .A2(new_n891), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n1076), .B2(new_n891), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n845), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1075), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n898), .B1(new_n894), .B2(new_n845), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n900), .A2(new_n902), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n715), .A2(new_n716), .A3(new_n867), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n845), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n891), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n804), .B2(new_n806), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n897), .B1(new_n1091), .B2(new_n1081), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n1053), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1093), .A2(new_n1087), .A3(new_n1082), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1073), .B1(new_n1095), .B2(new_n778), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n812), .A2(G330), .A3(new_n801), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n843), .A3(new_n844), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1087), .A2(new_n1098), .B1(new_n807), .B2(new_n891), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1087), .A2(new_n1098), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT117), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT117), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1099), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n615), .A2(new_n887), .A3(new_n880), .A4(new_n409), .ZN(new_n1106));
  OAI21_X1  g0906(.A(KEYINPUT118), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1100), .A2(new_n894), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1080), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1103), .B1(new_n1087), .B2(new_n1098), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1106), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT118), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1107), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1087), .B1(new_n1093), .B2(new_n1082), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1074), .B1(new_n1102), .B2(new_n845), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1088), .B(new_n1118), .C1(new_n1092), .C2(new_n1053), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n675), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1095), .A2(new_n1107), .A3(new_n1115), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1096), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(G378));
  OAI22_X1  g0924(.A1(new_n739), .A2(new_n818), .B1(new_n724), .B2(new_n817), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n727), .A2(G128), .B1(new_n760), .B2(new_n1055), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n730), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1125), .B(new_n1128), .C1(G132), .C2(new_n751), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT59), .ZN(new_n1130));
  AOI21_X1  g0930(.A(G41), .B1(new_n756), .B2(G124), .ZN(new_n1131));
  AOI21_X1  g0931(.A(G33), .B1(new_n743), .B2(G159), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(G50), .B1(new_n251), .B2(new_n266), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n727), .A2(G107), .B1(G58), .B2(new_n743), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n758), .B2(new_n745), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G97), .B2(new_n751), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1003), .B1(new_n206), .B2(new_n730), .C1(new_n411), .C2(new_n724), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G68), .B2(new_n740), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1137), .A2(new_n266), .A3(new_n362), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT58), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1134), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT120), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1142), .A2(KEYINPUT120), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1133), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(new_n721), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n781), .B1(new_n321), .B2(new_n838), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT121), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n653), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n400), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n405), .A2(new_n409), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1152), .B1(new_n405), .B2(new_n409), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT55), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1155), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT55), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n1153), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT56), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1156), .A2(new_n1159), .A3(KEYINPUT56), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1148), .B(new_n1150), .C1(new_n1164), .C2(new_n774), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1162), .A2(KEYINPUT122), .A3(new_n1163), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n884), .B2(G330), .ZN(new_n1167));
  AND4_X1   g0967(.A1(G330), .A2(new_n871), .A3(new_n1166), .A4(new_n878), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n904), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n879), .A2(KEYINPUT122), .A3(new_n1164), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n884), .A2(G330), .A3(new_n1166), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n905), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1165), .B1(new_n1173), .B2(new_n779), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1095), .B1(new_n1115), .B2(new_n1107), .ZN(new_n1175));
  OAI211_X1 g0975(.A(KEYINPUT57), .B(new_n1173), .C1(new_n1175), .C2(new_n1106), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n674), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1105), .A2(KEYINPUT118), .A3(new_n1106), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1114), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1120), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n1113), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT57), .B1(new_n1181), .B2(new_n1173), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1174), .B1(new_n1177), .B2(new_n1182), .ZN(G375));
  NAND2_X1  g0983(.A1(new_n1081), .A2(new_n774), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n734), .A2(new_n746), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n751), .A2(new_n1055), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n770), .B2(new_n817), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G128), .C2(new_n756), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n724), .A2(new_n818), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n258), .B1(new_n742), .B2(new_n930), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(G50), .C2(new_n740), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1188), .B(new_n1191), .C1(new_n825), .C2(new_n730), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n770), .A2(new_n758), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n362), .B1(new_n742), .B2(new_n202), .C1(new_n206), .C2(new_n736), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n482), .B2(new_n740), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n730), .A2(new_n764), .B1(new_n734), .B2(new_n212), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n725), .B2(G107), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(new_n830), .C2(new_n745), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1192), .B1(new_n1193), .B2(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1199), .A2(new_n720), .B1(new_n210), .B2(new_n838), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1184), .A2(new_n780), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1112), .B2(new_n779), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1107), .A2(new_n1115), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n976), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1202), .B1(new_n1204), .B2(new_n1205), .ZN(G381));
  INV_X1    g1006(.A(G375), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1123), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G384), .ZN(new_n1210));
  INV_X1    g1010(.A(G390), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G393), .A2(G396), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(G387), .A2(G381), .A3(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1214), .ZN(G407));
  OAI211_X1 g1015(.A(G407), .B(G213), .C1(G343), .C2(new_n1208), .ZN(G409));
  NAND2_X1  g1016(.A1(G375), .A2(G378), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1204), .A2(KEYINPUT60), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT60), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1203), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n674), .A3(new_n1220), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1221), .A2(G384), .A3(new_n1202), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G384), .B1(new_n1221), .B2(new_n1202), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(G213), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(G343), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1180), .A2(new_n674), .A3(new_n1122), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1096), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n1174), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT123), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1167), .A2(new_n1168), .A3(new_n904), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n905), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1180), .B2(new_n1113), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1235), .A2(new_n976), .B1(new_n1174), .B2(KEYINPUT123), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1226), .B1(new_n1231), .B2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1217), .A2(new_n1224), .A3(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT62), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(KEYINPUT62), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT61), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1221), .A2(new_n1202), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1210), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1221), .A2(G384), .A3(new_n1202), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1226), .A2(G2897), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1245), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1226), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT123), .B1(new_n1123), .B2(new_n1174), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1174), .A2(KEYINPUT123), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1173), .B1(new_n1175), .B2(new_n1106), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1251), .B1(new_n1205), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1249), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT57), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1106), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n1234), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n674), .A3(new_n1176), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1123), .B1(new_n1258), .B2(new_n1174), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1246), .B(new_n1248), .C1(new_n1254), .C2(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G390), .B(new_n943), .C1(new_n977), .C2(new_n988), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT124), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G393), .A2(G396), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1213), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G387), .A2(new_n1211), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1262), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1212), .B1(new_n1262), .B2(KEYINPUT124), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1269), .A2(new_n1262), .A3(new_n1266), .A4(new_n1264), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1261), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1260), .B2(new_n1238), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1254), .A2(new_n1259), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT63), .B1(new_n1275), .B2(new_n1224), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1268), .A2(new_n1241), .A3(new_n1270), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(new_n1274), .A2(new_n1276), .A3(KEYINPUT125), .A4(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1248), .A2(new_n1246), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1238), .B1(new_n1275), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT63), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1277), .B1(new_n1273), .B2(new_n1238), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1279), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1272), .B1(new_n1278), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1272), .B(KEYINPUT126), .C1(new_n1278), .C2(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(new_n1208), .A2(new_n1217), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1224), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1291), .B(new_n1271), .Z(G402));
endmodule


