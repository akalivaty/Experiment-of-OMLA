

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, n1043, G284, G297, G282, G295, n520, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n718), .A2(n717), .ZN(n719) );
  BUF_X1 U554 ( .A(n1043), .Z(G164) );
  NOR2_X1 U555 ( .A1(n789), .A2(n640), .ZN(n620) );
  XNOR2_X1 U556 ( .A(n522), .B(KEYINPUT102), .ZN(n608) );
  NAND2_X1 U557 ( .A1(n631), .A2(G1996), .ZN(n604) );
  INV_X1 U558 ( .A(KEYINPUT64), .ZN(n520) );
  NOR2_X1 U559 ( .A1(n1043), .A2(G1384), .ZN(n721) );
  NOR2_X1 U560 ( .A1(n544), .A2(n543), .ZN(n1043) );
  AND2_X1 U561 ( .A1(n531), .A2(G2104), .ZN(n889) );
  NOR2_X2 U562 ( .A1(G2104), .A2(G2105), .ZN(n530) );
  XNOR2_X2 U563 ( .A(n603), .B(n520), .ZN(n631) );
  NAND2_X1 U564 ( .A1(n606), .A2(n605), .ZN(n522) );
  NOR2_X1 U565 ( .A1(n700), .A2(KEYINPUT33), .ZN(n704) );
  AND2_X1 U566 ( .A1(n526), .A2(G2105), .ZN(n894) );
  OR2_X1 U567 ( .A1(n675), .A2(n674), .ZN(n676) );
  OR2_X1 U568 ( .A1(n643), .A2(n642), .ZN(n647) );
  XNOR2_X1 U569 ( .A(n672), .B(KEYINPUT31), .ZN(n684) );
  OR2_X1 U570 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U571 ( .A(KEYINPUT23), .B(KEYINPUT67), .ZN(n524) );
  XNOR2_X1 U572 ( .A(n699), .B(n698), .ZN(n700) );
  INV_X1 U573 ( .A(KEYINPUT65), .ZN(n698) );
  NOR2_X1 U574 ( .A1(n536), .A2(n535), .ZN(G160) );
  OR2_X1 U575 ( .A1(n702), .A2(n713), .ZN(n523) );
  INV_X1 U576 ( .A(KEYINPUT27), .ZN(n632) );
  NOR2_X1 U577 ( .A1(n687), .A2(n665), .ZN(n666) );
  INV_X1 U578 ( .A(n631), .ZN(n664) );
  BUF_X1 U579 ( .A(n664), .Z(n656) );
  NAND2_X1 U580 ( .A1(n523), .A2(n999), .ZN(n703) );
  INV_X1 U581 ( .A(G2105), .ZN(n531) );
  INV_X1 U582 ( .A(G2104), .ZN(n526) );
  AND2_X1 U583 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U584 ( .A1(G543), .A2(G651), .ZN(n805) );
  NOR2_X1 U585 ( .A1(G651), .A2(n577), .ZN(n809) );
  XNOR2_X1 U586 ( .A(n525), .B(n524), .ZN(n529) );
  NAND2_X1 U587 ( .A1(G101), .A2(n889), .ZN(n525) );
  NAND2_X1 U588 ( .A1(G125), .A2(n894), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(KEYINPUT66), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n536) );
  XOR2_X2 U591 ( .A(KEYINPUT17), .B(n530), .Z(n890) );
  NAND2_X1 U592 ( .A1(G137), .A2(n890), .ZN(n534) );
  NAND2_X1 U593 ( .A1(G2105), .A2(G2104), .ZN(n532) );
  XOR2_X1 U594 ( .A(KEYINPUT68), .B(n532), .Z(n726) );
  NAND2_X1 U595 ( .A1(G113), .A2(n726), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U597 ( .A1(n890), .A2(G138), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n889), .A2(G102), .ZN(n537) );
  XOR2_X1 U599 ( .A(KEYINPUT89), .B(n537), .Z(n538) );
  NAND2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U601 ( .A(n540), .B(KEYINPUT90), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n894), .A2(G126), .ZN(n542) );
  NAND2_X1 U603 ( .A1(G114), .A2(n726), .ZN(n541) );
  NAND2_X1 U604 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U605 ( .A(G543), .B(KEYINPUT0), .Z(n577) );
  NAND2_X1 U606 ( .A1(G52), .A2(n809), .ZN(n547) );
  INV_X1 U607 ( .A(G651), .ZN(n548) );
  NOR2_X1 U608 ( .A1(G543), .A2(n548), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT1), .B(n545), .Z(n810) );
  NAND2_X1 U610 ( .A1(G64), .A2(n810), .ZN(n546) );
  NAND2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G90), .A2(n805), .ZN(n550) );
  NOR2_X1 U613 ( .A1(n577), .A2(n548), .ZN(n806) );
  NAND2_X1 U614 ( .A1(G77), .A2(n806), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n551), .Z(n552) );
  NOR2_X1 U617 ( .A1(n553), .A2(n552), .ZN(G171) );
  NAND2_X1 U618 ( .A1(G50), .A2(n809), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G62), .A2(n810), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(KEYINPUT83), .B(n556), .ZN(n560) );
  NAND2_X1 U622 ( .A1(G88), .A2(n805), .ZN(n558) );
  NAND2_X1 U623 ( .A1(G75), .A2(n806), .ZN(n557) );
  AND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(G303) );
  NAND2_X1 U626 ( .A1(n806), .A2(G76), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT72), .B(n561), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n805), .A2(G89), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT4), .B(n562), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT5), .ZN(n571) );
  XNOR2_X1 U632 ( .A(KEYINPUT73), .B(KEYINPUT6), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G51), .A2(n809), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G63), .A2(n810), .ZN(n566) );
  NAND2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT7), .B(n572), .ZN(G168) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U640 ( .A1(G49), .A2(n809), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G74), .A2(G651), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U643 ( .A1(n810), .A2(n575), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n576), .B(KEYINPUT80), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G87), .A2(n577), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U647 ( .A(KEYINPUT81), .B(n580), .Z(G288) );
  NAND2_X1 U648 ( .A1(G48), .A2(n809), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n581), .B(KEYINPUT82), .ZN(n588) );
  NAND2_X1 U650 ( .A1(G86), .A2(n805), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G61), .A2(n810), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n806), .A2(G73), .ZN(n584) );
  XOR2_X1 U654 ( .A(KEYINPUT2), .B(n584), .Z(n585) );
  NOR2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(G305) );
  NAND2_X1 U657 ( .A1(G85), .A2(n805), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G72), .A2(n806), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U660 ( .A1(G47), .A2(n809), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G60), .A2(n810), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n593) );
  OR2_X1 U663 ( .A1(n594), .A2(n593), .ZN(G290) );
  NAND2_X1 U664 ( .A1(G54), .A2(n809), .ZN(n596) );
  NAND2_X1 U665 ( .A1(G66), .A2(n810), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G92), .A2(n805), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G79), .A2(n806), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U670 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U671 ( .A(n601), .B(KEYINPUT15), .Z(n984) );
  INV_X1 U672 ( .A(n984), .ZN(n789) );
  NAND2_X1 U673 ( .A1(G160), .A2(G40), .ZN(n720) );
  INV_X1 U674 ( .A(n720), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n602), .A2(n721), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n604), .B(KEYINPUT26), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G1341), .A2(n664), .ZN(n605) );
  INV_X1 U678 ( .A(n608), .ZN(n619) );
  NAND2_X1 U679 ( .A1(G81), .A2(n805), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n609), .B(KEYINPUT12), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT70), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G68), .A2(n806), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n613), .B(KEYINPUT13), .ZN(n615) );
  NAND2_X1 U685 ( .A1(G43), .A2(n809), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U687 ( .A1(n810), .A2(G56), .ZN(n616) );
  XOR2_X1 U688 ( .A(KEYINPUT14), .B(n616), .Z(n617) );
  NOR2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n994) );
  NAND2_X1 U690 ( .A1(n619), .A2(n994), .ZN(n640) );
  XNOR2_X1 U691 ( .A(n620), .B(KEYINPUT103), .ZN(n639) );
  INV_X1 U692 ( .A(n664), .ZN(n652) );
  NAND2_X1 U693 ( .A1(n652), .A2(G2067), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT104), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n656), .A2(G1348), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n637) );
  NAND2_X1 U697 ( .A1(G53), .A2(n809), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G65), .A2(n810), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U700 ( .A1(G91), .A2(n805), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G78), .A2(n806), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U704 ( .A(n630), .B(KEYINPUT69), .Z(n777) );
  NAND2_X1 U705 ( .A1(n631), .A2(G2072), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n664), .A2(G1956), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U709 ( .A(KEYINPUT101), .B(n636), .ZN(n644) );
  NAND2_X1 U710 ( .A1(n777), .A2(n644), .ZN(n641) );
  AND2_X1 U711 ( .A1(n637), .A2(n641), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n649) );
  NAND2_X1 U713 ( .A1(n640), .A2(n789), .ZN(n643) );
  INV_X1 U714 ( .A(n641), .ZN(n642) );
  NOR2_X1 U715 ( .A1(n644), .A2(n777), .ZN(n645) );
  XOR2_X1 U716 ( .A(n645), .B(KEYINPUT28), .Z(n646) );
  AND2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n651) );
  XNOR2_X1 U719 ( .A(KEYINPUT105), .B(KEYINPUT29), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(n682) );
  XNOR2_X1 U721 ( .A(G2078), .B(KEYINPUT25), .ZN(n1021) );
  NAND2_X1 U722 ( .A1(n652), .A2(n1021), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n653), .B(KEYINPUT100), .ZN(n655) );
  INV_X1 U724 ( .A(G1961), .ZN(n867) );
  NAND2_X1 U725 ( .A1(n656), .A2(n867), .ZN(n654) );
  NAND2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n669) );
  NAND2_X1 U727 ( .A1(n669), .A2(G171), .ZN(n683) );
  NOR2_X1 U728 ( .A1(n656), .A2(G2090), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n656), .A2(G8), .ZN(n713) );
  NOR2_X1 U730 ( .A1(G1971), .A2(n713), .ZN(n657) );
  NOR2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n659), .A2(G303), .ZN(n673) );
  INV_X1 U733 ( .A(n673), .ZN(n660) );
  OR2_X1 U734 ( .A1(n660), .A2(G286), .ZN(n662) );
  AND2_X1 U735 ( .A1(n683), .A2(n662), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n682), .A2(n661), .ZN(n677) );
  INV_X1 U737 ( .A(n662), .ZN(n675) );
  INV_X1 U738 ( .A(G8), .ZN(n665) );
  NOR2_X1 U739 ( .A1(n665), .A2(G1966), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n664), .A2(n663), .ZN(n686) );
  NOR2_X1 U741 ( .A1(n664), .A2(G2084), .ZN(n687) );
  NAND2_X1 U742 ( .A1(n686), .A2(n666), .ZN(n667) );
  XNOR2_X1 U743 ( .A(KEYINPUT30), .B(n667), .ZN(n668) );
  NOR2_X1 U744 ( .A1(G168), .A2(n668), .ZN(n671) );
  NOR2_X1 U745 ( .A1(G171), .A2(n669), .ZN(n670) );
  AND2_X1 U746 ( .A1(n684), .A2(n673), .ZN(n674) );
  NAND2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U748 ( .A1(n678), .A2(G8), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n679), .B(KEYINPUT32), .ZN(n706) );
  NAND2_X1 U750 ( .A1(G1976), .A2(G288), .ZN(n992) );
  INV_X1 U751 ( .A(n713), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n992), .A2(n680), .ZN(n695) );
  INV_X1 U753 ( .A(n695), .ZN(n681) );
  AND2_X1 U754 ( .A1(n706), .A2(n681), .ZN(n693) );
  NAND2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n691) );
  INV_X1 U757 ( .A(n686), .ZN(n689) );
  AND2_X1 U758 ( .A1(G8), .A2(n687), .ZN(n688) );
  NOR2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U761 ( .A(KEYINPUT106), .B(n692), .ZN(n705) );
  NAND2_X1 U762 ( .A1(n693), .A2(n705), .ZN(n697) );
  NOR2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n701) );
  NOR2_X1 U764 ( .A1(G1971), .A2(G303), .ZN(n694) );
  NOR2_X1 U765 ( .A1(n701), .A2(n694), .ZN(n1006) );
  OR2_X1 U766 ( .A1(n695), .A2(n1006), .ZN(n696) );
  NAND2_X1 U767 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n701), .A2(KEYINPUT33), .ZN(n702) );
  XOR2_X1 U769 ( .A(G1981), .B(G305), .Z(n999) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n718) );
  NAND2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n709) );
  NOR2_X1 U772 ( .A1(G2090), .A2(G303), .ZN(n707) );
  NAND2_X1 U773 ( .A1(G8), .A2(n707), .ZN(n708) );
  NAND2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U775 ( .A1(n710), .A2(n713), .ZN(n716) );
  NOR2_X1 U776 ( .A1(G1981), .A2(G305), .ZN(n711) );
  XNOR2_X1 U777 ( .A(n711), .B(KEYINPUT24), .ZN(n712) );
  XNOR2_X1 U778 ( .A(n712), .B(KEYINPUT99), .ZN(n714) );
  OR2_X1 U779 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U781 ( .A(n719), .B(KEYINPUT107), .ZN(n758) );
  NOR2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n771) );
  NAND2_X1 U783 ( .A1(n890), .A2(G140), .ZN(n722) );
  XNOR2_X1 U784 ( .A(n722), .B(KEYINPUT92), .ZN(n724) );
  NAND2_X1 U785 ( .A1(G104), .A2(n889), .ZN(n723) );
  NAND2_X1 U786 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U787 ( .A(KEYINPUT34), .B(n725), .ZN(n731) );
  NAND2_X1 U788 ( .A1(n894), .A2(G128), .ZN(n728) );
  NAND2_X1 U789 ( .A1(G116), .A2(n726), .ZN(n727) );
  NAND2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U791 ( .A(KEYINPUT35), .B(n729), .Z(n730) );
  NOR2_X1 U792 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U793 ( .A(KEYINPUT36), .B(n732), .ZN(n904) );
  XOR2_X1 U794 ( .A(G2067), .B(KEYINPUT37), .Z(n733) );
  XNOR2_X1 U795 ( .A(KEYINPUT91), .B(n733), .ZN(n769) );
  NOR2_X1 U796 ( .A1(n904), .A2(n769), .ZN(n942) );
  NAND2_X1 U797 ( .A1(n771), .A2(n942), .ZN(n766) );
  XNOR2_X1 U798 ( .A(KEYINPUT95), .B(G1991), .ZN(n1022) );
  NAND2_X1 U799 ( .A1(G119), .A2(n894), .ZN(n740) );
  NAND2_X1 U800 ( .A1(G95), .A2(n889), .ZN(n735) );
  NAND2_X1 U801 ( .A1(G131), .A2(n890), .ZN(n734) );
  NAND2_X1 U802 ( .A1(n735), .A2(n734), .ZN(n738) );
  NAND2_X1 U803 ( .A1(G107), .A2(n726), .ZN(n736) );
  XNOR2_X1 U804 ( .A(KEYINPUT93), .B(n736), .ZN(n737) );
  NOR2_X1 U805 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U806 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U807 ( .A(n741), .B(KEYINPUT94), .Z(n909) );
  NOR2_X1 U808 ( .A1(n1022), .A2(n909), .ZN(n742) );
  XNOR2_X1 U809 ( .A(n742), .B(KEYINPUT96), .ZN(n753) );
  NAND2_X1 U810 ( .A1(n894), .A2(G129), .ZN(n744) );
  NAND2_X1 U811 ( .A1(G117), .A2(n726), .ZN(n743) );
  NAND2_X1 U812 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U813 ( .A(KEYINPUT97), .B(n745), .ZN(n751) );
  NAND2_X1 U814 ( .A1(G105), .A2(n889), .ZN(n746) );
  XOR2_X1 U815 ( .A(KEYINPUT38), .B(n746), .Z(n749) );
  NAND2_X1 U816 ( .A1(n890), .A2(G141), .ZN(n747) );
  XOR2_X1 U817 ( .A(KEYINPUT98), .B(n747), .Z(n748) );
  NOR2_X1 U818 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U819 ( .A1(n751), .A2(n750), .ZN(n903) );
  AND2_X1 U820 ( .A1(G1996), .A2(n903), .ZN(n752) );
  NOR2_X1 U821 ( .A1(n753), .A2(n752), .ZN(n950) );
  INV_X1 U822 ( .A(n950), .ZN(n754) );
  NAND2_X1 U823 ( .A1(n754), .A2(n771), .ZN(n759) );
  AND2_X1 U824 ( .A1(n766), .A2(n759), .ZN(n756) );
  XNOR2_X1 U825 ( .A(G1986), .B(G290), .ZN(n991) );
  NAND2_X1 U826 ( .A1(n991), .A2(n771), .ZN(n755) );
  NAND2_X1 U827 ( .A1(n758), .A2(n757), .ZN(n774) );
  NOR2_X1 U828 ( .A1(G1996), .A2(n903), .ZN(n940) );
  INV_X1 U829 ( .A(n759), .ZN(n762) );
  NOR2_X1 U830 ( .A1(G1986), .A2(G290), .ZN(n760) );
  AND2_X1 U831 ( .A1(n1022), .A2(n909), .ZN(n948) );
  NOR2_X1 U832 ( .A1(n760), .A2(n948), .ZN(n761) );
  NOR2_X1 U833 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U834 ( .A1(n940), .A2(n763), .ZN(n764) );
  XNOR2_X1 U835 ( .A(KEYINPUT108), .B(n764), .ZN(n765) );
  XNOR2_X1 U836 ( .A(n765), .B(KEYINPUT39), .ZN(n767) );
  NAND2_X1 U837 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U838 ( .A(KEYINPUT109), .B(n768), .Z(n770) );
  NAND2_X1 U839 ( .A1(n904), .A2(n769), .ZN(n944) );
  NAND2_X1 U840 ( .A1(n770), .A2(n944), .ZN(n772) );
  NAND2_X1 U841 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U842 ( .A1(n774), .A2(n773), .ZN(n776) );
  XNOR2_X1 U843 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n775) );
  XNOR2_X1 U844 ( .A(n776), .B(n775), .ZN(G329) );
  INV_X1 U845 ( .A(n777), .ZN(G299) );
  AND2_X1 U846 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U847 ( .A1(n726), .A2(G111), .ZN(n784) );
  NAND2_X1 U848 ( .A1(G99), .A2(n889), .ZN(n779) );
  NAND2_X1 U849 ( .A1(G135), .A2(n890), .ZN(n778) );
  NAND2_X1 U850 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U851 ( .A1(n894), .A2(G123), .ZN(n780) );
  XOR2_X1 U852 ( .A(KEYINPUT18), .B(n780), .Z(n781) );
  NOR2_X1 U853 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U854 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U855 ( .A(n785), .B(KEYINPUT78), .ZN(n945) );
  XNOR2_X1 U856 ( .A(n945), .B(G2096), .ZN(n786) );
  OR2_X1 U857 ( .A1(G2100), .A2(n786), .ZN(G156) );
  INV_X1 U858 ( .A(G120), .ZN(G236) );
  INV_X1 U859 ( .A(G69), .ZN(G235) );
  INV_X1 U860 ( .A(G108), .ZN(G238) );
  INV_X1 U861 ( .A(G171), .ZN(G301) );
  NAND2_X1 U862 ( .A1(G7), .A2(G661), .ZN(n787) );
  XOR2_X1 U863 ( .A(n787), .B(KEYINPUT10), .Z(n846) );
  NAND2_X1 U864 ( .A1(n846), .A2(G567), .ZN(n788) );
  XOR2_X1 U865 ( .A(KEYINPUT11), .B(n788), .Z(G234) );
  XOR2_X1 U866 ( .A(G860), .B(KEYINPUT71), .Z(n797) );
  NAND2_X1 U867 ( .A1(n994), .A2(n797), .ZN(G153) );
  NAND2_X1 U868 ( .A1(G868), .A2(G301), .ZN(n791) );
  INV_X1 U869 ( .A(G868), .ZN(n827) );
  NAND2_X1 U870 ( .A1(n789), .A2(n827), .ZN(n790) );
  NAND2_X1 U871 ( .A1(n791), .A2(n790), .ZN(G284) );
  XOR2_X1 U872 ( .A(KEYINPUT74), .B(G868), .Z(n792) );
  NOR2_X1 U873 ( .A1(G286), .A2(n792), .ZN(n793) );
  XOR2_X1 U874 ( .A(KEYINPUT75), .B(n793), .Z(n796) );
  NOR2_X1 U875 ( .A1(G868), .A2(G299), .ZN(n794) );
  XNOR2_X1 U876 ( .A(KEYINPUT76), .B(n794), .ZN(n795) );
  NOR2_X1 U877 ( .A1(n796), .A2(n795), .ZN(G297) );
  INV_X1 U878 ( .A(n797), .ZN(n798) );
  NAND2_X1 U879 ( .A1(n798), .A2(G559), .ZN(n799) );
  NAND2_X1 U880 ( .A1(n799), .A2(n984), .ZN(n800) );
  XNOR2_X1 U881 ( .A(n800), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U882 ( .A1(G559), .A2(n827), .ZN(n801) );
  NAND2_X1 U883 ( .A1(n984), .A2(n801), .ZN(n803) );
  NAND2_X1 U884 ( .A1(n994), .A2(n827), .ZN(n802) );
  NAND2_X1 U885 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U886 ( .A(KEYINPUT77), .B(n804), .ZN(G282) );
  NAND2_X1 U887 ( .A1(G93), .A2(n805), .ZN(n808) );
  NAND2_X1 U888 ( .A1(G80), .A2(n806), .ZN(n807) );
  NAND2_X1 U889 ( .A1(n808), .A2(n807), .ZN(n814) );
  NAND2_X1 U890 ( .A1(G55), .A2(n809), .ZN(n812) );
  NAND2_X1 U891 ( .A1(G67), .A2(n810), .ZN(n811) );
  NAND2_X1 U892 ( .A1(n812), .A2(n811), .ZN(n813) );
  OR2_X1 U893 ( .A1(n814), .A2(n813), .ZN(n826) );
  NAND2_X1 U894 ( .A1(G559), .A2(n984), .ZN(n815) );
  XOR2_X1 U895 ( .A(n994), .B(n815), .Z(n823) );
  NOR2_X1 U896 ( .A1(G860), .A2(n823), .ZN(n816) );
  XOR2_X1 U897 ( .A(KEYINPUT79), .B(n816), .Z(n817) );
  XOR2_X1 U898 ( .A(n826), .B(n817), .Z(G145) );
  XOR2_X1 U899 ( .A(n826), .B(G305), .Z(n818) );
  XNOR2_X1 U900 ( .A(n818), .B(G288), .ZN(n819) );
  XNOR2_X1 U901 ( .A(KEYINPUT19), .B(n819), .ZN(n821) );
  XOR2_X1 U902 ( .A(G290), .B(G299), .Z(n820) );
  XNOR2_X1 U903 ( .A(n821), .B(n820), .ZN(n822) );
  XOR2_X1 U904 ( .A(G303), .B(n822), .Z(n916) );
  XNOR2_X1 U905 ( .A(n916), .B(n823), .ZN(n824) );
  NAND2_X1 U906 ( .A1(n824), .A2(G868), .ZN(n825) );
  XNOR2_X1 U907 ( .A(n825), .B(KEYINPUT84), .ZN(n829) );
  NAND2_X1 U908 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U909 ( .A1(n829), .A2(n828), .ZN(G295) );
  NAND2_X1 U910 ( .A1(G2078), .A2(G2084), .ZN(n830) );
  XOR2_X1 U911 ( .A(KEYINPUT20), .B(n830), .Z(n831) );
  NAND2_X1 U912 ( .A1(G2090), .A2(n831), .ZN(n832) );
  XNOR2_X1 U913 ( .A(KEYINPUT21), .B(n832), .ZN(n833) );
  NAND2_X1 U914 ( .A1(n833), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U915 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U916 ( .A1(G235), .A2(G236), .ZN(n834) );
  XNOR2_X1 U917 ( .A(n834), .B(KEYINPUT87), .ZN(n835) );
  NOR2_X1 U918 ( .A1(G238), .A2(n835), .ZN(n836) );
  NAND2_X1 U919 ( .A1(G57), .A2(n836), .ZN(n851) );
  NAND2_X1 U920 ( .A1(n851), .A2(G567), .ZN(n843) );
  XOR2_X1 U921 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n838) );
  NAND2_X1 U922 ( .A1(G132), .A2(G82), .ZN(n837) );
  XNOR2_X1 U923 ( .A(n838), .B(n837), .ZN(n839) );
  NOR2_X1 U924 ( .A1(G218), .A2(n839), .ZN(n840) );
  NAND2_X1 U925 ( .A1(G96), .A2(n840), .ZN(n841) );
  XNOR2_X1 U926 ( .A(KEYINPUT86), .B(n841), .ZN(n852) );
  NAND2_X1 U927 ( .A1(n852), .A2(G2106), .ZN(n842) );
  NAND2_X1 U928 ( .A1(n843), .A2(n842), .ZN(n853) );
  NAND2_X1 U929 ( .A1(G661), .A2(G483), .ZN(n844) );
  XNOR2_X1 U930 ( .A(KEYINPUT88), .B(n844), .ZN(n845) );
  NOR2_X1 U931 ( .A1(n853), .A2(n845), .ZN(n850) );
  NAND2_X1 U932 ( .A1(n850), .A2(G36), .ZN(G176) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n846), .ZN(G217) );
  INV_X1 U934 ( .A(n846), .ZN(G223) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U936 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n848) );
  XOR2_X1 U938 ( .A(KEYINPUT111), .B(n848), .Z(n849) );
  NAND2_X1 U939 ( .A1(n850), .A2(n849), .ZN(G188) );
  INV_X1 U941 ( .A(G132), .ZN(G219) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G82), .ZN(G220) );
  NOR2_X1 U944 ( .A1(n852), .A2(n851), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  INV_X1 U946 ( .A(n853), .ZN(G319) );
  XOR2_X1 U947 ( .A(G2100), .B(G2096), .Z(n855) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U950 ( .A(KEYINPUT43), .B(G2090), .Z(n857) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U952 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U953 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2084), .ZN(n860) );
  XNOR2_X1 U955 ( .A(n861), .B(n860), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1976), .B(G1971), .Z(n863) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1966), .ZN(n862) );
  XNOR2_X1 U958 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U959 ( .A(n864), .B(G2474), .Z(n866) );
  XNOR2_X1 U960 ( .A(G1956), .B(G1981), .ZN(n865) );
  XNOR2_X1 U961 ( .A(n866), .B(n865), .ZN(n871) );
  XNOR2_X1 U962 ( .A(KEYINPUT41), .B(n867), .ZN(n869) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n868) );
  XNOR2_X1 U964 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U965 ( .A(n871), .B(n870), .ZN(G229) );
  XOR2_X1 U966 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n873) );
  NAND2_X1 U967 ( .A1(G124), .A2(n894), .ZN(n872) );
  XNOR2_X1 U968 ( .A(n873), .B(n872), .ZN(n880) );
  NAND2_X1 U969 ( .A1(G100), .A2(n889), .ZN(n875) );
  NAND2_X1 U970 ( .A1(G112), .A2(n726), .ZN(n874) );
  NAND2_X1 U971 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U972 ( .A(n876), .B(KEYINPUT113), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G136), .A2(n890), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U975 ( .A1(n880), .A2(n879), .ZN(G162) );
  NAND2_X1 U976 ( .A1(n894), .A2(G130), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G118), .A2(n726), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n882), .A2(n881), .ZN(n887) );
  NAND2_X1 U979 ( .A1(G106), .A2(n889), .ZN(n884) );
  NAND2_X1 U980 ( .A1(G142), .A2(n890), .ZN(n883) );
  NAND2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n885), .Z(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U984 ( .A(G162), .B(n888), .ZN(n908) );
  NAND2_X1 U985 ( .A1(G103), .A2(n889), .ZN(n892) );
  NAND2_X1 U986 ( .A1(G139), .A2(n890), .ZN(n891) );
  NAND2_X1 U987 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U988 ( .A(KEYINPUT114), .B(n893), .ZN(n899) );
  NAND2_X1 U989 ( .A1(n894), .A2(G127), .ZN(n896) );
  NAND2_X1 U990 ( .A1(G115), .A2(n726), .ZN(n895) );
  NAND2_X1 U991 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U993 ( .A1(n899), .A2(n898), .ZN(n934) );
  XOR2_X1 U994 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n901) );
  XNOR2_X1 U995 ( .A(G160), .B(n945), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n934), .B(n902), .ZN(n906) );
  XOR2_X1 U998 ( .A(n904), .B(n903), .Z(n905) );
  XNOR2_X1 U999 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n908), .B(n907), .ZN(n911) );
  XNOR2_X1 U1001 ( .A(n909), .B(G164), .ZN(n910) );
  XNOR2_X1 U1002 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n912), .ZN(G395) );
  XOR2_X1 U1004 ( .A(G301), .B(G286), .Z(n914) );
  XOR2_X1 U1005 ( .A(n984), .B(n994), .Z(n913) );
  XNOR2_X1 U1006 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1007 ( .A(n916), .B(n915), .Z(n917) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n917), .ZN(n918) );
  XOR2_X1 U1009 ( .A(KEYINPUT115), .B(n918), .Z(G397) );
  XOR2_X1 U1010 ( .A(G2451), .B(G2430), .Z(n920) );
  XNOR2_X1 U1011 ( .A(G2438), .B(G2443), .ZN(n919) );
  XNOR2_X1 U1012 ( .A(n920), .B(n919), .ZN(n926) );
  XOR2_X1 U1013 ( .A(G2435), .B(G2454), .Z(n922) );
  XNOR2_X1 U1014 ( .A(G1348), .B(G1341), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(n922), .B(n921), .ZN(n924) );
  XOR2_X1 U1016 ( .A(G2446), .B(G2427), .Z(n923) );
  XNOR2_X1 U1017 ( .A(n924), .B(n923), .ZN(n925) );
  XOR2_X1 U1018 ( .A(n926), .B(n925), .Z(n927) );
  NAND2_X1 U1019 ( .A1(G14), .A2(n927), .ZN(n933) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n933), .ZN(n930) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n928), .ZN(n929) );
  NOR2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n932) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n931) );
  NAND2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G303), .ZN(G166) );
  INV_X1 U1028 ( .A(G57), .ZN(G237) );
  INV_X1 U1029 ( .A(n933), .ZN(G401) );
  XNOR2_X1 U1030 ( .A(G164), .B(G2078), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(G2072), .B(n934), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(KEYINPUT116), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(n938), .B(KEYINPUT50), .ZN(n956) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n941), .Z(n954) );
  INV_X1 U1038 ( .A(n942), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n952) );
  XNOR2_X1 U1040 ( .A(G160), .B(G2084), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n957), .ZN(n958) );
  INV_X1 U1048 ( .A(KEYINPUT55), .ZN(n1035) );
  NAND2_X1 U1049 ( .A1(n958), .A2(n1035), .ZN(n959) );
  NAND2_X1 U1050 ( .A1(n959), .A2(G29), .ZN(n1014) );
  XOR2_X1 U1051 ( .A(G5), .B(G1961), .Z(n979) );
  XOR2_X1 U1052 ( .A(G1981), .B(G6), .Z(n961) );
  XOR2_X1 U1053 ( .A(G1341), .B(G19), .Z(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G20), .B(G1956), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT124), .B(n964), .ZN(n968) );
  XOR2_X1 U1058 ( .A(KEYINPUT125), .B(G4), .Z(n966) );
  XNOR2_X1 U1059 ( .A(G1348), .B(KEYINPUT59), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n966), .B(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(n969), .B(KEYINPUT60), .ZN(n977) );
  XNOR2_X1 U1063 ( .A(G1986), .B(G24), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(G23), .B(G1976), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1066 ( .A(G1971), .B(KEYINPUT126), .Z(n972) );
  XNOR2_X1 U1067 ( .A(G22), .B(n972), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(KEYINPUT58), .B(n975), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G21), .B(G1966), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1074 ( .A(KEYINPUT61), .B(n982), .Z(n983) );
  NOR2_X1 U1075 ( .A1(G16), .A2(n983), .ZN(n1011) );
  XOR2_X1 U1076 ( .A(G16), .B(KEYINPUT56), .Z(n1009) );
  XOR2_X1 U1077 ( .A(G1348), .B(n984), .Z(n987) );
  XNOR2_X1 U1078 ( .A(G1956), .B(G299), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(KEYINPUT122), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(G1971), .A2(G303), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n998) );
  XOR2_X1 U1084 ( .A(G301), .B(G1961), .Z(n993) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n996) );
  XOR2_X1 U1086 ( .A(n994), .B(G1341), .Z(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G168), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(n1001), .B(KEYINPUT57), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT121), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1007), .B(KEYINPUT123), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1098 ( .A(KEYINPUT127), .B(n1012), .Z(n1013) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1040) );
  XOR2_X1 U1100 ( .A(G29), .B(KEYINPUT119), .Z(n1037) );
  XNOR2_X1 U1101 ( .A(G2067), .B(G26), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G33), .B(G2072), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(G28), .A2(n1017), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT118), .B(G1996), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(G32), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1026) );
  XOR2_X1 U1108 ( .A(n1021), .B(G27), .Z(n1024) );
  XOR2_X1 U1109 ( .A(n1022), .B(G25), .Z(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1027), .B(KEYINPUT53), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(G2084), .B(G34), .Z(n1028) );
  XNOR2_X1 U1114 ( .A(KEYINPUT54), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1033) );
  XOR2_X1 U1116 ( .A(KEYINPUT117), .B(G2090), .Z(n1031) );
  XNOR2_X1 U1117 ( .A(G35), .B(n1031), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1119 ( .A(n1035), .B(n1034), .ZN(n1036) );
  NOR2_X1 U1120 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1121 ( .A(n1038), .B(KEYINPUT120), .ZN(n1039) );
  NOR2_X1 U1122 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NAND2_X1 U1123 ( .A1(n1041), .A2(G11), .ZN(n1042) );
  XNOR2_X1 U1124 ( .A(KEYINPUT62), .B(n1042), .ZN(G150) );
  INV_X1 U1125 ( .A(G150), .ZN(G311) );
endmodule

