//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  XOR2_X1   g016(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT68), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n452), .B(new_n453), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  AND2_X1   g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n463), .B1(new_n459), .B2(new_n460), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(KEYINPUT71), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n471), .A2(new_n476), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n467), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n473), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n482));
  INV_X1    g057(.A(G137), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n479), .A2(new_n484), .ZN(G160));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g062(.A(KEYINPUT72), .B(new_n467), .C1(new_n469), .C2(new_n470), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G112), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(G124), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n469), .C2(new_n470), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n500), .A2(new_n502), .A3(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  NOR3_X1   g080(.A1(new_n505), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n471), .A2(new_n476), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(G138), .B(new_n467), .C1(new_n469), .C2(new_n470), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G62), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT73), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n511), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(G75), .A2(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(G651), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n514), .A2(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G88), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n513), .B1(new_n520), .B2(new_n521), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n519), .A2(new_n523), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n514), .A2(new_n516), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n520), .A2(new_n521), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(G51), .A2(new_n524), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AOI22_X1  g115(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n522), .A2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n524), .A2(G52), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n544), .A2(KEYINPUT75), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(KEYINPUT75), .B1(new_n544), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g125(.A(KEYINPUT76), .B(new_n543), .C1(new_n546), .C2(new_n547), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(G171));
  AOI22_X1  g127(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n542), .ZN(new_n554));
  XNOR2_X1  g129(.A(KEYINPUT77), .B(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n524), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n532), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  AOI22_X1  g139(.A1(new_n530), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n542), .B1(new_n565), .B2(KEYINPUT79), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n566), .B1(KEYINPUT79), .B2(new_n565), .ZN(new_n567));
  INV_X1    g142(.A(new_n524), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  OAI21_X1  g145(.A(G53), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n568), .A2(new_n571), .B1(KEYINPUT78), .B2(KEYINPUT9), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n524), .A2(new_n569), .A3(new_n570), .A4(G53), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n572), .A2(new_n573), .B1(G91), .B2(new_n522), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n567), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  AOI22_X1  g151(.A1(new_n522), .A2(G87), .B1(new_n524), .B2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G288));
  AOI22_X1  g154(.A1(new_n522), .A2(G86), .B1(new_n524), .B2(G48), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n514), .B2(new_n516), .ZN(new_n582));
  AND2_X1   g157(.A1(G73), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n580), .A2(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n522), .A2(G85), .B1(new_n524), .B2(G47), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n542), .B2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(new_n522), .A2(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n514), .B2(new_n516), .ZN(new_n593));
  AND2_X1   g168(.A1(G79), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n524), .A2(G54), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(KEYINPUT80), .B1(new_n595), .B2(new_n596), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  MUX2_X1   g176(.A(new_n601), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g177(.A(new_n601), .B(G301), .S(G868), .Z(G321));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G168), .A2(new_n605), .ZN(new_n606));
  AOI211_X1 g181(.A(new_n604), .B(new_n606), .C1(new_n605), .C2(G299), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(new_n604), .B2(new_n606), .ZN(G297));
  XOR2_X1   g183(.A(G297), .B(KEYINPUT82), .Z(G280));
  INV_X1    g184(.A(new_n601), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  NOR2_X1   g187(.A1(new_n559), .A2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n610), .A2(new_n611), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n490), .A2(G135), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT84), .ZN(new_n619));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n620), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n495), .A2(G123), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT85), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n619), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2096), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n471), .A2(new_n476), .A3(new_n480), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n625), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT86), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2430), .Z(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n641), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT87), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n642), .A2(new_n648), .A3(new_n644), .A4(new_n645), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(G14), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n642), .A2(new_n645), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(new_n643), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n650), .A2(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT17), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2084), .B(G2090), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT88), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n661), .B(new_n658), .C1(new_n655), .C2(new_n657), .ZN(new_n662));
  INV_X1    g237(.A(new_n658), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n655), .A3(new_n657), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT90), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(KEYINPUT89), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(KEYINPUT89), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n675), .A2(new_n674), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(new_n672), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(new_n678), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n678), .A3(new_n676), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n688), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n691), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(new_n687), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n694), .B1(new_n696), .B2(new_n689), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n670), .B1(new_n693), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n691), .B1(new_n690), .B2(new_n692), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n696), .A2(new_n694), .A3(new_n689), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n699), .A2(new_n669), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  NAND2_X1  g278(.A1(G290), .A2(G16), .ZN(new_n704));
  INV_X1    g279(.A(G24), .ZN(new_n705));
  OR3_X1    g280(.A1(new_n705), .A2(KEYINPUT92), .A3(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(KEYINPUT92), .B1(new_n705), .B2(G16), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(G1986), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n495), .A2(G119), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT91), .ZN(new_n711));
  OR2_X1    g286(.A1(G95), .A2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n490), .A2(G131), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G29), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G25), .B2(G29), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT35), .B(G1991), .Z(new_n720));
  OAI21_X1  g295(.A(new_n709), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n719), .B2(new_n720), .ZN(new_n722));
  OR2_X1    g297(.A1(G6), .A2(G16), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(G305), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT32), .B(G1981), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n724), .A2(G22), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G166), .B2(new_n724), .ZN(new_n732));
  INV_X1    g307(.A(G1971), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n724), .A2(G23), .ZN(new_n735));
  INV_X1    g310(.A(G288), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(new_n724), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT33), .B(G1976), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n729), .A2(new_n730), .A3(new_n734), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(KEYINPUT34), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(KEYINPUT34), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n722), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT36), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n480), .A2(G105), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT26), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n745), .B(new_n747), .C1(G129), .C2(new_n495), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n490), .A2(G141), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G29), .ZN(new_n752));
  NOR2_X1   g327(.A1(G29), .A2(G32), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(KEYINPUT97), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT97), .B2(new_n752), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(G28), .ZN(new_n759));
  INV_X1    g334(.A(G29), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n758), .B2(G28), .ZN(new_n761));
  AND2_X1   g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  NOR2_X1   g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n759), .A2(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n624), .B2(G29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n755), .B2(new_n756), .ZN(new_n766));
  NOR2_X1   g341(.A1(G16), .A2(G19), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n559), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1341), .ZN(new_n769));
  NOR2_X1   g344(.A1(G27), .A2(G29), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G164), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT98), .B(G2078), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n766), .A2(new_n769), .A3(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G34), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(KEYINPUT24), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(KEYINPUT24), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n760), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G160), .B2(new_n760), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G2084), .Z(new_n780));
  NAND3_X1  g355(.A1(new_n471), .A2(new_n476), .A3(G127), .ZN(new_n781));
  INV_X1    g356(.A(G115), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n473), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G2105), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n490), .A2(G139), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G29), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n760), .A2(G33), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G2072), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  AND4_X1   g371(.A1(new_n757), .A2(new_n774), .A3(new_n780), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n760), .A2(G35), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G162), .B2(new_n760), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT29), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G2090), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n724), .A2(G4), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n610), .B2(new_n724), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1348), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G21), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G168), .B2(G16), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(G1966), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(G1966), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n801), .A2(new_n804), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n797), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G5), .A2(G16), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G171), .B2(G16), .ZN(new_n812));
  INV_X1    g387(.A(G1961), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n800), .A2(G2090), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n724), .A2(G20), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT23), .Z(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G299), .B2(G16), .ZN(new_n819));
  INV_X1    g394(.A(G1956), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n815), .B2(KEYINPUT99), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n760), .A2(G26), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT95), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT28), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n490), .A2(KEYINPUT94), .A3(G140), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n827));
  INV_X1    g402(.A(G140), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n489), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n831));
  INV_X1    g406(.A(G116), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(G2105), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G128), .B2(new_n495), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n825), .B1(new_n836), .B2(new_n760), .ZN(new_n837));
  INV_X1    g412(.A(G2067), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  AND4_X1   g414(.A1(new_n814), .A2(new_n816), .A3(new_n822), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n744), .A2(new_n810), .A3(new_n840), .ZN(G150));
  INV_X1    g416(.A(G150), .ZN(G311));
  XNOR2_X1  g417(.A(KEYINPUT101), .B(G860), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n610), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT38), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(new_n542), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n522), .A2(G93), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n524), .A2(G55), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n850), .B1(new_n849), .B2(new_n851), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n848), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n559), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n559), .B(new_n848), .C1(new_n853), .C2(new_n852), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n846), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n844), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n854), .A2(new_n844), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n497), .B(G160), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n624), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n716), .B(new_n627), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n490), .A2(G142), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  INV_X1    g446(.A(G118), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(G2105), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(G130), .B2(new_n495), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n869), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n836), .A2(G164), .ZN(new_n878));
  AOI21_X1  g453(.A(G164), .B1(new_n830), .B2(new_n834), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n751), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n507), .A2(new_n509), .ZN(new_n882));
  INV_X1    g457(.A(new_n504), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n835), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n750), .B1(new_n885), .B2(new_n879), .ZN(new_n886));
  AOI211_X1 g461(.A(new_n877), .B(new_n791), .C1(new_n881), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n791), .A2(new_n877), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n789), .A2(new_n790), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT102), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n881), .A2(new_n886), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n876), .A2(new_n887), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n875), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n869), .B(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n881), .A2(new_n886), .A3(new_n888), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(KEYINPUT102), .A3(new_n889), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n897), .B2(new_n891), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n868), .B1(new_n893), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n876), .B1(new_n887), .B2(new_n892), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n895), .A3(new_n891), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n867), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g480(.A1(new_n856), .A2(new_n857), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n614), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n601), .A2(G299), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n601), .A2(G299), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT41), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n910), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n912), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n907), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n912), .A2(new_n908), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(new_n907), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  XNOR2_X1  g493(.A(G290), .B(G288), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n919), .A2(KEYINPUT103), .ZN(new_n920));
  XNOR2_X1  g495(.A(G305), .B(G303), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n919), .B2(KEYINPUT103), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n920), .B(new_n922), .Z(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n915), .B(new_n925), .C1(new_n916), .C2(new_n907), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n918), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n924), .B1(new_n918), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n854), .A2(new_n605), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(G295));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n930), .ZN(G331));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n911), .A2(new_n914), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n550), .A2(KEYINPUT104), .A3(new_n551), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n906), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n937));
  AOI21_X1  g512(.A(G286), .B1(G171), .B2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n858), .A2(KEYINPUT104), .A3(new_n551), .A4(new_n550), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n936), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n936), .A2(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n916), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(G37), .B1(new_n948), .B2(new_n924), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n942), .A2(new_n947), .A3(new_n923), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n933), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(KEYINPUT44), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(G397));
  XNOR2_X1  g534(.A(new_n835), .B(new_n838), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(G1996), .B2(new_n750), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT105), .B(G1384), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT45), .B1(new_n884), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G40), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n479), .A2(new_n964), .A3(new_n484), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(G1996), .A3(new_n750), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(KEYINPUT106), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(KEYINPUT106), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n961), .A2(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n717), .A2(new_n720), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n717), .A2(new_n720), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(G290), .B(G1986), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n610), .A2(KEYINPUT60), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(G164), .A2(G1384), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n965), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n983));
  NAND3_X1  g558(.A1(new_n884), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n965), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1348), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n838), .A2(new_n981), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT60), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n601), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT117), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n981), .A2(new_n838), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n986), .A2(new_n987), .ZN(new_n993));
  AND4_X1   g568(.A1(KEYINPUT117), .A2(new_n992), .A3(new_n993), .A4(new_n990), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n979), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n993), .A3(new_n990), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n988), .A2(KEYINPUT117), .A3(new_n990), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n978), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT61), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n884), .B2(new_n982), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n477), .A2(new_n478), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G2105), .ZN(new_n1005));
  INV_X1    g580(.A(new_n484), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(G40), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n884), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT56), .B(G2072), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(G164), .B2(G1384), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1010), .A2(new_n965), .A3(new_n1014), .A4(new_n1011), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT115), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n983), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(G164), .B2(G1384), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n965), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OR3_X1    g596(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n965), .B2(new_n1019), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n820), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n1026));
  XNOR2_X1  g601(.A(G299), .B(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1017), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1017), .B2(new_n1025), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1002), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1017), .A2(new_n1025), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1027), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1017), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(KEYINPUT61), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT58), .B(G1341), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1010), .A2(new_n965), .A3(new_n1014), .ZN(new_n1037));
  OAI22_X1  g612(.A1(new_n981), .A2(new_n1036), .B1(new_n1037), .B2(G1996), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n559), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT59), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1001), .A2(new_n1030), .A3(new_n1035), .A4(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n988), .A2(new_n601), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT116), .B1(new_n1043), .B2(new_n1028), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1034), .B(new_n1045), .C1(new_n1029), .C2(new_n1042), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n1037), .B2(G2078), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n986), .A2(new_n813), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n884), .A2(KEYINPUT45), .A3(new_n982), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1049), .A2(G2078), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n965), .A3(new_n1014), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT121), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1052), .A2(new_n1058), .A3(new_n1055), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1051), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT122), .B1(new_n1060), .B2(G301), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1059), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1058), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1050), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1065), .A3(G171), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1051), .A2(G171), .ZN(new_n1067));
  INV_X1    g642(.A(new_n963), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(new_n965), .A3(new_n1010), .A4(new_n1054), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1052), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1061), .A2(new_n1066), .A3(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  INV_X1    g649(.A(G1981), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n580), .A2(new_n1075), .A3(new_n584), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1075), .B1(new_n580), .B2(new_n584), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G305), .A2(G1981), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(KEYINPUT49), .A3(new_n1076), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n965), .A2(new_n980), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .A4(G8), .ZN(new_n1083));
  INV_X1    g658(.A(G1976), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(G288), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n736), .A2(G1976), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1082), .A2(new_n1085), .A3(G8), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1082), .A2(G8), .A3(new_n1086), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT52), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT109), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT109), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1092), .A3(KEYINPUT52), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1088), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1037), .A2(new_n733), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(G2090), .B2(new_n986), .ZN(new_n1096));
  NAND2_X1  g671(.A1(G303), .A2(G8), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1101));
  OR3_X1    g676(.A1(new_n1100), .A2(KEYINPUT108), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT108), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1096), .A2(new_n1102), .A3(G8), .A4(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1094), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1067), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1050), .A2(new_n1052), .A3(new_n1069), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(G171), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G8), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1024), .ZN(new_n1112));
  INV_X1    g687(.A(G2090), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n1022), .A4(new_n1021), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1111), .B1(new_n1114), .B2(new_n1095), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1105), .A2(new_n1110), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1053), .A2(new_n965), .A3(new_n1014), .ZN(new_n1120));
  INV_X1    g695(.A(G1966), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT112), .B(G2084), .Z(new_n1123));
  NAND4_X1  g698(.A1(new_n984), .A2(new_n965), .A3(new_n985), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1122), .A2(KEYINPUT118), .A3(new_n1124), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(G168), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(G8), .B1(KEYINPUT119), .B2(KEYINPUT51), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(KEYINPUT119), .B2(KEYINPUT51), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1125), .A2(G8), .ZN(new_n1133));
  NOR2_X1   g708(.A1(G168), .A2(new_n1111), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(KEYINPUT51), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1132), .A2(new_n1136), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1119), .A2(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1048), .A2(new_n1073), .A3(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1094), .B(new_n1104), .C1(new_n1117), .C2(new_n1115), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1137), .A2(new_n1134), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1129), .A2(new_n1131), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1145), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT62), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1142), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1125), .A2(G8), .A3(G168), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1141), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT113), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1117), .B1(new_n1096), .B2(G8), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1125), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1094), .A2(new_n1104), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1154), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1105), .A2(KEYINPUT113), .A3(new_n1157), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1153), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1083), .A2(new_n1084), .A3(new_n736), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1076), .ZN(new_n1164));
  AOI211_X1 g739(.A(new_n1111), .B(new_n981), .C1(new_n1164), .C2(KEYINPUT110), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1164), .A2(KEYINPUT110), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1104), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1165), .A2(new_n1166), .B1(new_n1167), .B2(new_n1094), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1150), .A2(new_n1162), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n977), .B1(new_n1140), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n966), .B1(new_n960), .B2(new_n751), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n966), .A2(G1996), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT46), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT125), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1174), .B(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n972), .B(KEYINPUT123), .Z(new_n1178));
  AOI22_X1  g753(.A1(new_n1178), .A2(new_n971), .B1(new_n838), .B2(new_n836), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1177), .B1(new_n1179), .B2(new_n966), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n971), .A2(KEYINPUT126), .A3(new_n974), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT126), .B1(new_n971), .B2(new_n974), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n966), .A2(G1986), .A3(G290), .ZN(new_n1183));
  XOR2_X1   g758(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1184));
  XNOR2_X1  g759(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1181), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1180), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1170), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g763(.A1(G227), .A2(new_n465), .ZN(new_n1190));
  AOI21_X1  g764(.A(new_n1190), .B1(new_n650), .B2(new_n653), .ZN(new_n1191));
  AND2_X1   g765(.A1(new_n1191), .A2(new_n702), .ZN(new_n1192));
  OAI211_X1 g766(.A(new_n904), .B(new_n1192), .C1(new_n952), .C2(new_n953), .ZN(G225));
  INV_X1    g767(.A(G225), .ZN(G308));
endmodule


