//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1193, new_n1194, new_n1195,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n202), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT64), .B(G50), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n217), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n207), .A2(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G50), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G150), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n208), .A2(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n260), .B1(G20), .B2(new_n204), .ZN(new_n261));
  INV_X1    g0061(.A(new_n252), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n255), .B1(G50), .B2(new_n249), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT9), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  INV_X1    g0065(.A(new_n217), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G226), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n275), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT3), .B(G33), .Z(new_n281));
  AOI22_X1  g0081(.A1(new_n280), .A2(G223), .B1(G77), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G222), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g0086(.A(new_n274), .B(new_n277), .C1(new_n286), .C2(new_n275), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G190), .ZN(new_n288));
  INV_X1    g0088(.A(G200), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n264), .B(new_n288), .C1(new_n289), .C2(new_n287), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT10), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n263), .B1(new_n287), .B2(G169), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G97), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n299), .B1(new_n285), .B2(new_n276), .C1(new_n233), .C2(new_n279), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n275), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n275), .A2(new_n272), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n274), .B1(G238), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT13), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(KEYINPUT13), .A3(new_n303), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(G169), .A3(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n308), .A2(KEYINPUT14), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(KEYINPUT14), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT66), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n301), .A2(new_n303), .B1(KEYINPUT66), .B2(KEYINPUT13), .ZN(new_n313));
  OAI21_X1  g0113(.A(G179), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n309), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n250), .A2(new_n203), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT12), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n221), .B2(new_n259), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n253), .A2(G68), .A3(new_n254), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT11), .B1(new_n319), .B2(new_n252), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n315), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n306), .A2(new_n307), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n324), .B1(new_n326), .B2(G200), .ZN(new_n327));
  OAI21_X1  g0127(.A(G190), .B1(new_n312), .B2(new_n313), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT3), .ZN(new_n332));
  INV_X1    g0132(.A(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT67), .B(G33), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(new_n332), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G223), .A2(G1698), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n276), .B2(G1698), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n336), .A2(new_n338), .B1(G33), .B2(G87), .ZN(new_n339));
  INV_X1    g0139(.A(new_n275), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n302), .A2(G232), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n273), .B2(new_n269), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n341), .A2(G190), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n341), .A2(new_n343), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT69), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT69), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n341), .B2(new_n343), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n344), .B1(new_n349), .B2(new_n289), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT17), .ZN(new_n351));
  INV_X1    g0151(.A(new_n253), .ZN(new_n352));
  INV_X1    g0152(.A(new_n258), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n254), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n352), .A2(new_n354), .B1(new_n249), .B2(new_n353), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT7), .B1(new_n336), .B2(G20), .ZN(new_n357));
  NOR2_X1   g0157(.A1(KEYINPUT3), .A2(G33), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n333), .A2(KEYINPUT67), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT67), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G33), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n358), .B1(new_n362), .B2(KEYINPUT3), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(new_n208), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n357), .A2(new_n365), .A3(G68), .ZN(new_n366));
  XNOR2_X1  g0166(.A(G58), .B(G68), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(G20), .B1(G159), .B2(new_n256), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n252), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT7), .B1(new_n334), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT68), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n373), .A2(new_n374), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n362), .A2(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(KEYINPUT7), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n375), .A2(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT16), .B1(new_n380), .B2(new_n368), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n356), .B1(new_n371), .B2(new_n381), .ZN(new_n382));
  OR3_X1    g0182(.A1(new_n350), .A2(new_n351), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G169), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n349), .A2(new_n384), .B1(new_n292), .B2(new_n345), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT18), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT18), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n385), .A2(new_n388), .A3(new_n382), .ZN(new_n389));
  INV_X1    g0189(.A(new_n369), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT16), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n380), .A2(new_n368), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n370), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n393), .A3(new_n252), .ZN(new_n394));
  AOI21_X1  g0194(.A(G200), .B1(new_n346), .B2(new_n348), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n394), .B(new_n356), .C1(new_n395), .C2(new_n344), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n351), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n383), .A2(new_n387), .A3(new_n389), .A4(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n280), .A2(G238), .B1(G107), .B2(new_n281), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n233), .B2(new_n285), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n275), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n274), .B1(G244), .B2(new_n302), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT65), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(KEYINPUT65), .A3(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G190), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n353), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT15), .B(G87), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n411), .A2(new_n259), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n262), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n253), .A2(G77), .A3(new_n254), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(G77), .B2(new_n249), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n409), .B(new_n416), .C1(new_n408), .C2(new_n289), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n416), .B1(new_n408), .B2(new_n292), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n406), .A2(new_n384), .A3(new_n407), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n298), .A2(new_n331), .A3(new_n399), .A4(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT24), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n332), .B1(new_n359), .B2(new_n361), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n208), .B(G87), .C1(new_n424), .C2(new_n358), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT78), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT78), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n336), .A2(new_n427), .A3(new_n208), .A4(G87), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(KEYINPUT22), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G87), .ZN(new_n430));
  OR4_X1    g0230(.A1(KEYINPUT22), .A2(new_n281), .A3(G20), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT75), .B(G116), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n335), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n208), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT79), .B1(new_n208), .B2(G107), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT23), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n423), .B1(new_n432), .B2(new_n439), .ZN(new_n440));
  AOI211_X1 g0240(.A(KEYINPUT24), .B(new_n438), .C1(new_n429), .C2(new_n431), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n252), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n262), .B(new_n249), .C1(G1), .C2(new_n333), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n223), .B1(KEYINPUT80), .B2(KEYINPUT25), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n445), .B1(new_n446), .B2(new_n249), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n250), .A2(KEYINPUT80), .A3(KEYINPUT25), .A4(new_n223), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n444), .A2(G107), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n271), .A2(G1), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT72), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(new_n270), .A3(KEYINPUT5), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT5), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT72), .B1(new_n453), .B2(G41), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(G41), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n450), .B(new_n452), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(G264), .A3(new_n340), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT81), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n207), .A2(G45), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n455), .B2(new_n451), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n268), .C1(new_n455), .C2(new_n454), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OR2_X1    g0263(.A1(G250), .A2(G1698), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(G257), .B2(new_n284), .ZN(new_n465));
  INV_X1    g0265(.A(G294), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n363), .A2(new_n465), .B1(new_n466), .B2(new_n335), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n463), .B1(new_n467), .B2(new_n275), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n289), .B1(new_n459), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n459), .A2(new_n468), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n471), .B2(G190), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n442), .A2(new_n449), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n449), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n432), .A2(new_n439), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT24), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n432), .A2(new_n423), .A3(new_n439), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n474), .B1(new_n478), .B2(new_n252), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n470), .A2(new_n384), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(G179), .B2(new_n470), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n473), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G116), .ZN(new_n483));
  INV_X1    g0283(.A(new_n433), .ZN(new_n484));
  OAI22_X1  g0284(.A1(new_n443), .A2(new_n483), .B1(new_n484), .B2(new_n249), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n433), .A2(G20), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n208), .C1(G33), .C2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n252), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT20), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n487), .A2(KEYINPUT20), .A3(new_n252), .A4(new_n490), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n384), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n224), .A2(G1698), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(G257), .B2(G1698), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n363), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G303), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n278), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n275), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n456), .A2(G270), .A3(new_n340), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n503), .A2(KEYINPUT77), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(KEYINPUT77), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n502), .A2(new_n504), .A3(new_n462), .A4(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT21), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n496), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n496), .B2(new_n506), .ZN(new_n509));
  INV_X1    g0309(.A(new_n495), .ZN(new_n510));
  OAI21_X1  g0310(.A(G179), .B1(new_n510), .B2(new_n485), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n508), .A2(new_n509), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(G200), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n510), .A2(new_n485), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G190), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT74), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n284), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(new_n488), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n222), .A2(G1698), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n363), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n523), .B1(new_n527), .B2(KEYINPUT71), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT4), .B1(new_n336), .B2(new_n525), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n340), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n456), .A2(G257), .A3(new_n340), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT73), .B1(new_n533), .B2(new_n462), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n462), .A3(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n520), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n521), .A2(new_n522), .A3(new_n488), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n529), .B2(new_n530), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n527), .A2(KEYINPUT71), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n275), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n536), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(new_n534), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT74), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n538), .A2(new_n545), .A3(G200), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n249), .A2(G97), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n444), .B2(G97), .ZN(new_n548));
  XNOR2_X1  g0348(.A(G97), .B(G107), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT70), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n550), .A2(KEYINPUT6), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  MUX2_X1   g0352(.A(new_n550), .B(G97), .S(KEYINPUT6), .Z(new_n553));
  OAI211_X1 g0353(.A(new_n552), .B(G20), .C1(new_n549), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n256), .A2(G77), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n379), .B2(G107), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n548), .B1(new_n557), .B2(new_n262), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n532), .A2(new_n537), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(G190), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n546), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n292), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n542), .A2(new_n544), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n384), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n564), .A3(new_n558), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n336), .A2(new_n208), .A3(G68), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G97), .A2(G107), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(new_n430), .B1(new_n299), .B2(new_n208), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n259), .A2(KEYINPUT19), .A3(new_n489), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n566), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(new_n252), .B1(new_n250), .B2(new_n411), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n443), .A2(new_n411), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n460), .A2(G250), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n340), .A2(new_n576), .B1(new_n268), .B2(new_n450), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G238), .A2(G1698), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n222), .B2(G1698), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n434), .B1(new_n336), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n580), .B2(new_n340), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n581), .A2(G179), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n384), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n575), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n443), .A2(new_n430), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n585), .B(KEYINPUT76), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(G200), .ZN(new_n587));
  OAI211_X1 g0387(.A(G190), .B(new_n577), .C1(new_n580), .C2(new_n340), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n586), .A2(new_n573), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n519), .A2(new_n561), .A3(new_n565), .A4(new_n591), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n422), .A2(new_n482), .A3(new_n592), .ZN(G372));
  INV_X1    g0393(.A(new_n422), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n511), .A2(new_n506), .ZN(new_n595));
  INV_X1    g0395(.A(new_n509), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n496), .A2(new_n506), .A3(new_n507), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n481), .B1(new_n442), .B2(new_n449), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(KEYINPUT82), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT82), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n601), .B(new_n481), .C1(new_n442), .C2(new_n449), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n598), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n473), .A2(new_n561), .A3(new_n591), .A4(new_n565), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT83), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT83), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n603), .A2(new_n608), .A3(new_n605), .ZN(new_n609));
  INV_X1    g0409(.A(new_n565), .ZN(new_n610));
  XNOR2_X1  g0410(.A(KEYINPUT84), .B(KEYINPUT26), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n591), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT26), .B1(new_n565), .B2(new_n590), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n584), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n607), .A2(new_n609), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n594), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n329), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n325), .B1(new_n618), .B2(new_n420), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n383), .A2(new_n397), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n387), .A2(new_n389), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n295), .B1(new_n623), .B2(new_n291), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n617), .A2(new_n624), .ZN(G369));
  INV_X1    g0425(.A(new_n482), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(G213), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(G343), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n626), .B1(new_n479), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n599), .A2(new_n632), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n519), .B1(new_n514), .B2(new_n633), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n512), .B(new_n632), .C1(new_n510), .C2(new_n485), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G330), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n600), .A2(new_n602), .A3(new_n632), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n598), .A2(new_n632), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n626), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(G399));
  NAND2_X1  g0446(.A1(new_n211), .A2(new_n270), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n567), .A2(new_n430), .A3(new_n483), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n647), .A2(G1), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n215), .B2(new_n647), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT28), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT29), .B1(new_n616), .B2(new_n633), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n610), .A2(new_n654), .A3(new_n591), .ZN(new_n655));
  INV_X1    g0455(.A(new_n611), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n565), .B2(new_n590), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n655), .A2(new_n584), .A3(new_n657), .ZN(new_n658));
  OAI211_X1 g0458(.A(KEYINPUT85), .B(new_n598), .C1(new_n479), .C2(new_n481), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT85), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n599), .B2(new_n512), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n604), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT86), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI211_X1 g0464(.A(KEYINPUT86), .B(new_n604), .C1(new_n661), .C2(new_n659), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n633), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT87), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g0468(.A(KEYINPUT87), .B(new_n633), .C1(new_n664), .C2(new_n665), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n653), .B1(new_n670), .B2(KEYINPUT29), .ZN(new_n671));
  INV_X1    g0471(.A(G330), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n674));
  OAI211_X1 g0474(.A(G179), .B(new_n577), .C1(new_n580), .C2(new_n340), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n471), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n673), .B1(new_n677), .B2(new_n563), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n559), .A2(KEYINPUT30), .A3(new_n471), .A4(new_n676), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n581), .A2(new_n292), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n563), .A2(new_n470), .A3(new_n506), .A4(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(KEYINPUT31), .A3(new_n632), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT31), .B1(new_n682), .B2(new_n632), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n561), .A2(new_n565), .A3(new_n591), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n626), .A2(new_n519), .A3(new_n687), .A4(new_n633), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n672), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n671), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n652), .B1(new_n690), .B2(G1), .ZN(G364));
  XNOR2_X1  g0491(.A(new_n640), .B(KEYINPUT88), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n208), .A2(G13), .A3(G45), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT89), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n647), .A2(G1), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n692), .B(new_n697), .C1(G330), .C2(new_n639), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n217), .B1(G20), .B2(new_n384), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n208), .A2(new_n292), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G200), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT91), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G190), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  XOR2_X1   g0505(.A(KEYINPUT33), .B(G317), .Z(new_n706));
  INV_X1    g0506(.A(G322), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n701), .A2(G190), .A3(new_n289), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n705), .A2(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT92), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n703), .A2(new_n516), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G326), .ZN(new_n714));
  NOR2_X1   g0514(.A1(G190), .A2(G200), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n701), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G311), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n281), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n516), .A2(G179), .A3(G200), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n208), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n208), .A2(G179), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n516), .A3(G200), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n721), .A2(G294), .B1(new_n724), .B2(G283), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(G190), .A3(G200), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n500), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n722), .A2(new_n715), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n718), .B(new_n727), .C1(G329), .C2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n711), .A2(new_n712), .A3(new_n714), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n723), .A2(new_n223), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT32), .ZN(new_n733));
  INV_X1    g0533(.A(G159), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n732), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n489), .B2(new_n720), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n278), .B1(new_n716), .B2(new_n221), .C1(new_n202), .C2(new_n708), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n735), .A2(new_n733), .B1(new_n430), .B2(new_n726), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n713), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n740), .B1(new_n201), .B2(new_n741), .C1(new_n203), .C2(new_n705), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n700), .B1(new_n731), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n699), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n363), .A2(new_n211), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n271), .B2(new_n216), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n244), .B2(new_n271), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n211), .A2(new_n278), .ZN(new_n752));
  INV_X1    g0552(.A(G355), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n752), .A2(new_n753), .B1(G116), .B2(new_n211), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT90), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n748), .B1(new_n751), .B2(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n743), .A2(new_n756), .A3(new_n697), .ZN(new_n757));
  INV_X1    g0557(.A(new_n746), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n639), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n698), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(G396));
  INV_X1    g0561(.A(new_n697), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n614), .B1(new_n606), .B2(KEYINPUT83), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n632), .B1(new_n763), .B2(new_n609), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n420), .A2(new_n632), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n632), .B1(new_n413), .B2(new_n415), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n417), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(new_n420), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n764), .B(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n689), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n762), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  INV_X1    g0572(.A(new_n708), .ZN(new_n773));
  INV_X1    g0573(.A(new_n716), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n773), .A2(G143), .B1(new_n774), .B2(G159), .ZN(new_n775));
  INV_X1    g0575(.A(G150), .ZN(new_n776));
  INV_X1    g0576(.A(G137), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n775), .B1(new_n705), .B2(new_n776), .C1(new_n777), .C2(new_n741), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT34), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n720), .A2(new_n202), .B1(new_n726), .B2(new_n201), .ZN(new_n782));
  INV_X1    g0582(.A(G132), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n336), .B1(new_n783), .B2(new_n728), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n782), .B(new_n784), .C1(G68), .C2(new_n724), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n780), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n430), .A2(new_n723), .B1(new_n726), .B2(new_n223), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n281), .B1(new_n728), .B2(new_n717), .C1(new_n433), .C2(new_n716), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(new_n704), .C2(G283), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT93), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n720), .A2(new_n489), .B1(new_n708), .B2(new_n466), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n713), .A2(G303), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n789), .B(new_n792), .C1(new_n790), .C2(new_n791), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n700), .B1(new_n794), .B2(KEYINPUT94), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(KEYINPUT94), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n699), .A2(new_n744), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n697), .B1(new_n221), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(new_n768), .C2(new_n745), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n772), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G384));
  OAI21_X1  g0601(.A(new_n552), .B1(new_n553), .B2(new_n549), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT35), .ZN(new_n803));
  OAI211_X1 g0603(.A(G116), .B(new_n218), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n803), .B2(new_n802), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT36), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n216), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n201), .A2(G68), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n207), .B(G13), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n630), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT96), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n390), .A2(KEYINPUT95), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT95), .ZN(new_n814));
  AOI21_X1  g0614(.A(KEYINPUT16), .B1(new_n369), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n371), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n812), .B1(new_n816), .B2(new_n355), .ZN(new_n817));
  OR3_X1    g0617(.A1(new_n816), .A2(new_n812), .A3(new_n355), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n398), .A2(new_n811), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT37), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n382), .A2(new_n811), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n386), .A2(new_n396), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT97), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n818), .B(new_n817), .C1(new_n385), .C2(new_n811), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n820), .B1(new_n824), .B2(new_n396), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n819), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n819), .B(KEYINPUT38), .C1(new_n823), .C2(new_n825), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n828), .A2(KEYINPUT39), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n386), .A2(new_n396), .A3(new_n821), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(KEYINPUT37), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n386), .A2(new_n396), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n833), .A2(KEYINPUT97), .A3(new_n820), .A4(new_n821), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT97), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n822), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n832), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n821), .B1(new_n620), .B2(new_n622), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n827), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n839), .A2(new_n829), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n830), .B1(new_n840), .B2(KEYINPUT39), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n315), .A2(new_n324), .A3(new_n633), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT98), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n622), .A2(new_n811), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n324), .B(new_n632), .C1(new_n618), .C2(new_n315), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n324), .A2(new_n632), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n325), .A2(new_n329), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n616), .A2(new_n633), .A3(new_n768), .ZN(new_n852));
  INV_X1    g0652(.A(new_n765), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n828), .A2(new_n829), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n846), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n624), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n671), .B2(new_n594), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n858), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n686), .A2(new_n688), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n862), .A2(new_n768), .A3(new_n850), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT40), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n855), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n839), .A2(new_n829), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n866), .A2(new_n863), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n867), .B2(new_n864), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n422), .B1(new_n688), .B2(new_n686), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n672), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n861), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT99), .ZN(new_n873));
  INV_X1    g0673(.A(G13), .ZN(new_n874));
  OAI21_X1  g0674(.A(G1), .B1(new_n874), .B2(G20), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n873), .B(new_n875), .C1(new_n861), .C2(new_n871), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n872), .A2(KEYINPUT99), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n810), .B1(new_n876), .B2(new_n877), .ZN(G367));
  INV_X1    g0678(.A(KEYINPUT102), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n610), .A2(new_n632), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT101), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n558), .A2(new_n632), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n561), .A2(new_n565), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n626), .A3(new_n644), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT42), .Z(new_n886));
  AOI21_X1  g0686(.A(new_n610), .B1(new_n884), .B2(new_n599), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n886), .B1(new_n632), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n633), .B1(new_n586), .B2(new_n573), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT100), .Z(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n584), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n591), .B2(new_n890), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT43), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n879), .B1(new_n888), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n888), .A2(new_n879), .A3(new_n894), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(new_n893), .A3(new_n892), .A4(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n641), .A2(new_n884), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n892), .A2(new_n893), .ZN(new_n900));
  INV_X1    g0700(.A(new_n897), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n900), .B1(new_n901), .B2(new_n895), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n899), .B1(new_n898), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n647), .B(KEYINPUT41), .ZN(new_n906));
  MUX2_X1   g0706(.A(new_n636), .B(new_n626), .S(new_n644), .Z(new_n907));
  NOR2_X1   g0707(.A1(new_n907), .A2(new_n640), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n692), .B2(new_n907), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n690), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT103), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n645), .A2(new_n884), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT45), .Z(new_n914));
  NOR2_X1   g0714(.A1(new_n645), .A2(new_n884), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT44), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n914), .A2(new_n642), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n916), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n641), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n911), .A2(new_n912), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n917), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT103), .B1(new_n921), .B2(new_n910), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n906), .B1(new_n923), .B2(new_n690), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n696), .A2(G1), .A3(new_n695), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT104), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n905), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n747), .B1(new_n211), .B2(new_n411), .C1(new_n239), .C2(new_n749), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n723), .A2(new_n489), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(G107), .B2(new_n721), .ZN(new_n930));
  INV_X1    g0730(.A(new_n726), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(KEYINPUT46), .A3(G116), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n363), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(KEYINPUT105), .B(G317), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n773), .A2(G303), .B1(new_n729), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(G283), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n936), .B1(new_n937), .B2(new_n716), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT46), .B1(new_n931), .B2(new_n484), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n933), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n940), .B1(new_n466), .B2(new_n705), .C1(new_n717), .C2(new_n741), .ZN(new_n941));
  AOI22_X1  g0741(.A1(G143), .A2(new_n713), .B1(new_n704), .B2(G159), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n716), .A2(new_n201), .B1(new_n728), .B2(new_n777), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n281), .B(new_n943), .C1(G150), .C2(new_n773), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n723), .A2(new_n221), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n720), .A2(new_n203), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n945), .B(new_n946), .C1(G58), .C2(new_n931), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n942), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT47), .Z(new_n950));
  OAI211_X1 g0750(.A(new_n762), .B(new_n928), .C1(new_n950), .C2(new_n700), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n892), .A2(new_n746), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n927), .A2(new_n954), .ZN(G387));
  NAND2_X1  g0755(.A1(new_n636), .A2(new_n746), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n752), .A2(new_n649), .B1(G107), .B2(new_n211), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT106), .Z(new_n958));
  OR2_X1    g0758(.A1(new_n236), .A2(new_n271), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n258), .A2(G50), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT50), .ZN(new_n961));
  AOI211_X1 g0761(.A(G45), .B(new_n648), .C1(G68), .C2(G77), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n749), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n958), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n762), .B1(new_n964), .B2(new_n748), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n704), .A2(new_n353), .B1(G68), .B2(new_n774), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT107), .Z(new_n967));
  OAI221_X1 g0767(.A(new_n336), .B1(new_n776), .B2(new_n728), .C1(new_n201), .C2(new_n708), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n726), .A2(new_n221), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n720), .A2(new_n411), .ZN(new_n970));
  NOR4_X1   g0770(.A1(new_n968), .A2(new_n929), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n967), .B(new_n971), .C1(new_n734), .C2(new_n741), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n773), .A2(new_n935), .B1(new_n774), .B2(G303), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n705), .B2(new_n717), .C1(new_n707), .C2(new_n741), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT48), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n721), .A2(G283), .B1(new_n931), .B2(G294), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT49), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(KEYINPUT108), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n723), .A2(new_n433), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n336), .B(new_n983), .C1(G326), .C2(new_n729), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT108), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n972), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n965), .B1(new_n987), .B2(new_n699), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n909), .A2(new_n926), .B1(new_n956), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n647), .B(KEYINPUT109), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n910), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n690), .A2(new_n909), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT110), .Z(G393));
  NAND2_X1  g0794(.A1(new_n921), .A2(new_n910), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT112), .ZN(new_n996));
  INV_X1    g0796(.A(new_n990), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n920), .B2(new_n922), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT113), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n996), .A2(new_n998), .A3(KEYINPUT113), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n919), .A2(new_n917), .A3(new_n926), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n747), .B1(new_n489), .B2(new_n211), .C1(new_n247), .C2(new_n749), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n1005), .A2(new_n762), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n704), .A2(G303), .B1(new_n484), .B2(new_n721), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n281), .B1(new_n728), .B2(new_n707), .C1(new_n466), .C2(new_n716), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n732), .B(new_n1011), .C1(G283), .C2(new_n931), .ZN(new_n1012));
  AND3_X1   g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n713), .A2(G317), .B1(G311), .B2(new_n773), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT52), .Z(new_n1015));
  AOI22_X1  g0815(.A1(new_n713), .A2(G150), .B1(G159), .B2(new_n773), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT51), .Z(new_n1017));
  NAND2_X1  g0817(.A1(new_n729), .A2(G143), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1018), .B(new_n336), .C1(new_n258), .C2(new_n716), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n721), .A2(G77), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n203), .B2(new_n726), .C1(new_n430), .C2(new_n723), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1019), .B(new_n1021), .C1(G50), .C2(new_n704), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n1013), .A2(new_n1015), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1006), .B1(new_n700), .B2(new_n1023), .C1(new_n884), .C2(new_n758), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1004), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1003), .A2(new_n1026), .ZN(G390));
  NOR2_X1   g0827(.A1(new_n770), .A2(new_n422), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n592), .A2(new_n482), .A3(new_n632), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n682), .A2(new_n632), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT31), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n683), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n768), .B(G330), .C1(new_n1030), .C2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT115), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n768), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1035), .B(new_n851), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1038), .B1(new_n1039), .B2(new_n1037), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n668), .A2(new_n669), .A3(new_n853), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n767), .A2(new_n420), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT114), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n765), .B1(new_n764), .B2(new_n768), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1035), .B(new_n850), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n852), .A2(new_n853), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n1039), .A3(KEYINPUT114), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n860), .B(new_n1029), .C1(new_n1044), .C2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1035), .A2(new_n851), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1041), .A2(new_n1042), .A3(new_n850), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n843), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n840), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n841), .B1(new_n854), .B2(new_n1056), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1054), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n1058), .A2(new_n1059), .A3(new_n1054), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1052), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n1053), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1058), .A2(new_n1059), .A3(new_n1054), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n859), .B(new_n1028), .C1(new_n671), .C2(new_n594), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1062), .A2(new_n990), .A3(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n713), .A2(G283), .B1(G97), .B2(new_n774), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n223), .B2(new_n705), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT117), .Z(new_n1073));
  OAI221_X1 g0873(.A(new_n281), .B1(new_n728), .B2(new_n466), .C1(new_n708), .C2(new_n483), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1020), .B1(new_n203), .B2(new_n723), .C1(new_n430), .C2(new_n726), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(G128), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1077), .A2(new_n741), .B1(new_n705), .B2(new_n777), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n726), .A2(new_n776), .ZN(new_n1079));
  XOR2_X1   g0879(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1080));
  XNOR2_X1  g0880(.A(new_n1079), .B(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n721), .A2(G159), .B1(new_n724), .B2(G50), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n773), .A2(G132), .B1(new_n729), .B2(G125), .ZN(new_n1083));
  XOR2_X1   g0883(.A(KEYINPUT54), .B(G143), .Z(new_n1084));
  AOI21_X1  g0884(.A(new_n281), .B1(new_n774), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1078), .A2(new_n1081), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n699), .B1(new_n1076), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n797), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1088), .B(new_n762), .C1(new_n353), .C2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n841), .B2(new_n744), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1061), .A2(new_n1060), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1091), .B1(new_n1092), .B2(new_n926), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1070), .A2(new_n1093), .ZN(G378));
  NAND2_X1  g0894(.A1(new_n1069), .A2(new_n1066), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(KEYINPUT121), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT121), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1069), .A2(new_n1097), .A3(new_n1066), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n844), .A2(new_n845), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT120), .B1(new_n1100), .B2(new_n856), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n297), .A2(KEYINPUT118), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n263), .A2(new_n811), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT119), .Z(new_n1105));
  NOR2_X1   g0905(.A1(new_n297), .A2(KEYINPUT118), .ZN(new_n1106));
  OR3_X1    g0906(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1105), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1108), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n868), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n672), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n868), .A3(G330), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1101), .B(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT57), .B1(new_n1099), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1116), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1112), .B1(new_n868), .B2(G330), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1100), .B(new_n856), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1115), .B(new_n1116), .C1(new_n846), .C2(new_n857), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1122), .A2(new_n1123), .A3(KEYINPUT57), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1069), .A2(new_n1097), .A3(new_n1066), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1097), .B1(new_n1069), .B2(new_n1066), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1124), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n990), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1119), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n363), .B2(new_n270), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G97), .A2(new_n704), .B1(new_n713), .B2(G116), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n969), .B(new_n946), .C1(G58), .C2(new_n724), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n716), .A2(new_n411), .B1(new_n728), .B2(new_n937), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n708), .A2(new_n223), .ZN(new_n1135));
  NOR4_X1   g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n336), .A4(G41), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT58), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1131), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n720), .A2(new_n776), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n708), .A2(new_n1077), .B1(new_n716), .B2(new_n777), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(new_n931), .C2(new_n1084), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n713), .A2(G125), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(new_n705), .C2(new_n783), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(KEYINPUT59), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n724), .A2(G159), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G33), .B(G41), .C1(new_n729), .C2(G124), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1144), .A2(KEYINPUT59), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1139), .B1(new_n1138), .B2(new_n1137), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n699), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n697), .B1(new_n201), .B2(new_n797), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(new_n1112), .C2(new_n745), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n1118), .B2(new_n926), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1129), .A2(new_n1155), .ZN(G375));
  XOR2_X1   g0956(.A(new_n926), .B(KEYINPUT122), .Z(new_n1157));
  NAND2_X1  g0957(.A1(new_n1068), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n697), .B1(new_n203), .B2(new_n797), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G294), .A2(new_n713), .B1(new_n704), .B2(new_n484), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n278), .B1(new_n773), .B2(G283), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G107), .A2(new_n774), .B1(new_n729), .B2(G303), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n945), .B(new_n970), .C1(G97), .C2(new_n931), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT123), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G132), .A2(new_n713), .B1(new_n704), .B2(new_n1084), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n716), .A2(new_n776), .B1(new_n728), .B2(new_n1077), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G137), .B2(new_n773), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n363), .B1(G58), .B2(new_n724), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n721), .A2(G50), .B1(new_n931), .B2(G159), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1164), .A2(KEYINPUT123), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1165), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1159), .B1(new_n700), .B2(new_n1173), .C1(new_n850), .C2(new_n745), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1158), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n906), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1052), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1176), .B1(new_n1178), .B2(new_n1179), .ZN(G381));
  AND3_X1   g0980(.A1(new_n1070), .A2(KEYINPUT124), .A3(new_n1093), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT124), .B1(new_n1070), .B2(new_n1093), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(G375), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n926), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n923), .A2(new_n690), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n906), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n953), .B1(new_n1188), .B2(new_n905), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1025), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1185), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(G407));
  NAND2_X1  g0992(.A1(new_n631), .A2(G213), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1185), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(G407), .A2(G213), .A3(new_n1195), .ZN(G409));
  NAND2_X1  g0996(.A1(G390), .A2(new_n1189), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(G387), .A2(new_n1190), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(G393), .B(new_n760), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(G378), .B(new_n1155), .C1(new_n1119), .C2(new_n1128), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1118), .B(new_n1177), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1122), .A2(new_n1123), .A3(new_n1157), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1207), .A2(new_n1153), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1183), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1194), .B1(new_n1205), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1179), .A2(KEYINPUT125), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT60), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1212), .A2(KEYINPUT60), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1052), .A2(new_n990), .ZN(new_n1217));
  OAI211_X1 g1017(.A(G384), .B(new_n1176), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1179), .A2(KEYINPUT125), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT60), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1217), .B1(new_n1221), .B2(new_n1213), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n800), .B1(new_n1222), .B2(new_n1175), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1218), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1211), .A2(KEYINPUT62), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT62), .B1(new_n1211), .B2(new_n1225), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT126), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1211), .A2(new_n1225), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT62), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1228), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1205), .A2(new_n1210), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1193), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1194), .A2(G2897), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1218), .A2(new_n1223), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1218), .B2(new_n1223), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT61), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1232), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1204), .B1(new_n1229), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT63), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1204), .B1(new_n1242), .B2(new_n1230), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1211), .A2(KEYINPUT63), .A3(new_n1225), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n1239), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1241), .A2(new_n1245), .ZN(G405));
  INV_X1    g1046(.A(new_n1203), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1200), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1224), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1202), .A2(new_n1225), .A3(new_n1203), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1184), .B1(new_n1129), .B2(new_n1155), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT127), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1205), .A2(KEYINPUT127), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1254), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1251), .B(new_n1256), .ZN(G402));
endmodule


