//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT67), .B(G116), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G119), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT2), .B(G113), .Z(new_n193));
  AOI21_X1  g007(.A(new_n188), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G116), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(G119), .ZN(new_n198));
  INV_X1    g012(.A(new_n190), .ZN(new_n199));
  AND4_X1   g013(.A1(new_n188), .A2(new_n193), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  OAI22_X1  g014(.A1(new_n194), .A2(new_n200), .B1(new_n192), .B2(new_n193), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n201), .B(KEYINPUT71), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT69), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n206), .A2(new_n209), .A3(new_n212), .A4(new_n207), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT64), .A2(G143), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(G146), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G143), .ZN(new_n221));
  AND2_X1   g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n220), .A2(G143), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT64), .B(G143), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(new_n220), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G128), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n203), .B1(new_n214), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT64), .A2(G143), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT64), .A2(G143), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n220), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n224), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n227), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n211), .A2(new_n213), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(KEYINPUT69), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n219), .A2(new_n221), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT65), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n219), .A2(new_n243), .A3(new_n221), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n233), .A2(new_n234), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(KEYINPUT66), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n242), .A2(new_n244), .B1(new_n245), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n207), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n205), .A2(G137), .ZN(new_n254));
  OAI21_X1  g068(.A(G131), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n213), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n229), .B(new_n238), .C1(new_n252), .C2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n202), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n202), .A2(new_n257), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n187), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n236), .A2(new_n237), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n252), .B2(new_n256), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n187), .B1(new_n202), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G101), .ZN(new_n267));
  INV_X1    g081(.A(G237), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G210), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n267), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n266), .A2(KEYINPUT29), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n263), .A2(new_n201), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n264), .B(new_n278), .C1(new_n259), .C2(new_n187), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(new_n273), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT70), .B1(new_n257), .B2(new_n281), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n214), .A2(new_n228), .A3(new_n203), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT69), .B1(new_n236), .B2(new_n237), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n242), .A2(new_n244), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n245), .A2(new_n251), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(new_n255), .A3(new_n213), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n285), .A2(new_n286), .A3(new_n290), .A4(KEYINPUT30), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n282), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n263), .A2(new_n281), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n201), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n274), .B1(new_n296), .B2(new_n259), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n280), .A2(KEYINPUT29), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G472), .B1(new_n277), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n279), .A2(new_n273), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n274), .B1(new_n202), .B2(new_n257), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n296), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n294), .B1(new_n282), .B2(new_n291), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT73), .B1(new_n306), .B2(new_n303), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n301), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT31), .B1(new_n296), .B2(new_n304), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n300), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT32), .ZN(new_n311));
  NOR2_X1   g125(.A1(G472), .A2(G902), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n312), .B(KEYINPUT74), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n310), .B2(new_n314), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n299), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G217), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(G234), .B2(new_n276), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT22), .B(G137), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n320), .B(new_n321), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n239), .A2(G119), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G119), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n249), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT24), .B(G110), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G110), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT66), .B(G128), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT23), .A3(G119), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT23), .B1(new_n239), .B2(G119), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(new_n324), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n330), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G125), .ZN(new_n338));
  INV_X1    g152(.A(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G140), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT75), .ZN(new_n341));
  OR3_X1    g155(.A1(new_n339), .A2(KEYINPUT75), .A3(G140), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT16), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT16), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G146), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n220), .B1(new_n343), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n336), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n327), .A2(new_n328), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n332), .A2(new_n334), .A3(new_n330), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n346), .A2(G146), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n338), .A2(new_n340), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n220), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n349), .A2(new_n350), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n350), .B1(new_n349), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n323), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n323), .B1(new_n349), .B2(new_n357), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT25), .B1(new_n363), .B2(new_n276), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n365), .B(G902), .C1(new_n360), .C2(new_n362), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n319), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n319), .A2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G104), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT3), .B1(new_n372), .B2(G107), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n374));
  INV_X1    g188(.A(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n372), .A2(G107), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G101), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT80), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n378), .A2(new_n382), .A3(new_n379), .A4(G101), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n378), .A2(G101), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT79), .B(G101), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(new_n376), .A3(new_n373), .A4(new_n377), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(KEYINPUT4), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n236), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT81), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n381), .A2(new_n383), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n236), .A4(new_n388), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT83), .B1(new_n375), .B2(G104), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT82), .B1(new_n372), .B2(G107), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n372), .A3(G107), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n375), .A3(G104), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n395), .A2(new_n396), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G101), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT10), .A3(new_n387), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n289), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT84), .B1(new_n252), .B2(new_n403), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(G146), .B1(new_n217), .B2(new_n218), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT1), .ZN(new_n410));
  OAI21_X1  g224(.A(G128), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n219), .A2(new_n221), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n287), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n402), .A2(new_n387), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n394), .A2(new_n408), .A3(new_n214), .A4(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n242), .A2(new_n244), .B1(new_n411), .B2(new_n412), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT86), .B1(new_n421), .B2(new_n415), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n287), .A2(new_n288), .A3(new_n415), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n252), .A2(new_n425), .A3(new_n415), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n214), .A2(KEYINPUT85), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT12), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n252), .A2(new_n415), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n417), .A2(KEYINPUT86), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT12), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n426), .A4(new_n427), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n420), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n269), .A2(G227), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT78), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G140), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n394), .A2(new_n408), .A3(new_n419), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n237), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n438), .A3(new_n420), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(G469), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G469), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(new_n276), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT87), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n450), .A3(new_n447), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n420), .A2(new_n429), .A3(new_n433), .A4(new_n438), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n438), .B1(new_n442), .B2(new_n420), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n445), .B(new_n276), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G952), .ZN(new_n457));
  AOI211_X1 g271(.A(G953), .B(new_n457), .C1(G234), .C2(G237), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(G898), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT96), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI211_X1 g275(.A(new_n276), .B(new_n269), .C1(G234), .C2(G237), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G214), .B1(G237), .B2(G902), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n252), .A2(new_n339), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n228), .A2(G125), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G224), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G953), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT7), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n201), .A2(new_n391), .A3(new_n388), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n193), .A2(new_n198), .A3(new_n199), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT68), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n192), .A2(KEYINPUT5), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n477), .B(G113), .C1(KEYINPUT5), .C2(new_n199), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n478), .A3(new_n416), .ZN(new_n479));
  XNOR2_X1  g293(.A(G110), .B(G122), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n466), .A2(KEYINPUT7), .A3(new_n471), .A4(new_n467), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n473), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n480), .B(KEYINPUT8), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n416), .B1(new_n476), .B2(new_n478), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n479), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI211_X1 g301(.A(KEYINPUT88), .B(new_n416), .C1(new_n476), .C2(new_n478), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(G902), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n474), .A2(new_n479), .ZN(new_n491));
  INV_X1    g305(.A(new_n480), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(KEYINPUT6), .A3(new_n481), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n468), .B(new_n470), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n496), .A3(new_n492), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G210), .B1(G237), .B2(G902), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n490), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n490), .B2(new_n498), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n464), .B(new_n465), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G478), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT9), .B(G234), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n506), .A2(new_n318), .A3(G953), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n231), .A2(new_n232), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G128), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT13), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n331), .A2(G143), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(KEYINPUT13), .A3(G128), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n515), .A2(KEYINPUT94), .A3(G134), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT94), .B1(new_n515), .B2(G134), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n513), .A3(new_n205), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n191), .A2(G122), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n189), .A2(G122), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n375), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n375), .B1(new_n519), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n516), .A2(new_n517), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n518), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n205), .B1(new_n510), .B2(new_n513), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n519), .A2(KEYINPUT14), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT95), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n519), .A2(KEYINPUT14), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT95), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n519), .A2(new_n532), .A3(KEYINPUT14), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n530), .A2(new_n531), .A3(new_n533), .A4(new_n520), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n528), .B1(G107), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n508), .B1(new_n525), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n515), .A2(G134), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n524), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n515), .A2(KEYINPUT94), .A3(G134), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n534), .A2(G107), .ZN(new_n543));
  INV_X1    g357(.A(new_n528), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n545), .A3(new_n507), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n536), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n505), .B1(new_n547), .B2(new_n276), .ZN(new_n548));
  AOI211_X1 g362(.A(G902), .B(new_n504), .C1(new_n536), .C2(new_n546), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n347), .A2(new_n348), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n268), .A2(new_n269), .A3(G214), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n217), .A3(new_n218), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n268), .A2(new_n269), .A3(G143), .A4(G214), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n212), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT17), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n553), .A2(new_n212), .A3(new_n554), .ZN(new_n557));
  OR3_X1    g371(.A1(new_n557), .A2(new_n555), .A3(KEYINPUT17), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G113), .B(G122), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(new_n372), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n341), .A2(new_n342), .A3(G146), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n356), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n553), .A2(new_n554), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT18), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n564), .A2(new_n565), .A3(new_n212), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n553), .A2(new_n554), .B1(KEYINPUT18), .B2(G131), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n559), .A2(new_n561), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n561), .B1(new_n559), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n276), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT93), .B(G475), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT90), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n557), .B2(new_n555), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n564), .A2(G131), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n553), .A2(new_n212), .A3(new_n554), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(KEYINPUT90), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT19), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n341), .B2(new_n342), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n355), .A2(KEYINPUT19), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n220), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n576), .A2(new_n579), .A3(new_n354), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(KEYINPUT91), .A3(new_n568), .ZN(new_n585));
  INV_X1    g399(.A(new_n561), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT91), .B1(new_n584), .B2(new_n568), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n569), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT20), .ZN(new_n591));
  NOR2_X1   g405(.A1(G475), .A2(G902), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n589), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n592), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n584), .A2(new_n568), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT91), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n586), .A3(new_n585), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n598), .B2(new_n569), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n600));
  OAI21_X1  g414(.A(new_n593), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n590), .B1(new_n599), .B2(new_n591), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n550), .B(new_n574), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n502), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(G221), .ZN(new_n605));
  INV_X1    g419(.A(new_n506), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n606), .B2(new_n276), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT77), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n456), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n317), .A2(new_n371), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT97), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(new_n386), .ZN(G3));
  INV_X1    g427(.A(new_n300), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n302), .B1(new_n296), .B2(new_n304), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n303), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT31), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n309), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT98), .B1(new_n619), .B2(G902), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n310), .A2(new_n621), .A3(new_n276), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(G472), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n420), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n390), .A2(new_n393), .B1(new_n417), .B2(new_n418), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n214), .B1(new_n625), .B2(new_n408), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n439), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n627), .B2(new_n452), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n448), .A2(KEYINPUT87), .B1(new_n628), .B2(new_n445), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n370), .B(new_n608), .C1(new_n629), .C2(new_n451), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n310), .A2(new_n314), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n623), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n574), .B1(new_n601), .B2(new_n602), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT99), .B1(new_n542), .B2(new_n545), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n546), .A3(new_n536), .ZN(new_n637));
  INV_X1    g451(.A(new_n546), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n507), .B1(new_n542), .B2(new_n545), .ZN(new_n639));
  OAI22_X1  g453(.A1(new_n638), .A2(new_n639), .B1(new_n634), .B2(new_n635), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n503), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n547), .A2(new_n503), .A3(new_n276), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n503), .B2(new_n276), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n633), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n502), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n632), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  XNOR2_X1  g463(.A(new_n574), .B(KEYINPUT100), .ZN(new_n650));
  INV_X1    g464(.A(new_n550), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n599), .B(new_n600), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n502), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n632), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT101), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT35), .B(G107), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  INV_X1    g472(.A(new_n359), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n349), .A2(new_n350), .A3(new_n357), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n323), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n368), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n367), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n622), .A2(G472), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n621), .B1(new_n310), .B2(new_n276), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n631), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n623), .A2(KEYINPUT102), .A3(new_n631), .A4(new_n666), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n610), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  AOI21_X1  g489(.A(new_n608), .B1(new_n629), .B2(new_n451), .ZN(new_n676));
  INV_X1    g490(.A(new_n465), .ZN(new_n677));
  INV_X1    g491(.A(new_n501), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n490), .A2(new_n498), .A3(new_n499), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n666), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n458), .B1(new_n462), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n650), .A2(new_n651), .A3(new_n652), .A4(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n317), .A2(new_n676), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  NAND2_X1  g502(.A1(new_n305), .A2(new_n307), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n274), .B1(new_n259), .B2(new_n260), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n276), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G472), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n315), .B2(new_n316), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n678), .A2(new_n679), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT38), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n633), .A2(new_n651), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(new_n677), .A3(new_n666), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n693), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n683), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n676), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT103), .Z(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n698), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n225), .ZN(G45));
  AND3_X1   g519(.A1(new_n633), .A2(new_n644), .A3(new_n684), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n681), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n317), .A2(new_n708), .A3(new_n676), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  NOR2_X1   g524(.A1(new_n628), .A2(new_n445), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n607), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n455), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n317), .A2(new_n371), .A3(new_n646), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n317), .A2(new_n371), .A3(new_n654), .A4(new_n715), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  NOR2_X1   g534(.A1(new_n714), .A2(new_n681), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n603), .A2(new_n463), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n317), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  XOR2_X1   g538(.A(KEYINPUT104), .B(G472), .Z(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n310), .B2(new_n276), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n617), .A2(new_n618), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n266), .A2(new_n274), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n313), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n465), .B1(new_n500), .B2(new_n501), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n714), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n696), .A2(new_n463), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n731), .A2(new_n733), .A3(new_n371), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT105), .B(G122), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G24));
  NAND3_X1  g551(.A1(new_n731), .A2(new_n721), .A3(new_n706), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  OAI21_X1  g553(.A(KEYINPUT32), .B1(new_n619), .B2(new_n313), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n370), .B1(new_n742), .B2(new_n299), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n500), .A2(new_n501), .A3(new_n677), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n633), .A3(new_n644), .A4(new_n684), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n455), .A2(new_n447), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n440), .A2(new_n747), .A3(new_n443), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n442), .A2(KEYINPUT106), .A3(new_n438), .A4(new_n420), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n445), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n713), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT42), .B1(new_n743), .B2(new_n752), .ZN(new_n753));
  AND4_X1   g567(.A1(KEYINPUT42), .A2(new_n317), .A3(new_n371), .A4(new_n752), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n212), .ZN(G33));
  INV_X1    g570(.A(new_n744), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n751), .A2(new_n685), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n743), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n444), .B1(new_n762), .B2(new_n445), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT107), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n748), .A2(new_n749), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT45), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n761), .B1(new_n768), .B2(new_n446), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(KEYINPUT46), .A3(new_n447), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n455), .A3(new_n770), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(new_n713), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n623), .A2(new_n631), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n633), .A2(new_n641), .A3(new_n643), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT43), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n666), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT44), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n744), .B(KEYINPUT108), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n772), .A2(new_n777), .A3(new_n699), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  XNOR2_X1  g594(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n772), .B(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n317), .A2(new_n371), .A3(new_n745), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(KEYINPUT110), .B(G140), .Z(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G42));
  NOR2_X1   g600(.A1(new_n693), .A2(new_n370), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n695), .A2(new_n608), .A3(new_n677), .ZN(new_n788));
  INV_X1    g602(.A(new_n455), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT49), .B1(new_n711), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n774), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n711), .A2(new_n789), .A3(KEYINPUT49), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n715), .A2(new_n458), .A3(new_n744), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n775), .ZN(new_n796));
  INV_X1    g610(.A(new_n743), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT48), .Z(new_n799));
  AND2_X1   g613(.A1(new_n787), .A2(new_n795), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n633), .A3(new_n644), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n371), .A2(new_n775), .A3(new_n458), .A4(new_n731), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n457), .B(G953), .C1(new_n802), .C2(new_n733), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n695), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n802), .A2(new_n677), .A3(new_n805), .A4(new_n715), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT50), .Z(new_n807));
  NOR2_X1   g621(.A1(new_n633), .A2(new_n644), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n800), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n308), .A2(new_n309), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n314), .B1(new_n810), .B2(new_n728), .ZN(new_n811));
  AOI21_X1  g625(.A(G902), .B1(new_n727), .B2(new_n300), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n666), .B(new_n811), .C1(new_n812), .C2(new_n725), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n807), .B(new_n809), .C1(new_n813), .C2(new_n796), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n711), .A2(new_n789), .A3(new_n609), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n782), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n802), .A2(new_n778), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n804), .B1(new_n818), .B2(KEYINPUT51), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(KEYINPUT51), .B2(new_n818), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n456), .A2(new_n609), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n742), .B2(new_n299), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n707), .A2(new_n681), .A3(new_n714), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n822), .A2(new_n686), .B1(new_n823), .B2(new_n731), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n680), .A2(new_n651), .A3(new_n633), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n361), .B1(new_n661), .B2(new_n323), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n365), .B1(new_n827), .B2(G902), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n363), .A2(KEYINPUT25), .A3(new_n276), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n830), .A2(new_n319), .B1(new_n368), .B2(new_n664), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n684), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n826), .A2(new_n832), .A3(new_n751), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n693), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n824), .A2(new_n825), .A3(new_n709), .A4(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n709), .A2(new_n687), .A3(new_n834), .A4(new_n738), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n835), .A2(new_n837), .A3(KEYINPUT113), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT113), .B1(new_n835), .B2(new_n837), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n623), .A2(new_n630), .A3(new_n631), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n651), .B(new_n574), .C1(new_n602), .C2(new_n601), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n502), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT111), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n646), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT111), .B1(new_n645), .B2(new_n502), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n611), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n610), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n669), .B2(new_n670), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n849), .B1(new_n672), .B2(new_n851), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n753), .A2(new_n754), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n716), .A2(new_n719), .A3(new_n723), .A4(new_n735), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT112), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n765), .A2(G469), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n446), .B1(new_n628), .B2(new_n445), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n607), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n706), .A3(new_n744), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n856), .B1(new_n813), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n731), .A2(new_n752), .A3(KEYINPUT112), .A4(new_n666), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n650), .A2(new_n550), .A3(new_n652), .A4(new_n684), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n864), .A2(new_n757), .A3(new_n831), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n822), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n863), .A2(new_n759), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n852), .A2(new_n853), .A3(new_n855), .A4(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT53), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n835), .A2(new_n837), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n841), .A2(new_n869), .B1(new_n872), .B2(KEYINPUT53), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n868), .B2(new_n870), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n846), .A2(new_n847), .ZN(new_n879));
  INV_X1    g693(.A(new_n844), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n632), .A2(new_n881), .B1(new_n743), .B2(new_n610), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n673), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n863), .A2(new_n759), .A3(new_n866), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n867), .A2(KEYINPUT114), .A3(new_n673), .A4(new_n882), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n755), .A2(new_n854), .A3(new_n875), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n876), .B(new_n877), .C1(new_n840), .C2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT115), .B1(new_n874), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n874), .A2(KEYINPUT115), .A3(new_n889), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n820), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(G952), .A2(G953), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n794), .B1(new_n892), .B2(new_n893), .ZN(G75));
  OAI21_X1  g708(.A(new_n876), .B1(new_n840), .B2(new_n888), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n895), .A2(G902), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(G210), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n896), .B2(G210), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n494), .A2(new_n497), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n495), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT55), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n899), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n897), .A2(new_n900), .A3(new_n898), .A4(new_n904), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n269), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n906), .A2(KEYINPUT117), .A3(new_n907), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(G51));
  XNOR2_X1  g728(.A(new_n446), .B(KEYINPUT57), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n895), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT119), .B1(new_n895), .B2(KEYINPUT54), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n840), .A2(new_n888), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n919), .A2(KEYINPUT118), .A3(new_n877), .A4(new_n876), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT118), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n889), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n915), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n627), .A2(new_n452), .ZN(new_n927));
  OAI211_X1 g741(.A(KEYINPUT120), .B(new_n915), .C1(new_n918), .C2(new_n923), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n896), .A2(new_n768), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n908), .B1(new_n929), .B2(new_n930), .ZN(G54));
  AND3_X1   g745(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n909), .B1(new_n932), .B2(new_n589), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n589), .B2(new_n932), .ZN(G60));
  NAND2_X1  g748(.A1(new_n637), .A2(new_n640), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n503), .A2(new_n276), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT59), .Z(new_n938));
  OAI211_X1 g752(.A(new_n936), .B(new_n938), .C1(new_n918), .C2(new_n923), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n909), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n891), .B2(new_n890), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n935), .B2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT60), .Z(new_n944));
  AND2_X1   g758(.A1(new_n895), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n908), .B1(new_n945), .B2(new_n664), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n827), .B(KEYINPUT121), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT61), .Z(G66));
  NAND2_X1  g763(.A1(new_n852), .A2(new_n855), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n269), .ZN(new_n951));
  OAI21_X1  g765(.A(G953), .B1(new_n461), .B2(new_n469), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT122), .Z(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT123), .ZN(new_n955));
  INV_X1    g769(.A(G898), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n902), .B1(new_n956), .B2(G953), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n955), .B(new_n957), .ZN(G69));
  NAND2_X1  g772(.A1(new_n292), .A2(new_n293), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n581), .A2(new_n582), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n959), .B(new_n960), .Z(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(G900), .B2(G953), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n797), .A2(new_n826), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n772), .A2(new_n699), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT125), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n824), .A2(new_n709), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n853), .A2(new_n966), .A3(new_n759), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n965), .A2(new_n784), .A3(new_n779), .A4(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n962), .B1(new_n968), .B2(G953), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n704), .A2(new_n966), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n757), .B1(new_n645), .B2(new_n843), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n701), .A2(new_n743), .A3(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n973), .A2(new_n779), .A3(new_n784), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n269), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n961), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n970), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n982), .B(new_n969), .C1(new_n978), .C2(KEYINPUT124), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n978), .A2(KEYINPUT124), .ZN(new_n984));
  OAI22_X1  g798(.A1(new_n980), .A2(new_n982), .B1(new_n983), .B2(new_n984), .ZN(G72));
  XOR2_X1   g799(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n986));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n976), .B2(new_n950), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n989), .B(new_n274), .C1(new_n258), .C2(new_n306), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n873), .B(new_n988), .C1(new_n689), .C2(new_n297), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n988), .B1(new_n968), .B2(new_n950), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n992), .A2(new_n273), .A3(new_n259), .A4(new_n296), .ZN(new_n993));
  AND4_X1   g807(.A1(new_n909), .A2(new_n990), .A3(new_n991), .A4(new_n993), .ZN(G57));
endmodule


