//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1193, new_n1194, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(G20), .A3(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT64), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n235), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G351));
  OAI21_X1  g0050(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n209), .A2(G33), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n251), .B1(new_n252), .B2(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n217), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n208), .B2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G50), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n260), .B(new_n262), .C1(G50), .C2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT9), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n218), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n266), .ZN(new_n272));
  INV_X1    g0072(.A(G226), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n280), .A2(G223), .B1(new_n283), .B2(G77), .ZN(new_n284));
  INV_X1    g0084(.A(G222), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n278), .A2(new_n279), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n275), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n274), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G200), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(G190), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n265), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n264), .B1(new_n290), .B2(G169), .ZN(new_n296));
  INV_X1    g0096(.A(G179), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G41), .ZN(new_n300));
  INV_X1    g0100(.A(G45), .ZN(new_n301));
  AOI21_X1  g0101(.A(G1), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n289), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n268), .B1(new_n303), .B2(G244), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT66), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n280), .A2(G238), .B1(new_n283), .B2(G107), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n286), .A2(G232), .A3(new_n275), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n306), .B(new_n307), .C1(new_n271), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G200), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n311), .ZN(new_n314));
  XOR2_X1   g0114(.A(KEYINPUT8), .B(G58), .Z(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n253), .B1(G20), .B2(G77), .ZN(new_n316));
  XOR2_X1   g0116(.A(KEYINPUT15), .B(G87), .Z(new_n317));
  INV_X1    g0117(.A(KEYINPUT67), .ZN(new_n318));
  INV_X1    g0118(.A(new_n255), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT15), .B(G87), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT67), .B1(new_n321), .B2(new_n255), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n316), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n259), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT68), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n263), .A2(G77), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n261), .B2(G77), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n314), .A2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n311), .A2(G179), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n311), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n329), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n295), .A2(new_n299), .A3(new_n330), .A4(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n269), .B1(new_n272), .B2(new_n222), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n286), .A2(G232), .A3(G1698), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(new_n287), .C2(new_n273), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n336), .B1(new_n339), .B2(new_n289), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n340), .A2(new_n341), .ZN(new_n343));
  OAI21_X1  g0143(.A(G169), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n344), .A2(KEYINPUT14), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(KEYINPUT14), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G179), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n345), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n319), .A2(G77), .B1(G20), .B2(new_n221), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n201), .B2(new_n254), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n353), .A2(new_n259), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n354), .A2(KEYINPUT11), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(KEYINPUT11), .ZN(new_n356));
  OR3_X1    g0156(.A1(new_n263), .A2(KEYINPUT12), .A3(G68), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT12), .B1(new_n263), .B2(G68), .ZN(new_n358));
  AOI22_X1  g0158(.A1(G68), .A2(new_n261), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT71), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n351), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(G200), .B1(new_n342), .B2(new_n343), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT70), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(KEYINPUT70), .B(G200), .C1(new_n342), .C2(new_n343), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n360), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n349), .A2(G190), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT7), .B1(new_n286), .B2(G20), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT7), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n283), .A2(new_n373), .A3(new_n209), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(G68), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT72), .B1(new_n254), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT72), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n253), .A2(new_n379), .A3(G159), .ZN(new_n380));
  XNOR2_X1  g0180(.A(G58), .B(G68), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n378), .A2(new_n380), .B1(G20), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n375), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n376), .B1(new_n375), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n259), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n256), .B1(new_n208), .B2(G20), .ZN(new_n386));
  INV_X1    g0186(.A(new_n263), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n259), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n386), .A2(new_n388), .B1(new_n387), .B2(new_n256), .ZN(new_n389));
  NOR2_X1   g0189(.A1(G223), .A2(G1698), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n273), .B2(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n286), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n271), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n269), .B1(new_n272), .B2(new_n237), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n291), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n394), .A2(new_n395), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n396), .A2(KEYINPUT73), .B1(new_n397), .B2(new_n313), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n268), .B1(new_n303), .B2(G232), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n391), .A2(new_n286), .B1(G33), .B2(G87), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n399), .B1(new_n271), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT73), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n401), .A2(new_n402), .A3(G190), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n385), .B(new_n389), .C1(new_n398), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n394), .A2(new_n395), .A3(G179), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n332), .B2(new_n401), .ZN(new_n408));
  INV_X1    g0208(.A(new_n259), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n375), .A2(new_n382), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n375), .A2(new_n376), .A3(new_n382), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n389), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n408), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT18), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n408), .B(new_n417), .C1(new_n413), .C2(new_n414), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n397), .A2(KEYINPUT73), .A3(new_n313), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n402), .B1(new_n401), .B2(new_n291), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n401), .A2(G190), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n422), .A2(KEYINPUT17), .A3(new_n385), .A4(new_n389), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n406), .A2(new_n416), .A3(new_n418), .A4(new_n423), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n335), .A2(new_n371), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT78), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT5), .B(G41), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n301), .A2(G1), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n428), .A2(new_n429), .B1(new_n218), .B2(new_n270), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G257), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n208), .A2(G45), .ZN(new_n432));
  OR2_X1    g0232(.A1(KEYINPUT5), .A2(G41), .ZN(new_n433));
  NAND2_X1  g0233(.A1(KEYINPUT5), .A2(G41), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n267), .B1(new_n218), .B2(new_n270), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT77), .ZN(new_n439));
  OAI211_X1 g0239(.A(G244), .B(new_n275), .C1(new_n281), .C2(new_n282), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT76), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  OAI211_X1 g0245(.A(G250), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT4), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n445), .B(new_n446), .C1(new_n440), .C2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n444), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n439), .B1(new_n450), .B2(new_n271), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n440), .A2(new_n442), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT76), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n440), .A2(new_n447), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n446), .A2(new_n445), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n443), .A4(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(KEYINPUT77), .A3(new_n289), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n438), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n427), .B1(new_n458), .B2(new_n291), .ZN(new_n459));
  INV_X1    g0259(.A(new_n438), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n456), .A2(KEYINPUT77), .A3(new_n289), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT77), .B1(new_n456), .B2(new_n289), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(KEYINPUT78), .A3(G200), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n372), .A2(G107), .A3(new_n374), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT74), .ZN(new_n466));
  INV_X1    g0266(.A(G107), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(KEYINPUT6), .A3(G97), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n467), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n205), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(KEYINPUT6), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT74), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n372), .A2(new_n374), .A3(new_n474), .A4(G107), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n466), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n259), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n387), .A2(new_n469), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n208), .A2(G33), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n263), .A2(new_n479), .A3(new_n217), .A4(new_n258), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n480), .B2(new_n469), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n460), .B1(new_n450), .B2(new_n271), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n313), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n459), .A2(new_n464), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n481), .B1(new_n476), .B2(new_n259), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n332), .B2(new_n484), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n297), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n430), .A2(G270), .B1(new_n435), .B2(new_n436), .ZN(new_n493));
  OAI211_X1 g0293(.A(G264), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n494));
  OAI211_X1 g0294(.A(G257), .B(new_n275), .C1(new_n281), .C2(new_n282), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n278), .A2(G303), .A3(new_n279), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n289), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G116), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n387), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n409), .A2(G116), .A3(new_n263), .A4(new_n479), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n258), .A2(new_n217), .B1(G20), .B2(new_n500), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n445), .B(new_n209), .C1(G33), .C2(new_n469), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n503), .A2(KEYINPUT20), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT20), .B1(new_n503), .B2(new_n504), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n501), .B(new_n502), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n499), .A2(new_n507), .A3(KEYINPUT21), .A4(G169), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT81), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n499), .A2(G169), .A3(new_n507), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT21), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n332), .B1(new_n493), .B2(new_n498), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT81), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT21), .A4(new_n507), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n493), .A2(new_n498), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(G179), .A3(new_n507), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n509), .A2(new_n512), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(G190), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n507), .B1(new_n499), .B2(G200), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n480), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n387), .A2(KEYINPUT25), .A3(new_n467), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT25), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n263), .B2(G107), .ZN(new_n527));
  AOI22_X1  g0327(.A1(G107), .A2(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT24), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n467), .A2(KEYINPUT23), .A3(G20), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT23), .B1(new_n467), .B2(G20), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n530), .A2(new_n531), .B1(G20), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n209), .B(G87), .C1(new_n281), .C2(new_n282), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT22), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n286), .A2(new_n536), .A3(new_n209), .A4(G87), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT82), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n529), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n533), .ZN(new_n541));
  AOI21_X1  g0341(.A(G20), .B1(new_n278), .B2(new_n279), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n536), .B1(new_n542), .B2(G87), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n534), .A2(KEYINPUT22), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT82), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(KEYINPUT82), .A3(new_n529), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n259), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n528), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(G250), .B(new_n275), .C1(new_n281), .C2(new_n282), .ZN(new_n551));
  OAI211_X1 g0351(.A(G257), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n552));
  INV_X1    g0352(.A(G294), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n551), .B(new_n552), .C1(new_n277), .C2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(KEYINPUT83), .A3(new_n289), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n428), .A2(new_n429), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(G264), .A3(new_n271), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n437), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT83), .B1(new_n554), .B2(new_n289), .ZN(new_n559));
  OAI21_X1  g0359(.A(G169), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(KEYINPUT84), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT84), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n430), .A2(new_n562), .A3(G264), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n554), .A2(new_n289), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n564), .A2(G179), .A3(new_n437), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n550), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n540), .A2(new_n546), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n259), .A3(new_n548), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n558), .A2(G190), .A3(new_n559), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n565), .A2(new_n561), .A3(new_n437), .A4(new_n563), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n572), .A2(new_n291), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n570), .B(new_n528), .C1(new_n571), .C2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G238), .B(new_n275), .C1(new_n281), .C2(new_n282), .ZN(new_n575));
  OAI211_X1 g0375(.A(G244), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n532), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n289), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n429), .A2(new_n224), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(new_n271), .B1(G274), .B2(new_n429), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n297), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT79), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n317), .A2(new_n263), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n209), .B1(new_n338), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(G87), .B2(new_n206), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n209), .B(G68), .C1(new_n281), .C2(new_n282), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n255), .B2(new_n469), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n584), .B1(new_n590), .B2(new_n259), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT80), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n524), .B2(new_n317), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n480), .A2(KEYINPUT80), .A3(new_n321), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n578), .A2(KEYINPUT79), .A3(new_n297), .A4(new_n580), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n578), .A2(new_n580), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n332), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n583), .A2(new_n595), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(G200), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n480), .A2(new_n223), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n584), .B(new_n601), .C1(new_n590), .C2(new_n259), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n600), .B(new_n602), .C1(new_n313), .C2(new_n597), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n523), .A2(new_n568), .A3(new_n574), .A4(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n426), .A2(new_n492), .A3(new_n605), .ZN(G372));
  INV_X1    g0406(.A(new_n299), .ZN(new_n607));
  INV_X1    g0407(.A(new_n334), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n370), .A2(new_n608), .B1(new_n351), .B2(new_n361), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n406), .A2(new_n423), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n416), .B(new_n418), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n607), .B1(new_n611), .B2(new_n295), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n602), .B1(new_n313), .B2(new_n597), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT85), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n578), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n577), .A2(KEYINPUT85), .A3(new_n289), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n580), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n613), .B1(G200), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n595), .A2(new_n581), .ZN(new_n620));
  INV_X1    g0420(.A(new_n580), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n615), .B2(new_n616), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(G169), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n620), .B1(new_n623), .B2(KEYINPUT86), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n622), .B2(G169), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n619), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n484), .A2(new_n332), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n490), .A2(new_n629), .A3(new_n483), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n618), .A2(KEYINPUT86), .A3(new_n332), .ZN(new_n632));
  INV_X1    g0432(.A(new_n620), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n626), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n604), .A2(new_n489), .A3(new_n490), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(KEYINPUT26), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n570), .A2(new_n528), .B1(new_n560), .B2(new_n566), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n627), .B(new_n574), .C1(new_n518), .C2(new_n639), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n631), .B(new_n638), .C1(new_n640), .C2(new_n492), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n612), .B1(new_n426), .B2(new_n642), .ZN(G369));
  NAND3_X1  g0443(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  XOR2_X1   g0445(.A(new_n645), .B(KEYINPUT87), .Z(new_n646));
  OAI21_X1  g0446(.A(G213), .B1(new_n644), .B2(KEYINPUT27), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G343), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n507), .ZN(new_n651));
  MUX2_X1   g0451(.A(new_n518), .B(new_n523), .S(new_n651), .Z(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(G330), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n550), .A2(new_n650), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n568), .A2(new_n654), .A3(new_n574), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n568), .B2(new_n649), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n518), .A2(new_n649), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT88), .Z(new_n659));
  AOI22_X1  g0459(.A1(new_n659), .A2(new_n656), .B1(new_n639), .B2(new_n649), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n212), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n215), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n641), .A2(new_n649), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(KEYINPUT29), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT90), .B1(new_n640), .B2(new_n492), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n488), .B1(new_n313), .B2(new_n484), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n463), .A2(G200), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(new_n427), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n630), .B1(new_n674), .B2(new_n464), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n574), .B1(new_n639), .B2(new_n518), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n622), .A2(new_n291), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n634), .A2(new_n635), .B1(new_n613), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT90), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n675), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n637), .A2(KEYINPUT26), .B1(new_n635), .B2(new_n634), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n628), .B1(new_n627), .B2(new_n630), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n671), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n649), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n670), .B1(KEYINPUT29), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n565), .A2(new_n561), .A3(new_n563), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n597), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n438), .B1(new_n456), .B2(new_n289), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n499), .A2(new_n297), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n689), .A2(new_n690), .A3(KEYINPUT30), .A4(new_n691), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(G179), .B1(new_n493), .B2(new_n498), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n618), .A2(new_n572), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n458), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT89), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n463), .A2(new_n572), .A3(new_n618), .A4(new_n697), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT89), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n702), .A3(new_n694), .A4(new_n695), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n700), .A2(new_n650), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n568), .A2(new_n574), .A3(new_n604), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n512), .A2(new_n517), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n521), .A3(new_n515), .A4(new_n509), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n675), .A2(new_n708), .A3(new_n649), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n704), .B1(new_n709), .B2(KEYINPUT31), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n696), .A2(new_n699), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n711), .A2(new_n712), .A3(new_n649), .ZN(new_n713));
  OAI21_X1  g0513(.A(G330), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n687), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n668), .B1(new_n715), .B2(G1), .ZN(G364));
  AND2_X1   g0516(.A1(new_n209), .A2(G13), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n208), .B1(new_n717), .B2(G45), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n663), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n653), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(G330), .B2(new_n652), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n217), .B1(G20), .B2(new_n332), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n297), .A2(new_n291), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n209), .A2(G190), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G179), .A2(G200), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n209), .B1(new_n728), .B2(G190), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n727), .A2(new_n221), .B1(new_n729), .B2(new_n469), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n209), .A2(new_n313), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n725), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n297), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n726), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI22_X1  g0537(.A1(G50), .A2(new_n734), .B1(new_n737), .B2(G77), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n732), .A2(new_n735), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n291), .A2(G179), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n726), .A2(new_n740), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n738), .B1(new_n202), .B2(new_n739), .C1(new_n467), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n732), .A2(new_n740), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n286), .B1(new_n743), .B2(new_n223), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT92), .Z(new_n745));
  NAND2_X1  g0545(.A1(new_n726), .A2(new_n728), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G159), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT32), .ZN(new_n749));
  OR4_X1    g0549(.A1(new_n731), .A2(new_n742), .A3(new_n745), .A4(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n741), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G283), .A2(new_n751), .B1(new_n747), .B2(G329), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT94), .ZN(new_n753));
  INV_X1    g0553(.A(new_n739), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G326), .A2(new_n734), .B1(new_n754), .B2(G322), .ZN(new_n755));
  INV_X1    g0555(.A(new_n743), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G303), .A2(new_n756), .B1(new_n737), .B2(G311), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT33), .B(G317), .Z(new_n758));
  OAI21_X1  g0558(.A(new_n283), .B1(new_n758), .B2(new_n727), .ZN(new_n759));
  INV_X1    g0559(.A(new_n729), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(G294), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n753), .A2(new_n755), .A3(new_n757), .A4(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n724), .B1(new_n750), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n723), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT91), .Z(new_n768));
  NOR2_X1   g0568(.A1(new_n662), .A2(new_n286), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(new_n301), .B2(new_n216), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n245), .B2(new_n301), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n662), .A2(new_n283), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n773), .A2(G355), .B1(new_n500), .B2(new_n662), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n768), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n763), .A2(new_n775), .A3(new_n663), .A4(new_n719), .ZN(new_n776));
  INV_X1    g0576(.A(new_n766), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n652), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n722), .A2(new_n778), .ZN(G396));
  NOR2_X1   g0579(.A1(new_n334), .A2(new_n650), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n329), .A2(new_n650), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n330), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(new_n782), .B2(new_n334), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n641), .A2(new_n649), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT99), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n641), .A2(KEYINPUT99), .A3(new_n649), .A4(new_n783), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n314), .A2(new_n329), .ZN(new_n788));
  INV_X1    g0588(.A(new_n781), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n334), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n780), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n786), .A2(new_n787), .B1(new_n669), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n714), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n720), .B1(new_n794), .B2(new_n714), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n792), .A2(new_n764), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n724), .A2(new_n765), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n720), .B1(G77), .B2(new_n799), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n743), .A2(new_n467), .B1(new_n736), .B2(new_n500), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n283), .B1(new_n729), .B2(new_n469), .C1(new_n553), .C2(new_n739), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n801), .B(new_n802), .C1(G303), .C2(new_n734), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n741), .A2(new_n223), .B1(new_n746), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT96), .Z(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n727), .A2(KEYINPUT95), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n727), .A2(KEYINPUT95), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n803), .B(new_n806), .C1(new_n807), .C2(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G143), .A2(new_n754), .B1(new_n737), .B2(G159), .ZN(new_n812));
  INV_X1    g0612(.A(G137), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n813), .B2(new_n733), .C1(new_n252), .C2(new_n727), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT34), .Z(new_n815));
  OAI21_X1  g0615(.A(new_n286), .B1(new_n743), .B2(new_n201), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n741), .A2(new_n221), .B1(new_n746), .B2(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n816), .B(new_n818), .C1(G58), .C2(new_n760), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT97), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n811), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(KEYINPUT98), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n724), .B1(new_n821), .B2(KEYINPUT98), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n800), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n796), .A2(new_n797), .B1(new_n798), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  AOI21_X1  g0626(.A(new_n780), .B1(new_n786), .B2(new_n787), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n361), .A2(new_n650), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n362), .A2(new_n370), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n369), .A2(new_n368), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n365), .B2(new_n366), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n361), .B(new_n650), .C1(new_n831), .C2(new_n351), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n827), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n648), .B1(new_n413), .B2(new_n414), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n424), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n404), .A2(new_n415), .A3(new_n836), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT37), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n415), .A2(new_n404), .A3(new_n836), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n838), .A2(new_n843), .A3(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n835), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n648), .B1(new_n416), .B2(new_n418), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT39), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n840), .A2(KEYINPUT102), .A3(new_n842), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT102), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n839), .A2(new_n854), .A3(KEYINPUT37), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(new_n838), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n845), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n847), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n852), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n351), .A2(new_n361), .A3(new_n649), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n850), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n849), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n612), .B1(new_n687), .B2(new_n426), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n863), .B(new_n864), .Z(new_n865));
  INV_X1    g0665(.A(KEYINPUT103), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n792), .B1(new_n829), .B2(new_n832), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n700), .A2(new_n650), .A3(new_n703), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(new_n712), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(new_n710), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n839), .A2(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n871), .A2(new_n872), .B1(new_n424), .B2(new_n837), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n873), .B2(new_n853), .ZN(new_n874));
  INV_X1    g0674(.A(new_n847), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT40), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n866), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n492), .A2(new_n605), .A3(new_n650), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n868), .B1(new_n878), .B2(new_n712), .ZN(new_n879));
  INV_X1    g0679(.A(new_n869), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n857), .B2(new_n847), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n881), .A2(new_n883), .A3(KEYINPUT103), .A4(new_n867), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n881), .A2(new_n848), .A3(new_n867), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n877), .A2(new_n884), .B1(new_n885), .B2(new_n882), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n881), .A2(new_n425), .ZN(new_n888));
  OAI21_X1  g0688(.A(G330), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n888), .B2(new_n887), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n865), .A2(new_n890), .B1(new_n208), .B2(new_n717), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n865), .B2(new_n890), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n217), .A2(new_n209), .A3(new_n500), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n472), .B(KEYINPUT100), .Z(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT35), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n896), .B2(new_n895), .ZN(new_n898));
  XOR2_X1   g0698(.A(KEYINPUT101), .B(KEYINPUT36), .Z(new_n899));
  XNOR2_X1  g0699(.A(new_n898), .B(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n216), .B(G77), .C1(new_n202), .C2(new_n221), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n201), .A2(G68), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n208), .B(G13), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  OR3_X1    g0703(.A1(new_n892), .A2(new_n900), .A3(new_n903), .ZN(G367));
  NOR2_X1   g0704(.A1(new_n649), .A2(new_n602), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT104), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n636), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n678), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT105), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n675), .B1(new_n488), .B2(new_n649), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n491), .B2(new_n649), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n656), .A3(new_n659), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT42), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n911), .A2(new_n568), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n650), .B1(new_n915), .B2(new_n491), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n910), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n917), .B(new_n918), .Z(new_n919));
  INV_X1    g0719(.A(new_n657), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n912), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n663), .B(KEYINPUT41), .Z(new_n923));
  NAND2_X1  g0723(.A1(new_n912), .A2(new_n660), .ZN(new_n924));
  XOR2_X1   g0724(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n925));
  XOR2_X1   g0725(.A(new_n924), .B(new_n925), .Z(new_n926));
  NOR2_X1   g0726(.A1(new_n912), .A2(new_n660), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT107), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT44), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(KEYINPUT44), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n920), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n657), .A3(new_n932), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n653), .B(new_n656), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(new_n659), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n934), .A2(new_n715), .A3(new_n935), .A4(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n923), .B1(new_n938), .B2(new_n715), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n922), .B1(new_n939), .B2(new_n719), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n235), .A2(new_n770), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n767), .B1(new_n212), .B2(new_n321), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n720), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n202), .A2(new_n743), .B1(new_n739), .B2(new_n252), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n283), .B(new_n944), .C1(G143), .C2(new_n734), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n760), .A2(G68), .ZN(new_n946));
  INV_X1    g0746(.A(new_n810), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(G159), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n746), .A2(new_n813), .ZN(new_n949));
  INV_X1    g0749(.A(G77), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n741), .A2(new_n950), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n949), .B(new_n951), .C1(G50), .C2(new_n737), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n945), .A2(new_n946), .A3(new_n948), .A4(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT108), .B1(new_n743), .B2(new_n500), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT46), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n553), .B2(new_n810), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G303), .A2(new_n754), .B1(new_n737), .B2(G283), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n734), .A2(G311), .B1(new_n747), .B2(G317), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n760), .A2(G107), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n286), .B1(new_n751), .B2(G97), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n957), .A2(new_n958), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n953), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n943), .B1(new_n964), .B2(new_n723), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n908), .B2(new_n777), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n940), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT110), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n940), .A2(KEYINPUT110), .A3(new_n966), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n970), .A2(new_n972), .ZN(G387));
  AOI22_X1  g0773(.A1(G317), .A2(new_n754), .B1(new_n737), .B2(G303), .ZN(new_n974));
  INV_X1    g0774(.A(G322), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n974), .B1(new_n975), .B2(new_n733), .C1(new_n810), .C2(new_n804), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT48), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(KEYINPUT48), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n756), .A2(G294), .B1(new_n760), .B2(G283), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT49), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n741), .A2(new_n500), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n286), .B(new_n985), .C1(G326), .C2(new_n747), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n743), .A2(new_n950), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n286), .B1(new_n741), .B2(new_n469), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G159), .C2(new_n734), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G68), .A2(new_n737), .B1(new_n747), .B2(G150), .ZN(new_n991));
  INV_X1    g0791(.A(new_n727), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G50), .A2(new_n754), .B1(new_n992), .B2(new_n315), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n729), .A2(new_n321), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n990), .A2(new_n991), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n724), .B1(new_n987), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n656), .A2(new_n777), .ZN(new_n998));
  INV_X1    g0798(.A(new_n773), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n999), .A2(new_n665), .B1(G107), .B2(new_n212), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n240), .A2(new_n301), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT111), .Z(new_n1002));
  INV_X1    g0802(.A(KEYINPUT112), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n665), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n665), .A2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n301), .B1(new_n221), .B2(new_n950), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n256), .A2(G50), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n770), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1000), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n720), .B1(new_n1011), .B2(new_n768), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n997), .A2(new_n998), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n937), .B2(new_n719), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n715), .A2(new_n937), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n663), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n715), .A2(new_n937), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT113), .Z(G393));
  INV_X1    g0819(.A(new_n935), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n657), .B1(new_n931), .B2(new_n932), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1015), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n938), .A3(new_n663), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n934), .A2(new_n719), .A3(new_n935), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n767), .B1(new_n469), .B2(new_n212), .C1(new_n770), .C2(new_n249), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1025), .A2(new_n720), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G317), .A2(new_n734), .B1(new_n754), .B2(G311), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT52), .Z(new_n1028));
  OAI22_X1  g0828(.A1(new_n743), .A2(new_n807), .B1(new_n746), .B2(new_n975), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n283), .B1(new_n729), .B2(new_n500), .C1(new_n467), .C2(new_n741), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(G294), .C2(new_n737), .ZN(new_n1031));
  INV_X1    g0831(.A(G303), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1028), .B(new_n1031), .C1(new_n1032), .C2(new_n810), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G68), .A2(new_n756), .B1(new_n747), .B2(G143), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1034), .B(new_n286), .C1(new_n223), .C2(new_n741), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT114), .Z(new_n1036));
  OAI22_X1  g0836(.A1(new_n733), .A2(new_n252), .B1(new_n739), .B2(new_n377), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT51), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n315), .A2(new_n737), .B1(new_n760), .B2(G77), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n201), .C2(new_n810), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1033), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT115), .Z(new_n1042));
  OAI221_X1 g0842(.A(new_n1026), .B1(new_n724), .B2(new_n1042), .C1(new_n912), .C2(new_n777), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1024), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1023), .A2(new_n1044), .ZN(G390));
  INV_X1    g0845(.A(G330), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n879), .B2(new_n880), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n425), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n612), .B(new_n1048), .C1(new_n687), .C2(new_n426), .ZN(new_n1049));
  OAI211_X1 g0849(.A(G330), .B(new_n783), .C1(new_n710), .C2(new_n713), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n833), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n881), .A2(G330), .A3(new_n783), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n834), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n685), .A2(new_n649), .A3(new_n790), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(KEYINPUT116), .A3(new_n791), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT116), .B1(new_n1055), .B2(new_n791), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1052), .B(new_n1054), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n881), .A2(G330), .A3(new_n867), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1051), .B2(new_n833), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n827), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1049), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT117), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1055), .A2(new_n791), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT116), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1069), .A2(new_n833), .A3(new_n1056), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n861), .B1(new_n857), .B2(new_n847), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n860), .B1(new_n827), .B2(new_n834), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n859), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1075), .A3(new_n1052), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1070), .A2(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n1060), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1066), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1076), .ZN(new_n1081));
  OAI211_X1 g0881(.A(KEYINPUT117), .B(new_n1065), .C1(new_n1081), .C2(new_n1078), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1082), .A3(new_n663), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1081), .A2(new_n1078), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1074), .A2(new_n764), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n720), .B1(new_n315), .B2(new_n799), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n741), .A2(new_n221), .B1(new_n746), .B2(new_n553), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n286), .B(new_n1087), .C1(G87), .C2(new_n756), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n947), .A2(G107), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n760), .A2(G77), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n733), .A2(new_n807), .B1(new_n736), .B2(new_n469), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G116), .B2(new_n754), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(G125), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n286), .B1(new_n729), .B2(new_n377), .C1(new_n1094), .C2(new_n746), .ZN(new_n1095));
  INV_X1    g0895(.A(G128), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n733), .A2(new_n1096), .B1(new_n739), .B2(new_n817), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n201), .A2(new_n741), .B1(new_n736), .B2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n1095), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n743), .A2(new_n252), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(new_n813), .C2(new_n810), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1093), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1086), .B1(new_n1104), .B2(new_n723), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1084), .A2(new_n719), .B1(new_n1085), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1083), .A2(new_n1106), .ZN(G378));
  OAI211_X1 g0907(.A(new_n1076), .B(new_n1064), .C1(new_n1077), .C2(new_n1060), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1049), .B(KEYINPUT121), .Z(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n886), .A2(G330), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n295), .A2(new_n299), .ZN(new_n1112));
  XOR2_X1   g0912(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT120), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1112), .B(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n264), .A2(new_n648), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT119), .Z(new_n1117));
  XNOR2_X1  g0917(.A(new_n1115), .B(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1111), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n863), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n886), .A2(G330), .A3(new_n1118), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n877), .A2(new_n884), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n885), .A2(new_n882), .ZN(new_n1125));
  AND4_X1   g0925(.A1(G330), .A2(new_n1124), .A3(new_n1125), .A4(new_n1118), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1118), .B1(new_n886), .B2(G330), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n863), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1110), .A2(KEYINPUT57), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT122), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1110), .A2(new_n1129), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT57), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT122), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1110), .A2(new_n1135), .A3(new_n1129), .A4(KEYINPUT57), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1131), .A2(new_n1134), .A3(new_n663), .A4(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n718), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1119), .A2(new_n764), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n720), .B1(G50), .B2(new_n799), .ZN(new_n1140));
  AOI21_X1  g0940(.A(G50), .B1(new_n279), .B2(new_n300), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n741), .A2(new_n202), .B1(new_n746), .B2(new_n807), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n1142), .A2(new_n988), .A3(G41), .A4(new_n286), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n734), .A2(G116), .B1(new_n737), .B2(new_n317), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G97), .A2(new_n992), .B1(new_n754), .B2(G107), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1143), .A2(new_n946), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT58), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1141), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(G33), .B(G41), .C1(new_n747), .C2(G124), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n727), .A2(new_n817), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n733), .A2(new_n1094), .B1(new_n736), .B2(new_n813), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G150), .C2(new_n760), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1096), .A2(new_n739), .B1(new_n743), .B2(new_n1098), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1149), .B1(new_n377), .B2(new_n741), .C1(new_n1155), .C2(KEYINPUT59), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1148), .B1(new_n1147), .B2(new_n1146), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1140), .B1(new_n1158), .B2(new_n723), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1139), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1138), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1137), .A2(new_n1162), .ZN(G375));
  NAND2_X1  g0963(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n1049), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n923), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n1065), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n833), .A2(new_n765), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT123), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n720), .B1(G68), .B2(new_n799), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n739), .A2(new_n807), .B1(new_n746), .B2(new_n1032), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n1172), .A2(new_n951), .A3(new_n994), .A4(new_n286), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n733), .A2(new_n553), .B1(new_n743), .B2(new_n469), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G107), .B2(new_n737), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(new_n500), .C2(new_n810), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G137), .A2(new_n754), .B1(new_n747), .B2(G128), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n283), .B1(new_n751), .B2(G58), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n201), .C2(new_n729), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G159), .A2(new_n756), .B1(new_n737), .B2(G150), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n817), .B2(new_n733), .C1(new_n810), .C2(new_n1098), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1176), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1171), .B1(new_n1182), .B2(new_n723), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1164), .A2(new_n719), .B1(new_n1170), .B2(new_n1183), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1168), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(G381));
  NOR2_X1   g0986(.A1(G375), .A2(G378), .ZN(new_n1187));
  OR2_X1    g0987(.A1(G393), .A2(G396), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1188), .A2(G384), .A3(G390), .A4(G381), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(new_n970), .C2(new_n972), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT124), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(G407));
  INV_X1    g0992(.A(G343), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1187), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(G407), .A2(G213), .A3(new_n1194), .ZN(G409));
  INV_X1    g0995(.A(KEYINPUT62), .ZN(new_n1196));
  INV_X1    g0996(.A(G378), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1137), .B2(new_n1162), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1193), .A2(G213), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1108), .A2(new_n1109), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1167), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1083), .A3(new_n1106), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1129), .A2(new_n719), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(KEYINPUT125), .A3(new_n1160), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT125), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1138), .B2(new_n1161), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1199), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT60), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1166), .B1(new_n1209), .B2(new_n1064), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1165), .A2(KEYINPUT60), .A3(new_n1049), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n663), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1184), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n825), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(G384), .A3(new_n1184), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1198), .A2(new_n1208), .A3(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1196), .B1(new_n1217), .B2(KEYINPUT127), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1201), .A2(new_n1083), .A3(new_n1106), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1219), .A2(new_n1220), .B1(G213), .B2(new_n1193), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1216), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1162), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n663), .B1(new_n1200), .B2(KEYINPUT57), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1135), .B1(new_n1200), .B2(KEYINPUT57), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1223), .B1(new_n1226), .B2(new_n1136), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1221), .B(new_n1222), .C1(new_n1227), .C2(new_n1197), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT127), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(KEYINPUT62), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1221), .B1(new_n1227), .B2(new_n1197), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1193), .A2(G213), .A3(G2897), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1214), .A2(new_n1215), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1232), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT61), .B1(new_n1231), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1218), .A2(new_n1230), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n940), .A2(new_n966), .A3(G390), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(G393), .B(G396), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n969), .A2(new_n971), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(G390), .B(KEYINPUT126), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n967), .A2(new_n1023), .A3(new_n1044), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1238), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1239), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1237), .A2(new_n1248), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1217), .A2(KEYINPUT63), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1217), .A2(KEYINPUT63), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1236), .A4(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1249), .A2(new_n1253), .ZN(G405));
  OR2_X1    g1054(.A1(new_n1187), .A2(new_n1198), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1222), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1187), .A2(new_n1198), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1216), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1248), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1258), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1257), .A2(new_n1216), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1251), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(G402));
endmodule


