//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  NAND2_X1  g000(.A1(KEYINPUT0), .A2(G128), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(KEYINPUT64), .A3(G143), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(G146), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n188), .B(new_n190), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  OR2_X1    g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n189), .A2(G143), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n187), .B(new_n196), .C1(new_n194), .C2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n190), .B(new_n202), .C1(new_n193), .C2(new_n194), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(G143), .B2(new_n189), .ZN(new_n205));
  OAI22_X1  g019(.A1(new_n205), .A2(new_n201), .B1(new_n194), .B2(new_n197), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G953), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G224), .ZN(new_n211));
  XOR2_X1   g025(.A(new_n209), .B(new_n211), .Z(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G116), .ZN(new_n214));
  INV_X1    g028(.A(G116), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G119), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT2), .B(G113), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT66), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G113), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT2), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT2), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G113), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G116), .B(G119), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(KEYINPUT5), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n229), .B(G113), .C1(KEYINPUT5), .C2(new_n214), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT82), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G107), .ZN(new_n234));
  INV_X1    g048(.A(G107), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT82), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n232), .B(G104), .C1(new_n234), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G101), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT83), .B1(new_n235), .B2(G104), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n240));
  INV_X1    g054(.A(G104), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(G107), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n235), .A2(G104), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n237), .A2(new_n238), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n235), .A2(KEYINPUT82), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n233), .A2(G107), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n244), .B1(new_n249), .B2(G104), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G101), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n231), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  XOR2_X1   g068(.A(G110), .B(G122), .Z(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n237), .A2(new_n243), .A3(new_n245), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G101), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n246), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT84), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT84), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n258), .A2(new_n261), .A3(KEYINPUT4), .A4(new_n246), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT85), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n264), .A2(KEYINPUT4), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(KEYINPUT4), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n257), .A2(G101), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n217), .A2(new_n218), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT66), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n226), .B1(new_n224), .B2(new_n225), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n254), .B(new_n256), .C1(new_n263), .C2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n255), .B(KEYINPUT89), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n260), .B2(new_n262), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(new_n253), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(KEYINPUT6), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n275), .C1(new_n276), .C2(new_n253), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n280), .A2(KEYINPUT90), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(KEYINPUT90), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n212), .B(new_n278), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n231), .B(new_n252), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n255), .B(KEYINPUT8), .Z(new_n285));
  INV_X1    g099(.A(KEYINPUT91), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT7), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n286), .A2(new_n287), .B1(new_n210), .B2(G224), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n209), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT92), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n209), .A2(KEYINPUT92), .A3(new_n289), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n284), .A2(new_n285), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n200), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n208), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(KEYINPUT93), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n274), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n298), .A2(KEYINPUT94), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT94), .B1(new_n298), .B2(new_n299), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n283), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n283), .B(new_n303), .C1(new_n300), .C2(new_n301), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(KEYINPUT95), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT94), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n276), .A2(new_n253), .A3(new_n255), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n284), .A2(new_n285), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n292), .A2(new_n293), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n309), .A2(new_n312), .A3(new_n296), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n308), .B1(new_n313), .B2(G902), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n298), .A2(KEYINPUT94), .A3(new_n299), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n303), .B1(new_n316), .B2(new_n283), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT95), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n210), .A2(G952), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(G234), .B2(G237), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT21), .B(G898), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(G234), .A2(G237), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(G902), .A3(G953), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n321), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(G214), .B1(G237), .B2(G902), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n307), .A2(new_n319), .A3(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT9), .B(G234), .Z(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G221), .B1(new_n333), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G469), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n260), .A2(new_n262), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n195), .A2(new_n198), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n268), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT11), .ZN(new_n340));
  INV_X1    g154(.A(G134), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(G137), .ZN(new_n342));
  INV_X1    g156(.A(G137), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT11), .A3(G134), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(G137), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G131), .ZN(new_n347));
  INV_X1    g161(.A(G131), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n342), .A2(new_n344), .A3(new_n348), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n252), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n203), .A2(new_n206), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n189), .A2(KEYINPUT64), .A3(G143), .ZN(new_n357));
  INV_X1    g171(.A(new_n194), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT64), .B1(new_n189), .B2(G143), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n205), .A2(new_n201), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n203), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n362), .A2(new_n251), .A3(new_n246), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n356), .B1(KEYINPUT10), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n339), .A2(new_n351), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n210), .A2(G227), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT81), .ZN(new_n368));
  XNOR2_X1  g182(.A(G110), .B(G140), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n252), .A2(new_n353), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n251), .A3(new_n246), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n351), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(KEYINPUT12), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT12), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n376), .B(new_n351), .C1(new_n372), .C2(new_n373), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT87), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n203), .A2(new_n206), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n246), .B2(new_n251), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n350), .B1(new_n363), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n376), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n374), .A2(KEYINPUT12), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n366), .A2(new_n371), .A3(new_n378), .A4(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT88), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n375), .A2(new_n377), .A3(KEYINPUT87), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n384), .B1(new_n382), .B2(new_n383), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n268), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n260), .B2(new_n262), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n364), .B1(new_n393), .B2(new_n338), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n370), .B1(new_n394), .B2(new_n351), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n395), .A3(KEYINPUT88), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  AOI211_X1 g211(.A(new_n199), .B(new_n392), .C1(new_n260), .C2(new_n262), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT86), .B1(new_n398), .B2(new_n364), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n339), .A2(new_n400), .A3(new_n365), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n350), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n371), .B1(new_n402), .B2(new_n366), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n336), .B(new_n299), .C1(new_n397), .C2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n336), .A2(new_n299), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n366), .B1(new_n377), .B2(new_n375), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n402), .A2(new_n395), .B1(new_n406), .B2(new_n370), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n405), .B1(new_n407), .B2(G469), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n335), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G125), .B(G140), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n411));
  INV_X1    g225(.A(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G125), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n413), .A2(KEYINPUT16), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n189), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(G146), .A3(new_n414), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G237), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n210), .A3(G214), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n192), .ZN(new_n421));
  NOR2_X1   g235(.A1(G237), .A2(G953), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(G143), .A3(G214), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT17), .A3(G131), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(G131), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n418), .B(new_n425), .C1(KEYINPUT17), .C2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G113), .B(G122), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(new_n241), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT96), .ZN(new_n430));
  INV_X1    g244(.A(new_n423), .ZN(new_n431));
  AOI21_X1  g245(.A(G143), .B1(new_n422), .B2(G214), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(KEYINPUT18), .A2(G131), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n421), .A2(KEYINPUT96), .A3(new_n423), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT97), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n410), .A2(KEYINPUT75), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n207), .A2(G140), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n413), .A2(new_n441), .A3(KEYINPUT75), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n189), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n410), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G146), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n431), .A2(new_n432), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n443), .A2(new_n445), .B1(new_n446), .B2(new_n434), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n433), .A2(KEYINPUT97), .A3(new_n435), .A4(new_n436), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n439), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n427), .A2(new_n429), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n429), .B1(new_n427), .B2(new_n449), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n299), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G475), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n444), .A2(KEYINPUT19), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n440), .A2(new_n442), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(KEYINPUT19), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n426), .B(new_n417), .C1(new_n458), .C2(G146), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n449), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n429), .B1(new_n460), .B2(KEYINPUT98), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT98), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n449), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n450), .ZN(new_n465));
  NOR2_X1   g279(.A1(G475), .A2(G902), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n455), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n451), .B1(new_n463), .B2(new_n461), .ZN(new_n468));
  INV_X1    g282(.A(new_n466), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n468), .A2(KEYINPUT20), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n454), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G217), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n333), .A2(new_n472), .A3(G953), .ZN(new_n473));
  XNOR2_X1  g287(.A(G128), .B(G143), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n341), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n475), .B(KEYINPUT99), .Z(new_n476));
  XNOR2_X1  g290(.A(G116), .B(G122), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n249), .B(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n341), .B1(new_n474), .B2(KEYINPUT13), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n192), .A2(G128), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(KEYINPUT13), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n476), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n474), .B(new_n341), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n215), .A2(KEYINPUT14), .A3(G122), .ZN(new_n484));
  INV_X1    g298(.A(new_n477), .ZN(new_n485));
  OAI211_X1 g299(.A(G107), .B(new_n484), .C1(new_n485), .C2(KEYINPUT14), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n249), .A2(new_n477), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n473), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n482), .A2(new_n488), .A3(new_n473), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G478), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n471), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n409), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n331), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT70), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n272), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n228), .A2(KEYINPUT67), .A3(new_n269), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n341), .A2(G137), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n343), .A2(G134), .ZN(new_n506));
  OAI21_X1  g320(.A(G131), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n349), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n338), .A2(new_n350), .B1(new_n508), .B2(new_n379), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT28), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n349), .A2(new_n507), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT65), .B1(new_n353), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n338), .A2(new_n350), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT65), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n379), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n272), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT69), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n228), .A2(KEYINPUT67), .A3(new_n269), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT67), .B1(new_n228), .B2(new_n269), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n509), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT69), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n516), .A2(new_n522), .A3(new_n272), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n518), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n510), .B1(new_n524), .B2(KEYINPUT28), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n422), .A2(G210), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(G101), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n529), .B(KEYINPUT68), .Z(new_n530));
  OAI21_X1  g344(.A(new_n500), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n516), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n508), .A2(new_n379), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n513), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n533), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n272), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n529), .B(new_n521), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT31), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n535), .A2(new_n532), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n532), .B2(new_n516), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n272), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n543), .A2(KEYINPUT31), .A3(new_n529), .A4(new_n521), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n530), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n547));
  INV_X1    g361(.A(new_n521), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(KEYINPUT69), .B2(new_n517), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n549), .B2(new_n523), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT70), .B(new_n546), .C1(new_n550), .C2(new_n510), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n531), .A2(new_n545), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(G472), .A2(G902), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT32), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n199), .B1(new_n347), .B2(new_n349), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n511), .B1(new_n206), .B2(new_n203), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n502), .B(new_n503), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n521), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT28), .ZN(new_n561));
  INV_X1    g375(.A(new_n510), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n561), .A2(KEYINPUT29), .A3(new_n529), .A4(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT71), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n510), .B1(new_n560), .B2(KEYINPUT28), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n566), .A2(KEYINPUT71), .A3(KEYINPUT29), .A4(new_n529), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n299), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT72), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT72), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n565), .A2(new_n570), .A3(new_n299), .A4(new_n567), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n534), .A2(KEYINPUT65), .B1(new_n338), .B2(new_n350), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n537), .B1(new_n572), .B2(new_n515), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n521), .B1(new_n573), .B2(new_n522), .ZN(new_n574));
  INV_X1    g388(.A(new_n523), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT28), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n562), .A3(new_n530), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT29), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n536), .A2(new_n537), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n548), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n577), .B(new_n578), .C1(new_n529), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n569), .A2(new_n571), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G472), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n552), .A2(KEYINPUT32), .A3(new_n553), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n556), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n201), .A2(G119), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT23), .ZN(new_n588));
  INV_X1    g402(.A(G110), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT23), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n213), .B2(G128), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n588), .B(new_n589), .C1(new_n587), .C2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT73), .B1(new_n213), .B2(G128), .ZN(new_n593));
  MUX2_X1   g407(.A(KEYINPUT73), .B(new_n593), .S(new_n586), .Z(new_n594));
  XOR2_X1   g408(.A(KEYINPUT24), .B(G110), .Z(new_n595));
  OAI21_X1  g409(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT74), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n592), .B(KEYINPUT74), .C1(new_n594), .C2(new_n595), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n598), .A2(new_n417), .A3(new_n599), .A4(new_n443), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n588), .B1(new_n587), .B2(new_n591), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n594), .A2(new_n595), .B1(new_n601), .B2(G110), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n416), .A2(new_n417), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT22), .B(G137), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n210), .A2(G221), .A3(G234), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n600), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(KEYINPUT76), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n600), .B2(new_n604), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT77), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n600), .A2(KEYINPUT77), .A3(new_n604), .A4(new_n607), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n299), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT25), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n612), .A2(KEYINPUT25), .A3(new_n299), .A4(new_n613), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n472), .B1(G234), .B2(new_n299), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT80), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n619), .A2(G902), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(KEYINPUT78), .Z(new_n623));
  NAND3_X1  g437(.A1(new_n612), .A2(new_n613), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT79), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n620), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n624), .B(KEYINPUT79), .ZN(new_n628));
  INV_X1    g442(.A(new_n619), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n616), .B2(new_n617), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT80), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n585), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n499), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  INV_X1    g450(.A(new_n327), .ZN(new_n637));
  INV_X1    g451(.A(new_n306), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n328), .B(new_n637), .C1(new_n638), .C2(new_n317), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n465), .A2(new_n455), .A3(new_n466), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT20), .B1(new_n468), .B2(new_n469), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n640), .A2(new_n641), .B1(G475), .B2(new_n453), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT101), .B1(new_n492), .B2(G478), .ZN(new_n643));
  INV_X1    g457(.A(new_n491), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n299), .B1(new_n644), .B2(new_n489), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n493), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT100), .B1(new_n482), .B2(new_n488), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n491), .A3(new_n490), .ZN(new_n652));
  OAI22_X1  g466(.A1(new_n644), .A2(new_n489), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n652), .A2(G478), .A3(new_n653), .A4(new_n299), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n642), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT102), .B1(new_n639), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n329), .B1(new_n305), .B2(new_n306), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n637), .A4(new_n656), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n552), .A2(new_n299), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n663), .A2(G472), .B1(new_n553), .B2(new_n552), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n409), .A2(new_n664), .A3(new_n632), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NAND2_X1  g482(.A1(new_n642), .A2(new_n496), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n639), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  AND3_X1   g487(.A1(new_n307), .A2(new_n319), .A3(new_n330), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n409), .A2(new_n497), .ZN(new_n675));
  INV_X1    g489(.A(new_n623), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT36), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n609), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT103), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n600), .A2(new_n604), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n676), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n618), .B2(new_n619), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n674), .A2(new_n675), .A3(new_n664), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  AOI211_X1 g502(.A(new_n329), .B(new_n684), .C1(new_n305), .C2(new_n306), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n321), .B1(new_n326), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n669), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n689), .A2(new_n585), .A3(new_n409), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  XNOR2_X1  g508(.A(new_n691), .B(KEYINPUT39), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n409), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT40), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n307), .A2(new_n319), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(KEYINPUT38), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT38), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n307), .B2(new_n319), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n580), .A2(new_n529), .B1(new_n560), .B2(new_n546), .ZN(new_n705));
  OAI21_X1  g519(.A(G472), .B1(new_n705), .B2(G902), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n556), .A2(new_n584), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT104), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n642), .A2(new_n495), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n328), .A3(new_n684), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n710), .B(KEYINPUT105), .Z(new_n711));
  NAND4_X1  g525(.A1(new_n699), .A2(new_n704), .A3(new_n708), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND2_X1  g527(.A1(new_n305), .A2(new_n306), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n642), .A2(new_n655), .A3(new_n691), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n714), .A2(new_n328), .A3(new_n685), .A4(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(KEYINPUT106), .A3(new_n585), .A4(new_n409), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n585), .A2(new_n409), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n659), .A2(new_n685), .A3(new_n715), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT107), .B(G146), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G48));
  OAI21_X1  g538(.A(new_n299), .B1(new_n397), .B2(new_n403), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n336), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  OAI221_X1 g542(.A(new_n299), .B1(new_n726), .B2(new_n336), .C1(new_n397), .C2(new_n403), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n334), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n633), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n662), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n670), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  AND3_X1   g550(.A1(new_n556), .A2(new_n583), .A3(new_n584), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n728), .A2(new_n729), .A3(new_n637), .A4(new_n334), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n659), .A2(new_n497), .A3(new_n685), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  AND2_X1   g556(.A1(new_n659), .A2(new_n709), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n728), .A2(new_n334), .A3(new_n729), .ZN(new_n744));
  INV_X1    g558(.A(G472), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n552), .B2(new_n299), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n566), .A2(new_n530), .ZN(new_n747));
  AOI211_X1 g561(.A(G472), .B(G902), .C1(new_n545), .C2(new_n747), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n746), .A2(new_n748), .A3(new_n630), .A4(new_n628), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n743), .A2(new_n637), .A3(new_n744), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NOR3_X1   g565(.A1(new_n746), .A2(new_n684), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n648), .A2(new_n654), .ZN(new_n753));
  INV_X1    g567(.A(new_n691), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n471), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT109), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n471), .A2(new_n757), .A3(new_n753), .A4(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n744), .A2(new_n659), .A3(new_n752), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  AOI21_X1  g575(.A(new_n329), .B1(new_n307), .B2(new_n319), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n762), .A2(new_n409), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n628), .A2(new_n630), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n585), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n764), .B1(new_n585), .B2(new_n765), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n763), .B(new_n759), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT42), .ZN(new_n769));
  INV_X1    g583(.A(new_n762), .ZN(new_n770));
  INV_X1    g584(.A(new_n409), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n770), .A2(new_n633), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n759), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n348), .ZN(G33));
  NAND2_X1  g590(.A1(new_n772), .A2(new_n692), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n642), .A2(KEYINPUT111), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n640), .A2(new_n641), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n753), .A2(new_n782), .A3(new_n454), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n642), .B(new_n753), .C1(KEYINPUT111), .C2(KEYINPUT43), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n664), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n784), .A2(KEYINPUT112), .A3(new_n785), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n685), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n779), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n407), .A2(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n407), .A2(KEYINPUT45), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(G469), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n405), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n404), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT46), .B1(new_n796), .B2(new_n797), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n334), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n695), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n770), .B1(new_n791), .B2(new_n792), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n790), .A2(new_n685), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n664), .B1(new_n786), .B2(new_n787), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(KEYINPUT113), .A3(new_n805), .A4(KEYINPUT44), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n793), .A2(new_n802), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G137), .ZN(G39));
  OR2_X1    g622(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n770), .A2(new_n632), .A3(new_n755), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n809), .A2(new_n737), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n809), .A2(new_n810), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n728), .A2(new_n729), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n334), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n321), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(new_n784), .B2(new_n785), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n749), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n770), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n814), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n704), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n730), .A2(new_n328), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n820), .B1(new_n824), .B2(KEYINPUT118), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n824), .A2(KEYINPUT118), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n823), .A2(new_n825), .A3(KEYINPUT50), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n828));
  INV_X1    g642(.A(new_n820), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n824), .A2(KEYINPUT118), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n701), .A2(new_n703), .B1(new_n824), .B2(KEYINPUT118), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n762), .A2(new_n744), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n632), .A2(new_n321), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n708), .A2(new_n834), .A3(new_n471), .A4(new_n835), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n827), .A2(new_n833), .B1(new_n836), .B2(new_n655), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n762), .A2(new_n744), .A3(new_n819), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n752), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n838), .B1(new_n837), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n822), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(KEYINPUT120), .B(new_n822), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OR4_X1    g661(.A1(new_n657), .A2(new_n708), .A3(new_n834), .A4(new_n835), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n766), .A2(new_n767), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n839), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT121), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT48), .ZN(new_n852));
  INV_X1    g666(.A(new_n816), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(KEYINPUT117), .A3(new_n335), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n815), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT117), .B1(new_n853), .B2(new_n335), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n821), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n840), .A3(new_n837), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n320), .B1(new_n858), .B2(new_n814), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n847), .A2(new_n848), .A3(new_n852), .A4(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n760), .A2(new_n693), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n771), .A2(new_n691), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n743), .A3(new_n684), .A4(new_n707), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n722), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT116), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n722), .A2(new_n861), .A3(new_n867), .A4(new_n863), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n669), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n665), .A2(new_n674), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n686), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n686), .B2(new_n871), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n731), .B1(new_n662), .B2(new_n670), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n634), .A2(new_n499), .B1(new_n739), .B2(new_n740), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n665), .A2(new_n674), .A3(new_n656), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n750), .A4(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n782), .A2(new_n495), .A3(new_n454), .A4(new_n754), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT115), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n881), .A2(KEYINPUT115), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n585), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n746), .A2(new_n748), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n759), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n684), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n772), .A2(new_n692), .B1(new_n887), .B2(new_n763), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n769), .A2(new_n774), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n864), .A2(KEYINPUT52), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n869), .A2(new_n880), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n865), .A2(new_n868), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT52), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n635), .A2(new_n741), .A3(new_n878), .A4(new_n750), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n896), .B(new_n876), .C1(new_n874), .C2(new_n873), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n769), .A2(new_n888), .A3(new_n774), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n895), .A2(new_n899), .A3(KEYINPUT53), .A4(new_n869), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n829), .A2(new_n659), .A3(new_n744), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n869), .A2(new_n889), .A3(new_n880), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n866), .B1(new_n865), .B2(new_n868), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n892), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n899), .A2(KEYINPUT53), .A3(new_n869), .A4(new_n890), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n902), .A2(new_n903), .A3(new_n909), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n860), .A2(new_n910), .B1(G952), .B2(G953), .ZN(new_n911));
  OR3_X1    g725(.A1(new_n704), .A2(new_n335), .A3(new_n783), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n816), .A2(KEYINPUT49), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n816), .A2(KEYINPUT49), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n765), .A3(new_n914), .ZN(new_n915));
  OR4_X1    g729(.A1(new_n329), .A2(new_n912), .A3(new_n708), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n916), .ZN(G75));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n906), .A2(new_n908), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(G902), .ZN(new_n920));
  INV_X1    g734(.A(G210), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n212), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT55), .Z(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n210), .A2(G952), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n925), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n918), .B(new_n929), .C1(new_n920), .C2(new_n921), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n926), .A2(new_n928), .A3(new_n930), .ZN(G51));
  NAND2_X1  g745(.A1(new_n797), .A2(KEYINPUT57), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n797), .A2(KEYINPUT57), .ZN(new_n933));
  INV_X1    g747(.A(new_n909), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n932), .B(new_n933), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n397), .A2(new_n403), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n299), .B1(new_n906), .B2(new_n908), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  INV_X1    g754(.A(new_n796), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n939), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n927), .B1(new_n938), .B2(new_n944), .ZN(G54));
  AND2_X1   g759(.A1(KEYINPUT58), .A2(G475), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n919), .A2(G902), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n468), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n939), .A2(new_n465), .A3(new_n946), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n928), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n948), .A2(new_n952), .A3(new_n928), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(G60));
  NAND2_X1  g768(.A1(G478), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT59), .Z(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n902), .B2(new_n909), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n652), .A2(new_n653), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT124), .Z(new_n959));
  OAI21_X1  g773(.A(new_n928), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n934), .A2(new_n935), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n961), .A2(new_n956), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n960), .B1(new_n959), .B2(new_n962), .ZN(G63));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT60), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n919), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n612), .A2(new_n613), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n681), .A2(new_n682), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n919), .A2(new_n969), .A3(new_n965), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n928), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n968), .A2(KEYINPUT61), .A3(new_n928), .A4(new_n970), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(G66));
  NAND2_X1  g789(.A1(new_n897), .A2(new_n210), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n322), .A2(G224), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n976), .B(KEYINPUT125), .C1(new_n210), .C2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(KEYINPUT125), .B2(new_n976), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n923), .B1(G898), .B2(new_n210), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n979), .B(new_n980), .Z(G69));
  XNOR2_X1  g795(.A(new_n542), .B(new_n458), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n777), .A2(new_n722), .A3(new_n861), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n793), .A2(new_n803), .A3(new_n806), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n849), .A2(new_n743), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n983), .B1(new_n986), .B2(new_n802), .ZN(new_n987));
  INV_X1    g801(.A(new_n775), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n987), .A2(new_n988), .A3(new_n812), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n982), .B1(new_n989), .B2(new_n210), .ZN(new_n990));
  OAI21_X1  g804(.A(G953), .B1(new_n690), .B2(G227), .ZN(new_n991));
  NAND3_X1  g805(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n712), .A2(new_n722), .A3(new_n861), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n712), .A2(new_n995), .A3(new_n722), .A4(new_n861), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n994), .A2(new_n812), .A3(new_n996), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n772), .B(new_n696), .C1(new_n656), .C2(new_n870), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n807), .A2(new_n210), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n992), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  AOI22_X1  g814(.A1(new_n990), .A2(new_n991), .B1(new_n1000), .B2(new_n982), .ZN(G72));
  NAND4_X1  g815(.A1(new_n987), .A2(new_n988), .A3(new_n812), .A4(new_n880), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT63), .Z(new_n1004));
  NAND2_X1  g818(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n579), .A2(new_n529), .A3(new_n548), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n880), .A2(new_n807), .A3(new_n998), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1004), .B1(new_n1008), .B2(new_n997), .ZN(new_n1009));
  INV_X1    g823(.A(new_n529), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n580), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n927), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1011), .A2(new_n1006), .ZN(new_n1015));
  AND4_X1   g829(.A1(new_n1014), .A2(new_n901), .A3(new_n1004), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1004), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(new_n893), .B2(new_n900), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1014), .B1(new_n1018), .B2(new_n1015), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1013), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n1013), .B(KEYINPUT127), .C1(new_n1016), .C2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1022), .A2(new_n1023), .ZN(G57));
endmodule


