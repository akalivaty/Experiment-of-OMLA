

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591;

  XNOR2_X1 U322 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n415) );
  XNOR2_X1 U323 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U324 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U325 ( .A(n381), .B(n380), .ZN(n479) );
  XNOR2_X1 U326 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U327 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U328 ( .A(G85GAT), .B(KEYINPUT72), .Z(n360) );
  XOR2_X1 U329 ( .A(G71GAT), .B(G120GAT), .Z(n291) );
  XNOR2_X1 U330 ( .A(G99GAT), .B(G176GAT), .ZN(n290) );
  XNOR2_X1 U331 ( .A(n291), .B(n290), .ZN(n440) );
  XNOR2_X1 U332 ( .A(n440), .B(KEYINPUT71), .ZN(n292) );
  XNOR2_X1 U333 ( .A(n292), .B(KEYINPUT32), .ZN(n295) );
  XOR2_X1 U334 ( .A(G57GAT), .B(KEYINPUT13), .Z(n343) );
  XNOR2_X1 U335 ( .A(n343), .B(KEYINPUT33), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n293), .B(KEYINPUT31), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n299) );
  XNOR2_X1 U338 ( .A(G106GAT), .B(G78GAT), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n296), .B(G148GAT), .ZN(n430) );
  XNOR2_X1 U340 ( .A(G204GAT), .B(G92GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n297), .B(G64GAT), .ZN(n327) );
  XNOR2_X1 U342 ( .A(n430), .B(n327), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n360), .B(n300), .ZN(n302) );
  NAND2_X1 U345 ( .A1(G230GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n302), .B(n301), .ZN(n340) );
  XNOR2_X1 U347 ( .A(KEYINPUT41), .B(n340), .ZN(n560) );
  XOR2_X1 U348 ( .A(KEYINPUT104), .B(n560), .Z(n542) );
  XOR2_X1 U349 ( .A(G162GAT), .B(G134GAT), .Z(n304) );
  XNOR2_X1 U350 ( .A(G113GAT), .B(G120GAT), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U352 ( .A(KEYINPUT91), .B(KEYINPUT4), .Z(n306) );
  XNOR2_X1 U353 ( .A(G141GAT), .B(G148GAT), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U355 ( .A(n308), .B(n307), .Z(n313) );
  XOR2_X1 U356 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n310) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U359 ( .A(KEYINPUT89), .B(n311), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n322) );
  XOR2_X1 U361 ( .A(G57GAT), .B(KEYINPUT90), .Z(n315) );
  XNOR2_X1 U362 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n320) );
  XNOR2_X1 U364 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n316), .B(KEYINPUT2), .ZN(n429) );
  XOR2_X1 U366 ( .A(G85GAT), .B(n429), .Z(n318) );
  XOR2_X1 U367 ( .A(KEYINPUT0), .B(G127GAT), .Z(n448) );
  XNOR2_X1 U368 ( .A(G29GAT), .B(n448), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U370 ( .A(n320), .B(n319), .Z(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n524) );
  XOR2_X1 U372 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n324) );
  XNOR2_X1 U373 ( .A(KEYINPUT93), .B(KEYINPUT95), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n335) );
  XOR2_X1 U375 ( .A(G190GAT), .B(G176GAT), .Z(n326) );
  NAND2_X1 U376 ( .A1(G226GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n328) );
  XOR2_X1 U378 ( .A(n328), .B(n327), .Z(n333) );
  XNOR2_X1 U379 ( .A(G36GAT), .B(G197GAT), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n329), .B(G8GAT), .ZN(n388) );
  XOR2_X1 U381 ( .A(G211GAT), .B(KEYINPUT21), .Z(n331) );
  XNOR2_X1 U382 ( .A(G218GAT), .B(KEYINPUT87), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n420) );
  XNOR2_X1 U384 ( .A(n388), .B(n420), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U387 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n337) );
  XNOR2_X1 U388 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(n338), .ZN(n452) );
  XNOR2_X1 U391 ( .A(n339), .B(n452), .ZN(n527) );
  BUF_X1 U392 ( .A(n340), .Z(n580) );
  XOR2_X1 U393 ( .A(G78GAT), .B(G127GAT), .Z(n342) );
  XNOR2_X1 U394 ( .A(G22GAT), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U396 ( .A(n344), .B(n343), .Z(n346) );
  XNOR2_X1 U397 ( .A(G15GAT), .B(G71GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n359) );
  XOR2_X1 U399 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n348) );
  NAND2_X1 U400 ( .A1(G231GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U402 ( .A(n349), .B(KEYINPUT75), .Z(n357) );
  XOR2_X1 U403 ( .A(G64GAT), .B(G211GAT), .Z(n351) );
  XNOR2_X1 U404 ( .A(G1GAT), .B(G155GAT), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U406 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n353) );
  XNOR2_X1 U407 ( .A(G8GAT), .B(KEYINPUT77), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U411 ( .A(n359), .B(n358), .Z(n407) );
  XOR2_X1 U412 ( .A(KEYINPUT74), .B(G162GAT), .Z(n421) );
  XNOR2_X1 U413 ( .A(n421), .B(n360), .ZN(n362) );
  AND2_X1 U414 ( .A1(G232GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n368) );
  INV_X1 U416 ( .A(n368), .ZN(n366) );
  XOR2_X1 U417 ( .A(G92GAT), .B(G106GAT), .Z(n364) );
  XNOR2_X1 U418 ( .A(G50GAT), .B(G99GAT), .ZN(n363) );
  XOR2_X1 U419 ( .A(n364), .B(n363), .Z(n367) );
  INV_X1 U420 ( .A(n367), .ZN(n365) );
  NAND2_X1 U421 ( .A1(n366), .A2(n365), .ZN(n370) );
  NAND2_X1 U422 ( .A1(n368), .A2(n367), .ZN(n369) );
  NAND2_X1 U423 ( .A1(n370), .A2(n369), .ZN(n375) );
  XOR2_X1 U424 ( .A(G190GAT), .B(G134GAT), .Z(n449) );
  XOR2_X1 U425 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n372) );
  XNOR2_X1 U426 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n449), .B(n373), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n375), .B(n374), .ZN(n381) );
  XOR2_X1 U430 ( .A(G29GAT), .B(KEYINPUT7), .Z(n377) );
  XNOR2_X1 U431 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n391) );
  XNOR2_X1 U433 ( .A(G43GAT), .B(n391), .ZN(n379) );
  INV_X1 U434 ( .A(G36GAT), .ZN(n378) );
  INV_X1 U435 ( .A(KEYINPUT101), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n479), .B(n382), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n383), .B(KEYINPUT36), .ZN(n491) );
  NOR2_X1 U438 ( .A1(n407), .A2(n491), .ZN(n385) );
  XNOR2_X1 U439 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n402) );
  XNOR2_X1 U441 ( .A(G43GAT), .B(G15GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n386), .B(G113GAT), .ZN(n441) );
  XNOR2_X1 U443 ( .A(G50GAT), .B(G22GAT), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n387), .B(G141GAT), .ZN(n424) );
  XNOR2_X1 U445 ( .A(n441), .B(n424), .ZN(n401) );
  XOR2_X1 U446 ( .A(G1GAT), .B(n388), .Z(n390) );
  NAND2_X1 U447 ( .A1(G229GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n391), .B(KEYINPUT30), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n392), .B(KEYINPUT66), .ZN(n393) );
  XOR2_X1 U451 ( .A(n394), .B(n393), .Z(n399) );
  XOR2_X1 U452 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n396) );
  XNOR2_X1 U453 ( .A(KEYINPUT67), .B(KEYINPUT65), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U455 ( .A(G169GAT), .B(n397), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U457 ( .A(n401), .B(n400), .Z(n576) );
  XNOR2_X1 U458 ( .A(n576), .B(KEYINPUT70), .ZN(n539) );
  NAND2_X1 U459 ( .A1(n402), .A2(n539), .ZN(n403) );
  NOR2_X1 U460 ( .A1(n580), .A2(n403), .ZN(n404) );
  XOR2_X1 U461 ( .A(KEYINPUT112), .B(n404), .Z(n413) );
  NOR2_X1 U462 ( .A1(n576), .A2(n560), .ZN(n406) );
  INV_X1 U463 ( .A(KEYINPUT46), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n409) );
  INV_X1 U465 ( .A(n479), .ZN(n564) );
  INV_X1 U466 ( .A(n407), .ZN(n585) );
  NOR2_X1 U467 ( .A1(n564), .A2(n585), .ZN(n408) );
  NAND2_X1 U468 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n410), .B(KEYINPUT47), .ZN(n411) );
  XNOR2_X1 U470 ( .A(KEYINPUT111), .B(n411), .ZN(n412) );
  NAND2_X1 U471 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n414), .B(KEYINPUT48), .ZN(n552) );
  NAND2_X1 U473 ( .A1(n527), .A2(n552), .ZN(n416) );
  NOR2_X1 U474 ( .A1(n524), .A2(n417), .ZN(n575) );
  XOR2_X1 U475 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n419) );
  XNOR2_X1 U476 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n434) );
  XOR2_X1 U478 ( .A(n420), .B(G204GAT), .Z(n423) );
  XNOR2_X1 U479 ( .A(G197GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n428) );
  XOR2_X1 U481 ( .A(KEYINPUT88), .B(n424), .Z(n426) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U484 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n469) );
  NAND2_X1 U488 ( .A1(n575), .A2(n469), .ZN(n436) );
  XOR2_X1 U489 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n454) );
  XOR2_X1 U491 ( .A(KEYINPUT80), .B(KEYINPUT82), .Z(n438) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U494 ( .A(n439), .B(KEYINPUT81), .Z(n443) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U497 ( .A(KEYINPUT79), .B(KEYINPUT20), .Z(n445) );
  XNOR2_X1 U498 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U500 ( .A(n447), .B(n446), .Z(n451) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n453), .B(n452), .ZN(n536) );
  AND2_X1 U504 ( .A1(n454), .A2(n536), .ZN(n455) );
  XNOR2_X2 U505 ( .A(n455), .B(KEYINPUT120), .ZN(n570) );
  NAND2_X1 U506 ( .A1(n542), .A2(n570), .ZN(n459) );
  XOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT57), .Z(n457) );
  XOR2_X1 U508 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n456) );
  XNOR2_X1 U509 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U510 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  NAND2_X1 U511 ( .A1(n570), .A2(n564), .ZN(n463) );
  XOR2_X1 U512 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n461) );
  INV_X1 U513 ( .A(G190GAT), .ZN(n460) );
  INV_X1 U514 ( .A(n524), .ZN(n507) );
  NOR2_X1 U515 ( .A1(n539), .A2(n580), .ZN(n464) );
  XOR2_X1 U516 ( .A(KEYINPUT73), .B(n464), .Z(n495) );
  XOR2_X1 U517 ( .A(KEYINPUT27), .B(n527), .Z(n472) );
  NOR2_X1 U518 ( .A1(n507), .A2(n472), .ZN(n551) );
  XNOR2_X1 U519 ( .A(KEYINPUT28), .B(n469), .ZN(n517) );
  NAND2_X1 U520 ( .A1(n551), .A2(n517), .ZN(n538) );
  XOR2_X1 U521 ( .A(n536), .B(KEYINPUT85), .Z(n465) );
  NOR2_X1 U522 ( .A1(n538), .A2(n465), .ZN(n477) );
  NAND2_X1 U523 ( .A1(n536), .A2(n527), .ZN(n466) );
  XOR2_X1 U524 ( .A(KEYINPUT97), .B(n466), .Z(n467) );
  NAND2_X1 U525 ( .A1(n467), .A2(n469), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n468), .B(KEYINPUT25), .ZN(n474) );
  NOR2_X1 U527 ( .A1(n536), .A2(n469), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT96), .B(n470), .Z(n471) );
  XOR2_X1 U529 ( .A(KEYINPUT26), .B(n471), .Z(n574) );
  INV_X1 U530 ( .A(n574), .ZN(n554) );
  NOR2_X1 U531 ( .A1(n472), .A2(n554), .ZN(n473) );
  NOR2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n475), .A2(n524), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT98), .B(n478), .Z(n493) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n481) );
  NAND2_X1 U537 ( .A1(n479), .A2(n585), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(n482) );
  AND2_X1 U539 ( .A1(n493), .A2(n482), .ZN(n506) );
  NAND2_X1 U540 ( .A1(n495), .A2(n506), .ZN(n488) );
  NOR2_X1 U541 ( .A1(n507), .A2(n488), .ZN(n483) );
  XOR2_X1 U542 ( .A(G1GAT), .B(n483), .Z(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(n484), .ZN(G1324GAT) );
  INV_X1 U544 ( .A(n527), .ZN(n511) );
  NOR2_X1 U545 ( .A1(n511), .A2(n488), .ZN(n485) );
  XOR2_X1 U546 ( .A(G8GAT), .B(n485), .Z(G1325GAT) );
  INV_X1 U547 ( .A(n536), .ZN(n513) );
  NOR2_X1 U548 ( .A1(n513), .A2(n488), .ZN(n487) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n517), .A2(n488), .ZN(n490) );
  XNOR2_X1 U552 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(G1327GAT) );
  XNOR2_X1 U554 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n500) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT100), .Z(n498) );
  NOR2_X1 U556 ( .A1(n585), .A2(n491), .ZN(n492) );
  NAND2_X1 U557 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U558 ( .A(KEYINPUT37), .B(n494), .ZN(n521) );
  NAND2_X1 U559 ( .A1(n495), .A2(n521), .ZN(n496) );
  XOR2_X1 U560 ( .A(KEYINPUT38), .B(n496), .Z(n504) );
  NAND2_X1 U561 ( .A1(n504), .A2(n524), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NAND2_X1 U564 ( .A1(n504), .A2(n527), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n504), .A2(n536), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  INV_X1 U569 ( .A(n517), .ZN(n531) );
  NAND2_X1 U570 ( .A1(n504), .A2(n531), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n505), .B(G50GAT), .ZN(G1331GAT) );
  AND2_X1 U572 ( .A1(n576), .A2(n542), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n522), .A2(n506), .ZN(n516) );
  NOR2_X1 U574 ( .A1(n507), .A2(n516), .ZN(n509) );
  XNOR2_X1 U575 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n511), .A2(n516), .ZN(n512) );
  XOR2_X1 U579 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U580 ( .A1(n513), .A2(n516), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n519) );
  XNOR2_X1 U584 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(KEYINPUT107), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n524), .A2(n532), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(KEYINPUT108), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n527), .A2(n532), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U594 ( .A(G99GAT), .B(KEYINPUT109), .Z(n530) );
  NAND2_X1 U595 ( .A1(n532), .A2(n536), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(G1338GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n534) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U600 ( .A(G106GAT), .B(n535), .Z(G1339GAT) );
  XOR2_X1 U601 ( .A(G113GAT), .B(KEYINPUT113), .Z(n541) );
  NAND2_X1 U602 ( .A1(n536), .A2(n552), .ZN(n537) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n548) );
  INV_X1 U604 ( .A(n539), .ZN(n568) );
  NAND2_X1 U605 ( .A1(n548), .A2(n568), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U608 ( .A1(n548), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(n545), .ZN(G1341GAT) );
  NAND2_X1 U611 ( .A1(n585), .A2(n548), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U615 ( .A1(n548), .A2(n564), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  XOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT115), .Z(n556) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n565) );
  INV_X1 U620 ( .A(n565), .ZN(n559) );
  OR2_X1 U621 ( .A1(n559), .A2(n576), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n562) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U627 ( .A(n562), .B(n561), .Z(G1345GAT) );
  NAND2_X1 U628 ( .A1(n585), .A2(n565), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U630 ( .A(G162GAT), .B(KEYINPUT117), .Z(n567) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n570), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G169GAT), .B(n569), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n585), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n588) );
  NOR2_X1 U640 ( .A1(n576), .A2(n588), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n582) );
  INV_X1 U645 ( .A(n588), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(KEYINPUT126), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n491), .A2(n588), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

