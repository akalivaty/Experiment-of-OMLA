

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X2 U324 ( .A(n455), .B(KEYINPUT41), .ZN(n552) );
  XNOR2_X1 U325 ( .A(n348), .B(G57GAT), .ZN(n437) );
  XNOR2_X1 U326 ( .A(G120GAT), .B(G148GAT), .ZN(n348) );
  NOR2_X1 U327 ( .A1(n584), .A2(n410), .ZN(n411) );
  XNOR2_X1 U328 ( .A(KEYINPUT97), .B(n403), .ZN(n546) );
  XOR2_X1 U329 ( .A(n346), .B(KEYINPUT3), .Z(n292) );
  NOR2_X1 U330 ( .A1(n457), .A2(n579), .ZN(n458) );
  XNOR2_X1 U331 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U332 ( .A(n437), .B(n436), .ZN(n439) );
  INV_X1 U333 ( .A(KEYINPUT73), .ZN(n445) );
  NOR2_X1 U334 ( .A1(n545), .A2(n521), .ZN(n469) );
  XNOR2_X1 U335 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U336 ( .A(n468), .B(n467), .ZN(n545) );
  XOR2_X1 U337 ( .A(n396), .B(n385), .Z(n472) );
  XNOR2_X1 U338 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U339 ( .A(n476), .B(n475), .ZN(n477) );
  NOR2_X1 U340 ( .A1(n523), .A2(n477), .ZN(n566) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n452) );
  XNOR2_X1 U342 ( .A(n451), .B(KEYINPUT38), .ZN(n503) );
  XNOR2_X1 U343 ( .A(n479), .B(G176GAT), .ZN(n480) );
  XNOR2_X1 U344 ( .A(n452), .B(KEYINPUT40), .ZN(n453) );
  XNOR2_X1 U345 ( .A(n481), .B(n480), .ZN(G1349GAT) );
  XNOR2_X1 U346 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n294) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n388) );
  XOR2_X1 U350 ( .A(G113GAT), .B(KEYINPUT0), .Z(n349) );
  XOR2_X1 U351 ( .A(n388), .B(n349), .Z(n296) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U354 ( .A(G71GAT), .B(KEYINPUT20), .Z(n298) );
  XNOR2_X1 U355 ( .A(G15GAT), .B(G120GAT), .ZN(n297) );
  XNOR2_X1 U356 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U357 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U358 ( .A(G99GAT), .B(G190GAT), .Z(n302) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G134GAT), .ZN(n301) );
  XNOR2_X1 U360 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U361 ( .A(G127GAT), .B(G176GAT), .Z(n304) );
  XNOR2_X1 U362 ( .A(KEYINPUT83), .B(G183GAT), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n523) );
  XNOR2_X1 U366 ( .A(G29GAT), .B(G134GAT), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n309), .B(KEYINPUT78), .ZN(n360) );
  XOR2_X1 U368 ( .A(n360), .B(G106GAT), .Z(n311) );
  NAND2_X1 U369 ( .A1(G232GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n311), .B(n310), .ZN(n327) );
  XOR2_X1 U371 ( .A(KEYINPUT77), .B(KEYINPUT65), .Z(n313) );
  XNOR2_X1 U372 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U374 ( .A(n314), .B(KEYINPUT9), .Z(n316) );
  XOR2_X1 U375 ( .A(G99GAT), .B(G85GAT), .Z(n438) );
  XNOR2_X1 U376 ( .A(G218GAT), .B(n438), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U378 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n318) );
  XNOR2_X1 U379 ( .A(G162GAT), .B(G92GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U381 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U382 ( .A(G43GAT), .B(G50GAT), .Z(n322) );
  XNOR2_X1 U383 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n429) );
  XNOR2_X1 U385 ( .A(G36GAT), .B(G190GAT), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n323), .B(KEYINPUT79), .ZN(n387) );
  XNOR2_X1 U387 ( .A(n429), .B(n387), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n559) );
  XNOR2_X1 U390 ( .A(KEYINPUT36), .B(n559), .ZN(n584) );
  XOR2_X1 U391 ( .A(KEYINPUT81), .B(G64GAT), .Z(n329) );
  XNOR2_X1 U392 ( .A(G155GAT), .B(G57GAT), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U394 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n331) );
  XNOR2_X1 U395 ( .A(KEYINPUT82), .B(KEYINPUT12), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n343) );
  XOR2_X1 U398 ( .A(G1GAT), .B(G127GAT), .Z(n356) );
  XNOR2_X1 U399 ( .A(G22GAT), .B(G15GAT), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n334), .B(KEYINPUT71), .ZN(n428) );
  XOR2_X1 U401 ( .A(n428), .B(KEYINPUT14), .Z(n336) );
  NAND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n356), .B(n337), .ZN(n341) );
  XOR2_X1 U405 ( .A(G71GAT), .B(KEYINPUT13), .Z(n444) );
  XOR2_X1 U406 ( .A(G8GAT), .B(G183GAT), .Z(n390) );
  XOR2_X1 U407 ( .A(n444), .B(n390), .Z(n339) );
  XNOR2_X1 U408 ( .A(G211GAT), .B(G78GAT), .ZN(n338) );
  XNOR2_X1 U409 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U411 ( .A(n343), .B(n342), .ZN(n579) );
  XOR2_X1 U412 ( .A(KEYINPUT91), .B(KEYINPUT2), .Z(n345) );
  XNOR2_X1 U413 ( .A(G162GAT), .B(KEYINPUT90), .ZN(n344) );
  XNOR2_X1 U414 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U415 ( .A(G141GAT), .B(G155GAT), .ZN(n347) );
  XNOR2_X1 U416 ( .A(n292), .B(n347), .ZN(n382) );
  XOR2_X1 U417 ( .A(n437), .B(n349), .Z(n351) );
  NAND2_X1 U418 ( .A1(G225GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U420 ( .A(n382), .B(n352), .ZN(n364) );
  XOR2_X1 U421 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n354) );
  XNOR2_X1 U422 ( .A(KEYINPUT5), .B(KEYINPUT94), .ZN(n353) );
  XNOR2_X1 U423 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U424 ( .A(n355), .B(KEYINPUT96), .Z(n358) );
  XNOR2_X1 U425 ( .A(n356), .B(G85GAT), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U427 ( .A(n359), .B(KEYINPUT95), .Z(n362) );
  XNOR2_X1 U428 ( .A(n360), .B(KEYINPUT1), .ZN(n361) );
  XNOR2_X1 U429 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U430 ( .A(n364), .B(n363), .ZN(n403) );
  XOR2_X1 U431 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n366) );
  XNOR2_X1 U432 ( .A(G218GAT), .B(KEYINPUT88), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U434 ( .A(n367), .B(G211GAT), .Z(n369) );
  XNOR2_X1 U435 ( .A(G197GAT), .B(G204GAT), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n396) );
  XOR2_X1 U437 ( .A(KEYINPUT92), .B(KEYINPUT23), .Z(n371) );
  XNOR2_X1 U438 ( .A(G22GAT), .B(KEYINPUT86), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U440 ( .A(KEYINPUT85), .B(KEYINPUT24), .Z(n373) );
  XNOR2_X1 U441 ( .A(KEYINPUT84), .B(G148GAT), .ZN(n372) );
  XNOR2_X1 U442 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U443 ( .A(n375), .B(n374), .Z(n384) );
  XOR2_X1 U444 ( .A(G106GAT), .B(G78GAT), .Z(n441) );
  XOR2_X1 U445 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n377) );
  XNOR2_X1 U446 ( .A(G50GAT), .B(KEYINPUT87), .ZN(n376) );
  XNOR2_X1 U447 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U448 ( .A(n441), .B(n378), .Z(n380) );
  NAND2_X1 U449 ( .A1(G228GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U450 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n384), .B(n383), .ZN(n385) );
  NAND2_X1 U453 ( .A1(n472), .A2(n523), .ZN(n386) );
  XNOR2_X1 U454 ( .A(n386), .B(KEYINPUT26), .ZN(n570) );
  XNOR2_X1 U455 ( .A(n388), .B(n387), .ZN(n394) );
  XNOR2_X1 U456 ( .A(G176GAT), .B(G92GAT), .ZN(n389) );
  XNOR2_X1 U457 ( .A(n389), .B(G64GAT), .ZN(n440) );
  XOR2_X1 U458 ( .A(n440), .B(n390), .Z(n392) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n521) );
  XNOR2_X1 U463 ( .A(KEYINPUT27), .B(n521), .ZN(n404) );
  NOR2_X1 U464 ( .A1(n570), .A2(n404), .ZN(n548) );
  XNOR2_X1 U465 ( .A(n548), .B(KEYINPUT98), .ZN(n401) );
  NOR2_X1 U466 ( .A1(n523), .A2(n521), .ZN(n397) );
  NOR2_X1 U467 ( .A1(n472), .A2(n397), .ZN(n398) );
  XNOR2_X1 U468 ( .A(n398), .B(KEYINPUT99), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n399), .B(KEYINPUT25), .ZN(n400) );
  NOR2_X1 U470 ( .A1(n401), .A2(n400), .ZN(n402) );
  NOR2_X1 U471 ( .A1(n403), .A2(n402), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n472), .B(KEYINPUT28), .ZN(n495) );
  NOR2_X1 U473 ( .A1(n546), .A2(n495), .ZN(n406) );
  INV_X1 U474 ( .A(n404), .ZN(n405) );
  NAND2_X1 U475 ( .A1(n406), .A2(n405), .ZN(n530) );
  INV_X1 U476 ( .A(n523), .ZN(n531) );
  NOR2_X1 U477 ( .A1(n530), .A2(n531), .ZN(n407) );
  NOR2_X1 U478 ( .A1(n408), .A2(n407), .ZN(n486) );
  NOR2_X1 U479 ( .A1(n579), .A2(n486), .ZN(n409) );
  XNOR2_X1 U480 ( .A(n409), .B(KEYINPUT105), .ZN(n410) );
  XOR2_X1 U481 ( .A(n411), .B(KEYINPUT37), .Z(n412) );
  XNOR2_X1 U482 ( .A(KEYINPUT106), .B(n412), .ZN(n519) );
  XOR2_X1 U483 ( .A(G141GAT), .B(G197GAT), .Z(n414) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(G36GAT), .ZN(n413) );
  XNOR2_X1 U485 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U486 ( .A(G8GAT), .B(G1GAT), .Z(n416) );
  XNOR2_X1 U487 ( .A(G169GAT), .B(G113GAT), .ZN(n415) );
  XNOR2_X1 U488 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U489 ( .A(n418), .B(n417), .Z(n423) );
  XOR2_X1 U490 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n420) );
  NAND2_X1 U491 ( .A1(G229GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U492 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U493 ( .A(KEYINPUT66), .B(n421), .ZN(n422) );
  XNOR2_X1 U494 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U495 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n425) );
  XNOR2_X1 U496 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n424) );
  XNOR2_X1 U497 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U498 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U499 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U500 ( .A(n431), .B(n430), .ZN(n550) );
  XOR2_X1 U501 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n433) );
  XNOR2_X1 U502 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n432) );
  XNOR2_X1 U503 ( .A(n433), .B(n432), .ZN(n450) );
  NAND2_X1 U504 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  INV_X1 U505 ( .A(KEYINPUT33), .ZN(n434) );
  XOR2_X1 U506 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U507 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U508 ( .A(n443), .B(n442), .ZN(n448) );
  XNOR2_X1 U509 ( .A(G204GAT), .B(n444), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n450), .B(n449), .ZN(n455) );
  BUF_X1 U512 ( .A(n455), .Z(n576) );
  NOR2_X1 U513 ( .A1(n550), .A2(n576), .ZN(n488) );
  NAND2_X1 U514 ( .A1(n519), .A2(n488), .ZN(n451) );
  NOR2_X1 U515 ( .A1(n523), .A2(n503), .ZN(n454) );
  NOR2_X1 U516 ( .A1(n550), .A2(n552), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n456), .B(KEYINPUT46), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n458), .B(KEYINPUT114), .ZN(n459) );
  NAND2_X1 U519 ( .A1(n459), .A2(n559), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT47), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n461), .B(KEYINPUT115), .ZN(n466) );
  INV_X1 U522 ( .A(n579), .ZN(n556) );
  NOR2_X1 U523 ( .A1(n584), .A2(n556), .ZN(n462) );
  XOR2_X1 U524 ( .A(KEYINPUT45), .B(n462), .Z(n463) );
  NOR2_X1 U525 ( .A1(n576), .A2(n463), .ZN(n464) );
  NAND2_X1 U526 ( .A1(n464), .A2(n550), .ZN(n465) );
  NAND2_X1 U527 ( .A1(n466), .A2(n465), .ZN(n468) );
  INV_X1 U528 ( .A(KEYINPUT48), .ZN(n467) );
  XNOR2_X1 U529 ( .A(KEYINPUT54), .B(n469), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n470), .A2(n546), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n471), .B(KEYINPUT64), .ZN(n571) );
  NOR2_X1 U532 ( .A1(n472), .A2(n571), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n474) );
  INV_X1 U534 ( .A(KEYINPUT55), .ZN(n473) );
  INV_X1 U535 ( .A(n552), .ZN(n478) );
  NAND2_X1 U536 ( .A1(n566), .A2(n478), .ZN(n481) );
  XOR2_X1 U537 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n479) );
  XOR2_X1 U538 ( .A(KEYINPUT101), .B(KEYINPUT34), .Z(n483) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(KEYINPUT102), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(n490) );
  INV_X1 U541 ( .A(n559), .ZN(n567) );
  NOR2_X1 U542 ( .A1(n567), .A2(n556), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NOR2_X1 U544 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT100), .B(n487), .ZN(n507) );
  NAND2_X1 U546 ( .A1(n488), .A2(n507), .ZN(n496) );
  NOR2_X1 U547 ( .A1(n546), .A2(n496), .ZN(n489) );
  XOR2_X1 U548 ( .A(n490), .B(n489), .Z(G1324GAT) );
  NOR2_X1 U549 ( .A1(n521), .A2(n496), .ZN(n491) );
  XOR2_X1 U550 ( .A(G8GAT), .B(n491), .Z(G1325GAT) );
  NOR2_X1 U551 ( .A1(n523), .A2(n496), .ZN(n493) );
  XNOR2_X1 U552 ( .A(KEYINPUT103), .B(KEYINPUT35), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U554 ( .A(G15GAT), .B(n494), .Z(G1326GAT) );
  INV_X1 U555 ( .A(n495), .ZN(n526) );
  NOR2_X1 U556 ( .A1(n526), .A2(n496), .ZN(n497) );
  XOR2_X1 U557 ( .A(KEYINPUT104), .B(n497), .Z(n498) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(n498), .ZN(G1327GAT) );
  NOR2_X1 U559 ( .A1(n503), .A2(n546), .ZN(n500) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U562 ( .A1(n503), .A2(n521), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1329GAT) );
  NOR2_X1 U565 ( .A1(n526), .A2(n503), .ZN(n504) );
  XOR2_X1 U566 ( .A(KEYINPUT108), .B(n504), .Z(n505) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(n505), .ZN(G1331GAT) );
  INV_X1 U568 ( .A(n550), .ZN(n572) );
  NOR2_X1 U569 ( .A1(n572), .A2(n552), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(KEYINPUT110), .ZN(n518) );
  NAND2_X1 U571 ( .A1(n518), .A2(n507), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n514), .A2(n546), .ZN(n511) );
  XOR2_X1 U573 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n509) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(KEYINPUT111), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n521), .A2(n514), .ZN(n512) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n523), .A2(n514), .ZN(n513) );
  XOR2_X1 U580 ( .A(G71GAT), .B(n513), .Z(G1334GAT) );
  NOR2_X1 U581 ( .A1(n526), .A2(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n525) );
  NOR2_X1 U586 ( .A1(n546), .A2(n525), .ZN(n520) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n521), .A2(n525), .ZN(n522) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n525), .ZN(n524) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U593 ( .A(KEYINPUT113), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n545), .A2(n530), .ZN(n532) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n541) );
  NOR2_X1 U598 ( .A1(n550), .A2(n541), .ZN(n533) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(n533), .Z(n534) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  NOR2_X1 U601 ( .A1(n552), .A2(n541), .ZN(n536) );
  XNOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT117), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  NOR2_X1 U605 ( .A1(n556), .A2(n541), .ZN(n539) );
  XNOR2_X1 U606 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n540), .Z(G1342GAT) );
  NOR2_X1 U609 ( .A1(n559), .A2(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(KEYINPUT51), .B(KEYINPUT119), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U612 ( .A(G134GAT), .B(n544), .Z(G1343GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(KEYINPUT120), .B(n549), .ZN(n560) );
  NOR2_X1 U616 ( .A1(n550), .A2(n560), .ZN(n551) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n551), .Z(G1344GAT) );
  XNOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n554) );
  NOR2_X1 U619 ( .A1(n552), .A2(n560), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n560), .A2(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n566), .A2(n572), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(G183GAT), .B(KEYINPUT125), .Z(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n579), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1351GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n582), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U642 ( .A1(n582), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n582), .A2(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  INV_X1 U647 ( .A(n582), .ZN(n583) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

