

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U550 ( .A(n774), .B(KEYINPUT108), .ZN(n777) );
  OR2_X1 U551 ( .A1(n762), .A2(n761), .ZN(n764) );
  XNOR2_X1 U552 ( .A(n752), .B(KEYINPUT32), .ZN(n753) );
  AND2_X1 U553 ( .A1(n691), .A2(n690), .ZN(n797) );
  NOR2_X2 U554 ( .A1(n733), .A2(n732), .ZN(n739) );
  NAND2_X2 U555 ( .A1(n797), .A2(n799), .ZN(n705) );
  XNOR2_X2 U556 ( .A(n692), .B(KEYINPUT102), .ZN(n744) );
  OR2_X1 U557 ( .A1(n757), .A2(n767), .ZN(n515) );
  AND2_X1 U558 ( .A1(n517), .A2(n822), .ZN(n516) );
  XNOR2_X1 U559 ( .A(KEYINPUT101), .B(n818), .ZN(n517) );
  OR2_X1 U560 ( .A1(n744), .A2(n776), .ZN(n518) );
  INV_X1 U561 ( .A(KEYINPUT26), .ZN(n697) );
  INV_X1 U562 ( .A(KEYINPUT28), .ZN(n713) );
  NAND2_X1 U563 ( .A1(n751), .A2(n750), .ZN(n752) );
  INV_X1 U564 ( .A(KEYINPUT5), .ZN(n538) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n799) );
  XNOR2_X1 U566 ( .A(n538), .B(KEYINPUT78), .ZN(n539) );
  NOR2_X1 U567 ( .A1(n523), .A2(G2105), .ZN(n549) );
  XNOR2_X1 U568 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U569 ( .A(n533), .B(KEYINPUT64), .ZN(n645) );
  INV_X1 U570 ( .A(n546), .ZN(n879) );
  XNOR2_X1 U571 ( .A(n601), .B(n600), .ZN(n972) );
  NOR2_X1 U572 ( .A1(n527), .A2(n526), .ZN(G164) );
  NOR2_X2 U573 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  XOR2_X1 U574 ( .A(KEYINPUT17), .B(n519), .Z(n545) );
  NAND2_X1 U575 ( .A1(n545), .A2(G138), .ZN(n520) );
  XOR2_X1 U576 ( .A(n520), .B(KEYINPUT93), .Z(n522) );
  XNOR2_X1 U577 ( .A(G2104), .B(KEYINPUT65), .ZN(n523) );
  BUF_X1 U578 ( .A(n549), .Z(n880) );
  NAND2_X1 U579 ( .A1(n880), .A2(G102), .ZN(n521) );
  NAND2_X1 U580 ( .A1(n522), .A2(n521), .ZN(n527) );
  AND2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n875) );
  NAND2_X1 U582 ( .A1(G114), .A2(n875), .ZN(n525) );
  AND2_X1 U583 ( .A1(n523), .A2(G2105), .ZN(n876) );
  NAND2_X1 U584 ( .A1(G126), .A2(n876), .ZN(n524) );
  NAND2_X1 U585 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n656) );
  NOR2_X2 U587 ( .A1(G651), .A2(n656), .ZN(n655) );
  NAND2_X1 U588 ( .A1(n655), .A2(G51), .ZN(n528) );
  XOR2_X1 U589 ( .A(KEYINPUT79), .B(n528), .Z(n531) );
  INV_X1 U590 ( .A(G651), .ZN(n535) );
  NOR2_X1 U591 ( .A1(G543), .A2(n535), .ZN(n529) );
  XOR2_X2 U592 ( .A(KEYINPUT1), .B(n529), .Z(n660) );
  NAND2_X1 U593 ( .A1(n660), .A2(G63), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U595 ( .A(KEYINPUT6), .B(n532), .ZN(n542) );
  NOR2_X1 U596 ( .A1(G543), .A2(G651), .ZN(n533) );
  NAND2_X1 U597 ( .A1(G89), .A2(n645), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(KEYINPUT4), .ZN(n537) );
  NOR2_X1 U599 ( .A1(n656), .A2(n535), .ZN(n648) );
  NAND2_X1 U600 ( .A1(G76), .A2(n648), .ZN(n536) );
  NAND2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n540) );
  NOR2_X1 U602 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U603 ( .A(n543), .B(KEYINPUT7), .Z(n544) );
  XNOR2_X1 U604 ( .A(KEYINPUT80), .B(n544), .ZN(G168) );
  XOR2_X1 U605 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  INV_X1 U606 ( .A(n545), .ZN(n546) );
  NAND2_X1 U607 ( .A1(G137), .A2(n879), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G113), .A2(n875), .ZN(n547) );
  AND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n689) );
  NAND2_X1 U610 ( .A1(G101), .A2(n549), .ZN(n550) );
  XNOR2_X1 U611 ( .A(KEYINPUT66), .B(n550), .ZN(n552) );
  INV_X1 U612 ( .A(KEYINPUT23), .ZN(n551) );
  XNOR2_X1 U613 ( .A(n552), .B(n551), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G125), .A2(n876), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U616 ( .A(n555), .B(KEYINPUT67), .ZN(n691) );
  AND2_X1 U617 ( .A1(n689), .A2(n691), .ZN(G160) );
  NAND2_X1 U618 ( .A1(n648), .A2(G72), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G85), .A2(n645), .ZN(n556) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G60), .A2(n660), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G47), .A2(n655), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  OR2_X1 U624 ( .A1(n561), .A2(n560), .ZN(G290) );
  AND2_X1 U625 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G132), .ZN(G219) );
  INV_X1 U628 ( .A(G82), .ZN(G220) );
  NAND2_X1 U629 ( .A1(n648), .A2(G75), .ZN(n563) );
  NAND2_X1 U630 ( .A1(G88), .A2(n645), .ZN(n562) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G62), .A2(n660), .ZN(n565) );
  NAND2_X1 U633 ( .A1(G50), .A2(n655), .ZN(n564) );
  NAND2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U635 ( .A(KEYINPUT89), .B(n566), .Z(n567) );
  NOR2_X1 U636 ( .A1(n568), .A2(n567), .ZN(G166) );
  NAND2_X1 U637 ( .A1(G64), .A2(n660), .ZN(n569) );
  XOR2_X1 U638 ( .A(KEYINPUT68), .B(n569), .Z(n576) );
  NAND2_X1 U639 ( .A1(n648), .A2(G77), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G90), .A2(n645), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U642 ( .A(n572), .B(KEYINPUT9), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G52), .A2(n655), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U645 ( .A1(n576), .A2(n575), .ZN(G171) );
  XOR2_X1 U646 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n578) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n577) );
  XNOR2_X1 U648 ( .A(n578), .B(n577), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n831) );
  NAND2_X1 U650 ( .A1(n831), .A2(G567), .ZN(n579) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  NAND2_X1 U652 ( .A1(G43), .A2(n655), .ZN(n580) );
  XNOR2_X1 U653 ( .A(n580), .B(KEYINPUT72), .ZN(n583) );
  NAND2_X1 U654 ( .A1(G56), .A2(n660), .ZN(n581) );
  XNOR2_X1 U655 ( .A(n581), .B(KEYINPUT14), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n589) );
  NAND2_X1 U657 ( .A1(G81), .A2(n645), .ZN(n584) );
  XNOR2_X1 U658 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U659 ( .A1(G68), .A2(n648), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U661 ( .A(KEYINPUT13), .B(n587), .Z(n588) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n989) );
  NAND2_X1 U663 ( .A1(G860), .A2(n989), .ZN(n590) );
  XOR2_X1 U664 ( .A(KEYINPUT73), .B(n590), .Z(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G79), .A2(n648), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n660), .A2(G66), .ZN(n592) );
  NAND2_X1 U668 ( .A1(G92), .A2(n645), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U670 ( .A(KEYINPUT74), .B(n593), .ZN(n596) );
  NAND2_X1 U671 ( .A1(G54), .A2(n655), .ZN(n594) );
  XNOR2_X1 U672 ( .A(KEYINPUT75), .B(n594), .ZN(n595) );
  NOR2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n601) );
  XNOR2_X1 U675 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n599) );
  XNOR2_X1 U676 ( .A(n599), .B(KEYINPUT15), .ZN(n600) );
  NOR2_X1 U677 ( .A1(n972), .A2(G868), .ZN(n603) );
  INV_X1 U678 ( .A(G868), .ZN(n672) );
  NOR2_X1 U679 ( .A1(n672), .A2(G301), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U681 ( .A1(n655), .A2(G53), .ZN(n604) );
  XOR2_X1 U682 ( .A(KEYINPUT69), .B(n604), .Z(n606) );
  NAND2_X1 U683 ( .A1(n660), .A2(G65), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U685 ( .A(KEYINPUT70), .B(n607), .Z(n611) );
  NAND2_X1 U686 ( .A1(n645), .A2(G91), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n648), .A2(G78), .ZN(n608) );
  AND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(G299) );
  NAND2_X1 U690 ( .A1(G868), .A2(G286), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G299), .A2(n672), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(G297) );
  INV_X1 U693 ( .A(n972), .ZN(n640) );
  INV_X1 U694 ( .A(G860), .ZN(n642) );
  NAND2_X1 U695 ( .A1(G559), .A2(n642), .ZN(n614) );
  XOR2_X1 U696 ( .A(KEYINPUT81), .B(n614), .Z(n615) );
  NAND2_X1 U697 ( .A1(n640), .A2(n615), .ZN(n616) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT16), .ZN(n617) );
  XNOR2_X1 U699 ( .A(KEYINPUT82), .B(n617), .ZN(G148) );
  NAND2_X1 U700 ( .A1(G868), .A2(n640), .ZN(n618) );
  NOR2_X1 U701 ( .A1(G559), .A2(n618), .ZN(n620) );
  AND2_X1 U702 ( .A1(n672), .A2(n989), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U704 ( .A1(n880), .A2(G99), .ZN(n621) );
  XOR2_X1 U705 ( .A(KEYINPUT83), .B(n621), .Z(n623) );
  NAND2_X1 U706 ( .A1(n875), .A2(G111), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U708 ( .A(KEYINPUT84), .B(n624), .ZN(n629) );
  NAND2_X1 U709 ( .A1(G123), .A2(n876), .ZN(n625) );
  XNOR2_X1 U710 ( .A(n625), .B(KEYINPUT18), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n879), .A2(G135), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n925) );
  XNOR2_X1 U714 ( .A(G2096), .B(n925), .ZN(n631) );
  INV_X1 U715 ( .A(G2100), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n631), .A2(n630), .ZN(G156) );
  NAND2_X1 U717 ( .A1(n645), .A2(G93), .ZN(n632) );
  XNOR2_X1 U718 ( .A(n632), .B(KEYINPUT86), .ZN(n635) );
  NAND2_X1 U719 ( .A1(G80), .A2(n648), .ZN(n633) );
  XOR2_X1 U720 ( .A(KEYINPUT87), .B(n633), .Z(n634) );
  NAND2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G67), .A2(n660), .ZN(n637) );
  NAND2_X1 U723 ( .A1(G55), .A2(n655), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n638) );
  OR2_X1 U725 ( .A1(n639), .A2(n638), .ZN(n673) );
  NAND2_X1 U726 ( .A1(n640), .A2(G559), .ZN(n641) );
  XNOR2_X1 U727 ( .A(n641), .B(n989), .ZN(n670) );
  NAND2_X1 U728 ( .A1(n642), .A2(n670), .ZN(n643) );
  XNOR2_X1 U729 ( .A(n643), .B(KEYINPUT85), .ZN(n644) );
  XOR2_X1 U730 ( .A(n673), .B(n644), .Z(G145) );
  NAND2_X1 U731 ( .A1(n660), .A2(G61), .ZN(n647) );
  NAND2_X1 U732 ( .A1(G86), .A2(n645), .ZN(n646) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n648), .A2(G73), .ZN(n649) );
  XOR2_X1 U735 ( .A(KEYINPUT2), .B(n649), .Z(n650) );
  NOR2_X1 U736 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U737 ( .A1(n655), .A2(G48), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n653), .A2(n652), .ZN(G305) );
  NAND2_X1 U739 ( .A1(G74), .A2(G651), .ZN(n654) );
  XNOR2_X1 U740 ( .A(n654), .B(KEYINPUT88), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G49), .A2(n655), .ZN(n658) );
  NAND2_X1 U742 ( .A1(G87), .A2(n656), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U744 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U745 ( .A1(n662), .A2(n661), .ZN(G288) );
  XOR2_X1 U746 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n664) );
  XOR2_X1 U747 ( .A(KEYINPUT19), .B(n673), .Z(n663) );
  XNOR2_X1 U748 ( .A(n664), .B(n663), .ZN(n667) );
  INV_X1 U749 ( .A(G299), .ZN(n711) );
  XNOR2_X1 U750 ( .A(n711), .B(G305), .ZN(n665) );
  XNOR2_X1 U751 ( .A(n665), .B(G288), .ZN(n666) );
  XNOR2_X1 U752 ( .A(n667), .B(n666), .ZN(n669) );
  XNOR2_X1 U753 ( .A(G290), .B(G166), .ZN(n668) );
  XNOR2_X1 U754 ( .A(n669), .B(n668), .ZN(n899) );
  XOR2_X1 U755 ( .A(n899), .B(n670), .Z(n671) );
  NOR2_X1 U756 ( .A1(n672), .A2(n671), .ZN(n675) );
  NOR2_X1 U757 ( .A1(G868), .A2(n673), .ZN(n674) );
  NOR2_X1 U758 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U759 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U760 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U761 ( .A1(G2090), .A2(n677), .ZN(n679) );
  XNOR2_X1 U762 ( .A(KEYINPUT92), .B(KEYINPUT21), .ZN(n678) );
  XNOR2_X1 U763 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U764 ( .A1(G2072), .A2(n680), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n681) );
  XOR2_X1 U767 ( .A(KEYINPUT22), .B(n681), .Z(n682) );
  NOR2_X1 U768 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G96), .A2(n683), .ZN(n835) );
  NAND2_X1 U770 ( .A1(n835), .A2(G2106), .ZN(n687) );
  NAND2_X1 U771 ( .A1(G120), .A2(G69), .ZN(n684) );
  NOR2_X1 U772 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U773 ( .A1(G108), .A2(n685), .ZN(n836) );
  NAND2_X1 U774 ( .A1(n836), .A2(G567), .ZN(n686) );
  NAND2_X1 U775 ( .A1(n687), .A2(n686), .ZN(n837) );
  NAND2_X1 U776 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U777 ( .A1(n837), .A2(n688), .ZN(n834) );
  NAND2_X1 U778 ( .A1(n834), .A2(G36), .ZN(G176) );
  INV_X1 U779 ( .A(G166), .ZN(G303) );
  INV_X1 U780 ( .A(KEYINPUT33), .ZN(n758) );
  AND2_X1 U781 ( .A1(n689), .A2(G40), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n705), .A2(G8), .ZN(n692) );
  NOR2_X1 U783 ( .A1(n744), .A2(G1966), .ZN(n734) );
  NAND2_X1 U784 ( .A1(G1348), .A2(n705), .ZN(n694) );
  INV_X1 U785 ( .A(n705), .ZN(n718) );
  NAND2_X1 U786 ( .A1(G2067), .A2(n718), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n702) );
  NAND2_X1 U788 ( .A1(n972), .A2(n702), .ZN(n696) );
  NAND2_X1 U789 ( .A1(G1341), .A2(n705), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n701) );
  XOR2_X1 U791 ( .A(G1996), .B(KEYINPUT104), .Z(n957) );
  NOR2_X1 U792 ( .A1(n705), .A2(n957), .ZN(n698) );
  XNOR2_X1 U793 ( .A(n698), .B(n697), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n699), .A2(n989), .ZN(n700) );
  NOR2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n972), .A2(n702), .ZN(n703) );
  NOR2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n718), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U799 ( .A(n706), .B(KEYINPUT27), .ZN(n708) );
  AND2_X1 U800 ( .A1(G1956), .A2(n705), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n716) );
  NOR2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U805 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U807 ( .A(n717), .B(KEYINPUT29), .ZN(n723) );
  NOR2_X1 U808 ( .A1(n718), .A2(G1961), .ZN(n719) );
  XOR2_X1 U809 ( .A(KEYINPUT103), .B(n719), .Z(n721) );
  XOR2_X1 U810 ( .A(KEYINPUT25), .B(G2078), .Z(n948) );
  NOR2_X1 U811 ( .A1(n948), .A2(n705), .ZN(n720) );
  NOR2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n728) );
  NOR2_X1 U813 ( .A1(G301), .A2(n728), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n733) );
  NOR2_X1 U815 ( .A1(n705), .A2(G2084), .ZN(n735) );
  INV_X1 U816 ( .A(n735), .ZN(n724) );
  NAND2_X1 U817 ( .A1(G8), .A2(n724), .ZN(n725) );
  OR2_X1 U818 ( .A1(n734), .A2(n725), .ZN(n726) );
  XNOR2_X1 U819 ( .A(n726), .B(KEYINPUT30), .ZN(n727) );
  NOR2_X1 U820 ( .A1(G168), .A2(n727), .ZN(n730) );
  AND2_X1 U821 ( .A1(G301), .A2(n728), .ZN(n729) );
  NOR2_X1 U822 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U823 ( .A(n731), .B(KEYINPUT31), .ZN(n732) );
  NOR2_X1 U824 ( .A1(n734), .A2(n739), .ZN(n737) );
  NAND2_X1 U825 ( .A1(G8), .A2(n735), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U827 ( .A(KEYINPUT105), .B(n738), .ZN(n754) );
  INV_X1 U828 ( .A(n739), .ZN(n742) );
  AND2_X1 U829 ( .A1(G286), .A2(G8), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n751) );
  INV_X1 U831 ( .A(G8), .ZN(n749) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n705), .ZN(n743) );
  XNOR2_X1 U833 ( .A(n743), .B(KEYINPUT106), .ZN(n746) );
  NOR2_X1 U834 ( .A1(n744), .A2(G1971), .ZN(n745) );
  NOR2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n747), .A2(G303), .ZN(n748) );
  OR2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X2 U838 ( .A1(n754), .A2(n753), .ZN(n762) );
  NAND2_X1 U839 ( .A1(G8), .A2(G166), .ZN(n755) );
  NOR2_X1 U840 ( .A1(G2090), .A2(n755), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n762), .A2(n756), .ZN(n757) );
  INV_X1 U842 ( .A(n744), .ZN(n767) );
  NAND2_X1 U843 ( .A1(n758), .A2(n515), .ZN(n766) );
  NOR2_X1 U844 ( .A1(G288), .A2(G1976), .ZN(n759) );
  XOR2_X1 U845 ( .A(n759), .B(KEYINPUT107), .Z(n768) );
  NOR2_X1 U846 ( .A1(G1971), .A2(G303), .ZN(n760) );
  NOR2_X1 U847 ( .A1(n768), .A2(n760), .ZN(n984) );
  INV_X1 U848 ( .A(n984), .ZN(n761) );
  NAND2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n980) );
  AND2_X1 U850 ( .A1(n767), .A2(n980), .ZN(n763) );
  AND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n773) );
  XOR2_X1 U853 ( .A(G1981), .B(G305), .Z(n975) );
  AND2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U855 ( .A1(KEYINPUT33), .A2(n769), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n975), .A2(n770), .ZN(n771) );
  AND2_X1 U857 ( .A1(n515), .A2(n771), .ZN(n772) );
  OR2_X2 U858 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XOR2_X1 U860 ( .A(n775), .B(KEYINPUT24), .Z(n776) );
  NAND2_X1 U861 ( .A1(n777), .A2(n518), .ZN(n812) );
  NAND2_X1 U862 ( .A1(n875), .A2(G117), .ZN(n778) );
  XNOR2_X1 U863 ( .A(n778), .B(KEYINPUT96), .ZN(n780) );
  NAND2_X1 U864 ( .A1(G129), .A2(n876), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U866 ( .A(n781), .B(KEYINPUT97), .ZN(n783) );
  NAND2_X1 U867 ( .A1(G141), .A2(n879), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n880), .A2(G105), .ZN(n784) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U872 ( .A(KEYINPUT98), .B(n787), .Z(n892) );
  NAND2_X1 U873 ( .A1(G1996), .A2(n892), .ZN(n795) );
  NAND2_X1 U874 ( .A1(G95), .A2(n880), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G107), .A2(n875), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U877 ( .A1(G131), .A2(n879), .ZN(n791) );
  NAND2_X1 U878 ( .A1(G119), .A2(n876), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n792) );
  OR2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n872) );
  NAND2_X1 U881 ( .A1(G1991), .A2(n872), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U883 ( .A(KEYINPUT99), .B(n796), .Z(n931) );
  INV_X1 U884 ( .A(n797), .ZN(n798) );
  NOR2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n826) );
  NAND2_X1 U886 ( .A1(n931), .A2(n826), .ZN(n800) );
  XOR2_X1 U887 ( .A(KEYINPUT100), .B(n800), .Z(n818) );
  XNOR2_X1 U888 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NAND2_X1 U889 ( .A1(n880), .A2(G104), .ZN(n801) );
  XNOR2_X1 U890 ( .A(n801), .B(KEYINPUT94), .ZN(n803) );
  NAND2_X1 U891 ( .A1(G140), .A2(n879), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U893 ( .A(KEYINPUT34), .B(n804), .ZN(n810) );
  NAND2_X1 U894 ( .A1(n875), .A2(G116), .ZN(n805) );
  XOR2_X1 U895 ( .A(KEYINPUT95), .B(n805), .Z(n807) );
  NAND2_X1 U896 ( .A1(n876), .A2(G128), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U898 ( .A(KEYINPUT35), .B(n808), .Z(n809) );
  NOR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U900 ( .A(KEYINPUT36), .B(n811), .ZN(n893) );
  NOR2_X1 U901 ( .A1(n824), .A2(n893), .ZN(n924) );
  NAND2_X1 U902 ( .A1(n826), .A2(n924), .ZN(n822) );
  NAND2_X1 U903 ( .A1(n812), .A2(n516), .ZN(n813) );
  XNOR2_X1 U904 ( .A(n813), .B(KEYINPUT109), .ZN(n815) );
  XNOR2_X1 U905 ( .A(G1986), .B(G290), .ZN(n981) );
  NAND2_X1 U906 ( .A1(n981), .A2(n826), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n829) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n892), .ZN(n921) );
  NOR2_X1 U909 ( .A1(G1991), .A2(n872), .ZN(n926) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U911 ( .A1(n926), .A2(n816), .ZN(n817) );
  NOR2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U913 ( .A(n819), .B(KEYINPUT110), .ZN(n820) );
  NOR2_X1 U914 ( .A1(n921), .A2(n820), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n824), .A2(n893), .ZN(n935) );
  NAND2_X1 U918 ( .A1(n825), .A2(n935), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U921 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U924 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(G188) );
  XNOR2_X1 U927 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  NOR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n837), .ZN(G319) );
  XOR2_X1 U934 ( .A(G2096), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U935 ( .A(G2090), .B(KEYINPUT112), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U937 ( .A(n840), .B(G2678), .Z(n842) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2100), .Z(n844) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U944 ( .A(G1956), .B(G1966), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1981), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U947 ( .A(n849), .B(G2474), .Z(n851) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U950 ( .A(KEYINPUT41), .B(G1976), .Z(n853) );
  XNOR2_X1 U951 ( .A(G1961), .B(G1971), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G136), .A2(n879), .ZN(n857) );
  NAND2_X1 U955 ( .A1(G112), .A2(n875), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n863) );
  NAND2_X1 U957 ( .A1(G124), .A2(n876), .ZN(n858) );
  XOR2_X1 U958 ( .A(KEYINPUT113), .B(n858), .Z(n859) );
  XNOR2_X1 U959 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G100), .A2(n880), .ZN(n860) );
  NAND2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U962 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U963 ( .A1(G139), .A2(n879), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G103), .A2(n880), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U966 ( .A1(n876), .A2(G127), .ZN(n866) );
  XOR2_X1 U967 ( .A(KEYINPUT115), .B(n866), .Z(n868) );
  NAND2_X1 U968 ( .A1(n875), .A2(G115), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n937) );
  XNOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n872), .B(KEYINPUT116), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n888) );
  NAND2_X1 U975 ( .A1(G118), .A2(n875), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G130), .A2(n876), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n886) );
  NAND2_X1 U978 ( .A1(G142), .A2(n879), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G106), .A2(n880), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U981 ( .A(KEYINPUT114), .B(n883), .Z(n884) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(n884), .ZN(n885) );
  NOR2_X1 U983 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U984 ( .A(n888), .B(n887), .Z(n890) );
  XNOR2_X1 U985 ( .A(G164), .B(G162), .ZN(n889) );
  XNOR2_X1 U986 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n937), .B(n891), .ZN(n895) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U990 ( .A(n925), .B(G160), .Z(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G395) );
  XOR2_X1 U993 ( .A(KEYINPUT117), .B(n899), .Z(n901) );
  XNOR2_X1 U994 ( .A(G171), .B(n972), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n903) );
  XOR2_X1 U996 ( .A(G286), .B(n989), .Z(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G37), .A2(n904), .ZN(G397) );
  XOR2_X1 U999 ( .A(G2451), .B(G2430), .Z(n906) );
  XNOR2_X1 U1000 ( .A(G2438), .B(G2443), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n912) );
  XOR2_X1 U1002 ( .A(G2435), .B(G2454), .Z(n908) );
  XNOR2_X1 U1003 ( .A(G1348), .B(G1341), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1005 ( .A(G2446), .B(G2427), .Z(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1007 ( .A(n912), .B(n911), .Z(n913) );
  NAND2_X1 U1008 ( .A1(G14), .A2(n913), .ZN(n919) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n919), .ZN(G401) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n922), .Z(n933) );
  XOR2_X1 U1021 ( .A(G160), .B(G2084), .Z(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n929) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n927), .B(KEYINPUT118), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(n934), .B(KEYINPUT119), .ZN(n936) );
  NAND2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1030 ( .A(G2072), .B(n937), .Z(n939) );
  XOR2_X1 U1031 ( .A(G164), .B(G2078), .Z(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1033 ( .A(KEYINPUT50), .B(n940), .Z(n941) );
  NOR2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n943), .ZN(n945) );
  INV_X1 U1036 ( .A(KEYINPUT55), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1038 ( .A1(n946), .A2(G29), .ZN(n1026) );
  XOR2_X1 U1039 ( .A(G29), .B(KEYINPUT124), .Z(n970) );
  XOR2_X1 U1040 ( .A(G2090), .B(G35), .Z(n963) );
  XNOR2_X1 U1041 ( .A(KEYINPUT121), .B(G2072), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n947), .B(G33), .ZN(n956) );
  XNOR2_X1 U1043 ( .A(G1991), .B(G25), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G27), .B(n948), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(G28), .A2(n951), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT120), .B(G2067), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(G26), .B(n952), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1051 ( .A(G32), .B(n957), .Z(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1053 ( .A(KEYINPUT122), .B(n960), .Z(n961) );
  XNOR2_X1 U1054 ( .A(n961), .B(KEYINPUT53), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(G34), .B(G2084), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n964), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1059 ( .A(n967), .B(KEYINPUT123), .Z(n968) );
  XNOR2_X1 U1060 ( .A(n968), .B(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n971), .ZN(n1024) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1064 ( .A(G299), .B(G1956), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n972), .B(G1348), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n993) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G168), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n977), .B(KEYINPUT57), .ZN(n988) );
  XNOR2_X1 U1070 ( .A(G1961), .B(G171), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(G1971), .A2(G303), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n986) );
  INV_X1 U1073 ( .A(n980), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1078 ( .A(n989), .B(G1341), .Z(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n1022) );
  INV_X1 U1082 ( .A(G16), .ZN(n1020) );
  XNOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT59), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(n996), .B(G4), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G1341), .B(G19), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(KEYINPUT125), .B(G1956), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(G20), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(KEYINPUT60), .B(n1004), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G21), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G1961), .B(G5), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1016) );
  XNOR2_X1 U1097 ( .A(G1986), .B(G24), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(G1976), .B(KEYINPUT126), .Z(n1011) );
  XNOR2_X1 U1101 ( .A(G23), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1105 ( .A(n1017), .B(KEYINPUT61), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT127), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

