//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT27), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT26), .ZN(new_n192));
  OR2_X1    g006(.A1(new_n190), .A2(KEYINPUT27), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(KEYINPUT27), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(G101), .B1(new_n192), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n196), .A3(G101), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G137), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n203), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n207), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(G137), .ZN(new_n210));
  OAI21_X1  g024(.A(G131), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(G128), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT1), .B1(new_n213), .B2(G146), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(G146), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n212), .A2(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  AND4_X1   g033(.A1(new_n219), .A2(new_n216), .A3(new_n217), .A4(G128), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n208), .B(new_n211), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n203), .A2(new_n207), .A3(new_n205), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n223), .A2(new_n208), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G128), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n216), .A2(new_n217), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT0), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT0), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n229), .A2(new_n234), .A3(KEYINPUT64), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n226), .A2(KEYINPUT0), .A3(G128), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n228), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n221), .B1(new_n224), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT2), .A2(G113), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT2), .A2(G113), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT68), .ZN(new_n242));
  XNOR2_X1  g056(.A(G116), .B(G119), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  AND2_X1   g061(.A1(G116), .A2(G119), .ZN(new_n248));
  NOR2_X1   g062(.A1(G116), .A2(G119), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n247), .B1(new_n250), .B2(new_n245), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT69), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n242), .A2(new_n246), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n238), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n200), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n226), .A2(new_n219), .A3(G128), .ZN(new_n258));
  OR2_X1    g072(.A1(KEYINPUT66), .A2(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT66), .A2(G128), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n259), .A2(new_n260), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n258), .B1(new_n261), .B2(new_n226), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n208), .A4(new_n211), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT65), .B1(new_n224), .B2(new_n237), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n229), .A2(new_n232), .A3(new_n230), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT64), .B1(new_n229), .B2(new_n234), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n223), .A2(new_n208), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .A4(new_n235), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT30), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n237), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n270), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT30), .A3(new_n221), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n254), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n256), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n279), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT70), .B1(new_n279), .B2(KEYINPUT31), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n282), .B(new_n256), .C1(new_n274), .C2(new_n278), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n253), .B1(new_n265), .B2(new_n273), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n238), .B2(new_n254), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n276), .A2(KEYINPUT28), .A3(new_n253), .A4(new_n221), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n200), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n280), .A2(new_n281), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT32), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT71), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n295));
  INV_X1    g109(.A(new_n255), .ZN(new_n296));
  INV_X1    g110(.A(new_n199), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(new_n197), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n265), .A2(new_n273), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT30), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n278), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n295), .B1(new_n304), .B2(new_n282), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n279), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n283), .A2(new_n289), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT32), .A4(new_n292), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n294), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G472), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n298), .B1(new_n284), .B2(new_n288), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n298), .A2(new_n255), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n274), .B2(new_n278), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n253), .B1(new_n276), .B2(new_n221), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n288), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n200), .A2(new_n317), .ZN(new_n321));
  AOI21_X1  g135(.A(G902), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n312), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n292), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n281), .A2(new_n290), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(new_n306), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n324), .B1(new_n327), .B2(KEYINPUT32), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n187), .B1(new_n311), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n308), .A2(new_n292), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT32), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n323), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n332), .A2(KEYINPUT72), .A3(new_n294), .A4(new_n310), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G214), .B1(G237), .B2(G902), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT20), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT92), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(G143), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT18), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT92), .B(G143), .ZN(new_n342));
  OAI221_X1 g156(.A(new_n340), .B1(new_n341), .B2(new_n206), .C1(new_n338), .C2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G125), .ZN(new_n345));
  INV_X1    g159(.A(G125), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G140), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(KEYINPUT75), .A3(G140), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(new_n215), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n345), .A2(new_n347), .A3(new_n215), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n342), .A2(new_n338), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(KEYINPUT92), .B2(new_n213), .ZN(new_n356));
  OAI21_X1  g170(.A(G131), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI221_X1 g171(.A(new_n343), .B1(new_n352), .B2(new_n353), .C1(new_n341), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n351), .A2(KEYINPUT16), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n345), .A2(KEYINPUT16), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(G146), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT19), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n349), .B2(new_n350), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT19), .B1(new_n345), .B2(new_n347), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n215), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(KEYINPUT93), .A3(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n340), .B(new_n206), .C1(new_n338), .C2(new_n342), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n357), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT93), .B1(new_n362), .B2(new_n366), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n358), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G113), .B(G122), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT94), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n369), .B2(KEYINPUT17), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT16), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n349), .B2(new_n350), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n215), .B1(new_n381), .B2(new_n360), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n362), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT17), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n357), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n368), .A2(new_n357), .A3(KEYINPUT94), .A4(new_n385), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n379), .A2(new_n384), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n375), .A3(new_n358), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n377), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(G475), .A2(G902), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n337), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n391), .ZN(new_n393));
  AOI211_X1 g207(.A(KEYINPUT20), .B(new_n393), .C1(new_n377), .C2(new_n389), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G902), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n388), .A2(new_n375), .A3(new_n358), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n375), .B1(new_n388), .B2(new_n358), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G475), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n213), .A2(G128), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT13), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n259), .A2(G143), .A3(new_n260), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G134), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n202), .A3(new_n401), .ZN(new_n407));
  XNOR2_X1  g221(.A(G116), .B(G122), .ZN(new_n408));
  INV_X1    g222(.A(G107), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G122), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G116), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n409), .B1(new_n415), .B2(KEYINPUT14), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n413), .A2(new_n416), .B1(new_n409), .B2(new_n408), .ZN(new_n417));
  INV_X1    g231(.A(new_n407), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n202), .B1(new_n404), .B2(new_n401), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n411), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(KEYINPUT9), .B(G234), .Z(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT78), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(G217), .A3(new_n189), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n421), .A2(new_n424), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT96), .A3(new_n396), .ZN(new_n428));
  INV_X1    g242(.A(G478), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(KEYINPUT15), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n396), .B1(new_n425), .B2(new_n426), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT95), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(KEYINPUT95), .B(new_n396), .C1(new_n425), .C2(new_n426), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n428), .A2(new_n430), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  OAI22_X1  g249(.A1(new_n431), .A2(KEYINPUT96), .B1(KEYINPUT15), .B2(new_n429), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(G234), .A2(G237), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(G952), .A3(new_n189), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(G898), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(G902), .A3(G953), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n395), .A2(new_n400), .A3(new_n437), .A4(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n243), .A2(KEYINPUT5), .ZN(new_n446));
  INV_X1    g260(.A(G113), .ZN(new_n447));
  INV_X1    g261(.A(G116), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g263(.A(G119), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n250), .A2(new_n245), .A3(new_n247), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT69), .B1(new_n241), .B2(new_n243), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n409), .A2(G104), .ZN(new_n456));
  AND2_X1   g270(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n457));
  NOR2_X1   g271(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G101), .ZN(new_n460));
  XNOR2_X1  g274(.A(G104), .B(G107), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n459), .B(new_n460), .C1(new_n457), .C2(new_n461), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n461), .A2(new_n460), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n445), .B1(new_n455), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n462), .A2(new_n463), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n251), .A2(new_n252), .B1(new_n446), .B2(new_n451), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT86), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n455), .A2(new_n464), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G110), .B(G122), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT85), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n472), .B(KEYINPUT8), .Z(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n189), .A2(G224), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n237), .A2(G125), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n218), .A2(new_n220), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n346), .ZN(new_n478));
  AOI221_X4 g292(.A(KEYINPUT87), .B1(KEYINPUT7), .B2(new_n475), .C1(new_n476), .C2(new_n478), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n476), .A2(new_n478), .B1(KEYINPUT7), .B2(new_n475), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n474), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT7), .A4(new_n475), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT89), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n480), .B(new_n481), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n484), .B(KEYINPUT88), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n474), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n466), .A2(new_n467), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n462), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n494));
  OR2_X1    g308(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n495));
  NAND2_X1  g309(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n495), .A2(new_n496), .B1(G104), .B2(new_n409), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n374), .A2(G107), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n457), .B1(new_n456), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n494), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n459), .B(KEYINPUT81), .C1(new_n457), .C2(new_n461), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(G101), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT82), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n459), .B1(new_n461), .B2(new_n457), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n460), .B1(new_n505), .B2(new_n494), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT82), .A3(new_n501), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n493), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT4), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n509), .A3(new_n501), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n254), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n492), .B(new_n471), .C1(new_n508), .C2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n487), .A2(new_n491), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n476), .A2(new_n478), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n514), .B(new_n475), .Z(new_n515));
  OAI21_X1  g329(.A(new_n492), .B1(new_n508), .B2(new_n511), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n471), .B(KEYINPUT84), .Z(new_n517));
  AOI22_X1  g331(.A1(new_n512), .A2(KEYINPUT6), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n516), .A2(KEYINPUT6), .A3(new_n517), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n520), .A3(new_n396), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n513), .A2(new_n520), .A3(KEYINPUT90), .A4(new_n396), .ZN(new_n524));
  OAI21_X1  g338(.A(G210), .B1(G237), .B2(G902), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n525), .B(KEYINPUT91), .Z(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n513), .A2(new_n520), .A3(new_n396), .A4(new_n525), .ZN(new_n528));
  AOI211_X1 g342(.A(new_n336), .B(new_n444), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT22), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(G137), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n381), .A2(new_n360), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n353), .B1(new_n533), .B2(G146), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT76), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT23), .B1(new_n230), .B2(G119), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n450), .B2(G128), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n259), .A2(KEYINPUT23), .A3(G119), .A4(new_n260), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n535), .B1(new_n539), .B2(G110), .ZN(new_n540));
  MUX2_X1   g354(.A(new_n230), .B(new_n212), .S(G119), .Z(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT24), .B(G110), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT73), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n540), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n539), .A2(new_n535), .A3(G110), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n534), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n539), .A2(G110), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n548), .A2(KEYINPUT74), .B1(new_n541), .B2(new_n544), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n383), .C1(KEYINPUT74), .C2(new_n548), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT77), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n551), .B1(new_n547), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n532), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n532), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n547), .A2(new_n550), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(new_n556), .B2(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G217), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(G234), .B2(new_n396), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n558), .A2(G902), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n560), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n554), .A2(new_n396), .A3(new_n557), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n563), .B2(KEYINPUT25), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT25), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n554), .A2(new_n565), .A3(new_n396), .A4(new_n557), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n561), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n423), .A2(new_n396), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G221), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n569), .B(KEYINPUT79), .Z(new_n570));
  INV_X1    g384(.A(KEYINPUT10), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n464), .A2(new_n477), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n230), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n258), .B1(new_n226), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n466), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n572), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n510), .A2(new_n275), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n576), .B(new_n224), .C1(new_n508), .C2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(G110), .B(G140), .ZN(new_n580));
  INV_X1    g394(.A(G227), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G953), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n580), .B(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n576), .B1(new_n508), .B2(new_n577), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n270), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n464), .A2(new_n477), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n575), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n270), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT12), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(KEYINPUT12), .A3(new_n270), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n578), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n584), .A2(new_n586), .B1(new_n594), .B2(new_n583), .ZN(new_n595));
  OAI21_X1  g409(.A(G469), .B1(new_n595), .B2(G902), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT83), .B(G469), .Z(new_n597));
  INV_X1    g411(.A(new_n583), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n586), .B2(new_n578), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n593), .A2(new_n578), .A3(new_n598), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n396), .B(new_n597), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n570), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n334), .A2(new_n529), .A3(new_n567), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  OAI21_X1  g418(.A(G472), .B1(new_n291), .B2(G902), .ZN(new_n605));
  AND4_X1   g419(.A1(new_n330), .A2(new_n602), .A3(new_n567), .A4(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n525), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n521), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n528), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n335), .A3(new_n443), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n400), .B1(new_n392), .B2(new_n394), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n433), .A2(new_n434), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n429), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n411), .A2(new_n420), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT33), .B1(new_n614), .B2(KEYINPUT97), .ZN(new_n615));
  OR3_X1    g429(.A1(new_n615), .A2(new_n426), .A3(new_n425), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n427), .A2(new_n615), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(new_n617), .A3(G478), .A4(new_n396), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n606), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT98), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT34), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G104), .ZN(G6));
  AOI21_X1  g439(.A(new_n392), .B1(KEYINPUT99), .B2(new_n394), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(KEYINPUT99), .B2(new_n394), .ZN(new_n627));
  INV_X1    g441(.A(new_n437), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n400), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n610), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n606), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  AND3_X1   g447(.A1(new_n602), .A2(new_n330), .A3(new_n605), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n564), .A2(new_n566), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n555), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n556), .B(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n560), .A2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n529), .A2(new_n634), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  NOR2_X1   g457(.A1(new_n442), .A2(G900), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT100), .Z(new_n645));
  XOR2_X1   g459(.A(new_n439), .B(KEYINPUT101), .Z(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n627), .A2(new_n400), .A3(new_n628), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT102), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n564), .A2(new_n566), .B1(new_n638), .B2(new_n637), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n329), .B2(new_n333), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n336), .B1(new_n608), .B2(new_n528), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n602), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n649), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  NAND2_X1  g470(.A1(new_n527), .A2(new_n528), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT38), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n274), .A2(new_n278), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n200), .B1(new_n660), .B2(new_n296), .ZN(new_n661));
  INV_X1    g475(.A(new_n314), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n396), .B1(new_n662), .B2(new_n319), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n327), .B2(KEYINPUT32), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n311), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n628), .A2(new_n611), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n640), .A2(new_n336), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n658), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(KEYINPUT103), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n647), .B(KEYINPUT39), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n602), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT40), .Z(new_n674));
  NAND3_X1  g488(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  NAND3_X1  g490(.A1(new_n611), .A2(new_n619), .A3(new_n647), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT104), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n611), .A2(new_n619), .A3(new_n679), .A4(new_n647), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n651), .A2(new_n654), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT105), .B(G146), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G48));
  OR2_X1    g499(.A1(new_n508), .A2(new_n577), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n224), .B1(new_n686), .B2(new_n576), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n583), .B1(new_n687), .B2(new_n579), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n593), .A2(new_n578), .A3(new_n598), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(G469), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n601), .B(new_n569), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n396), .B1(new_n599), .B2(new_n600), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n696), .A2(KEYINPUT106), .A3(new_n601), .A4(new_n569), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n334), .A2(new_n567), .A3(new_n621), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND4_X1  g516(.A1(new_n334), .A2(new_n567), .A3(new_n630), .A4(new_n699), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT107), .B(G116), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G18));
  INV_X1    g519(.A(new_n444), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n706), .A2(new_n652), .A3(new_n694), .A4(new_n697), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n334), .A2(new_n707), .A3(new_n640), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  NAND3_X1  g523(.A1(new_n652), .A2(new_n611), .A3(new_n628), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n304), .A2(new_n282), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n283), .B1(new_n298), .B2(new_n320), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n292), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n567), .A2(new_n443), .A3(new_n605), .A4(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n710), .A2(new_n698), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n414), .ZN(G24));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n605), .A2(new_n713), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n717), .B1(new_n718), .B2(new_n650), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n640), .A2(new_n605), .A3(KEYINPUT108), .A4(new_n713), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n652), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n698), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n723), .A3(new_n682), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(new_n569), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n596), .B2(new_n601), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n528), .A2(new_n335), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n727), .A2(new_n527), .A3(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n334), .A2(new_n567), .A3(new_n682), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n567), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n308), .A2(KEYINPUT32), .A3(new_n292), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n733), .B1(new_n734), .B2(new_n332), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n729), .A3(new_n682), .A4(KEYINPUT42), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  AOI21_X1  g552(.A(new_n733), .B1(new_n329), .B2(new_n333), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n649), .A2(new_n739), .A3(new_n729), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  AND2_X1   g555(.A1(new_n595), .A2(KEYINPUT45), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n595), .B2(KEYINPUT45), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(G469), .B2(G902), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n601), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n569), .A3(new_n672), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT109), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n395), .A2(new_n400), .A3(new_n619), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT43), .Z(new_n752));
  AOI21_X1  g566(.A(new_n650), .B1(new_n330), .B2(new_n605), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(KEYINPUT44), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(KEYINPUT44), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n527), .A2(new_n728), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n750), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  NAND2_X1  g575(.A1(new_n748), .A2(new_n569), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT47), .Z(new_n763));
  NOR3_X1   g577(.A1(new_n334), .A2(new_n567), .A3(new_n681), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n757), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT110), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n344), .ZN(G42));
  OR3_X1    g581(.A1(new_n751), .A2(new_n336), .A3(new_n570), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n696), .A2(new_n601), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n733), .B(new_n768), .C1(KEYINPUT49), .C2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT111), .ZN(new_n771));
  INV_X1    g585(.A(new_n658), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n773));
  INV_X1    g587(.A(new_n769), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n666), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n771), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n710), .A2(new_n698), .A3(new_n714), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n700), .A2(new_n703), .A3(new_n708), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n715), .B1(new_n651), .B2(new_n707), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n700), .A4(new_n703), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT113), .B1(new_n611), .B2(new_n437), .ZN(new_n784));
  MUX2_X1   g598(.A(KEYINPUT113), .B(new_n784), .S(new_n620), .Z(new_n785));
  AOI21_X1  g599(.A(new_n336), .B1(new_n527), .B2(new_n528), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n606), .A2(new_n785), .A3(new_n786), .A4(new_n443), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n603), .A2(new_n641), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n758), .B1(new_n596), .B2(new_n601), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n726), .B(new_n681), .C1(new_n719), .C2(new_n720), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n570), .B1(new_n646), .B2(new_n645), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n627), .A2(new_n400), .A3(new_n437), .A4(new_n791), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n650), .B(new_n792), .C1(new_n329), .C2(new_n333), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n789), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n737), .A2(new_n788), .A3(new_n740), .A4(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n783), .A2(new_n795), .A3(KEYINPUT114), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n779), .A2(new_n782), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n737), .A2(new_n788), .A3(new_n740), .A4(new_n794), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n655), .A2(new_n724), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n650), .A2(new_n647), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT116), .ZN(new_n805));
  INV_X1    g619(.A(new_n710), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n666), .A3(new_n806), .A4(new_n727), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n655), .A2(KEYINPUT115), .A3(new_n724), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n803), .A2(new_n808), .A3(new_n683), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n807), .A2(new_n655), .A3(new_n683), .A4(new_n724), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n796), .A2(new_n800), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n811), .B(new_n812), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n796), .A2(new_n800), .A3(KEYINPUT53), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n815), .A2(KEYINPUT117), .A3(new_n816), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n778), .A2(new_n816), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n825), .B(new_n799), .C1(new_n810), .C2(new_n813), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n796), .A2(new_n800), .A3(new_n820), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(new_n816), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n823), .A2(KEYINPUT54), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n646), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n752), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n831), .A2(new_n733), .A3(new_n718), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n774), .A2(new_n570), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n757), .B(new_n832), .C1(new_n763), .C2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n832), .A2(new_n336), .A3(new_n772), .A4(new_n699), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT50), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n699), .A2(new_n757), .ZN(new_n838));
  OR4_X1    g652(.A1(new_n439), .A2(new_n838), .A3(new_n733), .A4(new_n666), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n611), .A3(new_n619), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n831), .A2(new_n838), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT119), .Z(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n721), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n835), .A2(new_n841), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n844), .A2(new_n735), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT48), .Z(new_n851));
  NAND2_X1  g665(.A1(new_n189), .A2(G952), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n832), .B2(new_n723), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n620), .B2(new_n839), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n829), .A2(new_n848), .A3(new_n849), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(G952), .A2(G953), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n776), .B1(new_n856), .B2(new_n857), .ZN(G75));
  NOR2_X1   g672(.A1(new_n189), .A2(G952), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n516), .A2(KEYINPUT6), .A3(new_n517), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n516), .A2(new_n517), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT120), .Z(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT55), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(new_n515), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n828), .A2(new_n396), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(G210), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n526), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n866), .A2(new_n869), .ZN(new_n872));
  AOI211_X1 g686(.A(new_n859), .B(new_n870), .C1(new_n871), .C2(new_n872), .ZN(G51));
  XNOR2_X1  g687(.A(new_n828), .B(new_n824), .ZN(new_n874));
  NAND2_X1  g688(.A1(G469), .A2(G902), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT57), .Z(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n599), .B2(new_n600), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n867), .A2(new_n744), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n859), .B1(new_n878), .B2(new_n879), .ZN(G54));
  NAND2_X1  g694(.A1(KEYINPUT58), .A2(G475), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT121), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n867), .A2(new_n390), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n390), .B1(new_n867), .B2(new_n882), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n884), .A3(new_n859), .ZN(G60));
  NAND2_X1  g699(.A1(G478), .A2(G902), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT59), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n822), .A2(new_n821), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT117), .B1(new_n815), .B2(new_n816), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT54), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n828), .A2(new_n824), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n617), .A2(new_n616), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT122), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT123), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n896));
  INV_X1    g710(.A(new_n894), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n896), .B(new_n897), .C1(new_n829), .C2(new_n887), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n887), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n859), .B1(new_n874), .B2(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n895), .A2(new_n898), .A3(new_n900), .ZN(G63));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT61), .ZN(new_n903));
  OAI22_X1  g717(.A1(new_n902), .A2(KEYINPUT61), .B1(new_n189), .B2(G952), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n827), .A2(new_n816), .ZN(new_n905));
  INV_X1    g719(.A(new_n826), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT60), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n907), .A2(KEYINPUT124), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n828), .B2(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n904), .B1(new_n914), .B2(new_n637), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n911), .A2(new_n558), .A3(new_n913), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n903), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT124), .B1(new_n907), .B2(new_n910), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n828), .A2(new_n912), .A3(new_n909), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n637), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n904), .ZN(new_n921));
  AND4_X1   g735(.A1(new_n903), .A2(new_n920), .A3(new_n916), .A4(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n917), .A2(new_n922), .ZN(G66));
  NAND3_X1  g737(.A1(new_n441), .A2(G224), .A3(G953), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n783), .A2(new_n788), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n864), .B1(G898), .B2(new_n189), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n926), .B(new_n927), .Z(G69));
  NAND2_X1  g742(.A1(new_n302), .A2(new_n277), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n364), .A2(new_n365), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n929), .B(new_n930), .Z(new_n931));
  NAND3_X1  g745(.A1(new_n750), .A2(new_n806), .A3(new_n735), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n765), .A2(new_n932), .A3(new_n760), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n803), .A2(new_n683), .A3(new_n809), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n933), .A2(new_n737), .A3(new_n740), .A4(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(G953), .ZN(new_n936));
  INV_X1    g750(.A(G900), .ZN(new_n937));
  OR3_X1    g751(.A1(new_n937), .A2(KEYINPUT126), .A3(G227), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n189), .B1(KEYINPUT126), .B2(new_n937), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n931), .B(new_n936), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n934), .A2(new_n675), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n765), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n673), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n739), .A2(new_n946), .A3(new_n757), .A4(new_n785), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n760), .A2(new_n189), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n941), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n940), .B1(new_n949), .B2(new_n931), .ZN(G72));
  NAND2_X1  g764(.A1(G472), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT63), .Z(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT127), .Z(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n935), .B2(new_n925), .ZN(new_n954));
  INV_X1    g768(.A(new_n315), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n859), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n760), .A2(new_n783), .A3(new_n788), .A4(new_n947), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n953), .B1(new_n945), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n661), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n952), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n661), .A2(new_n955), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n960), .B1(new_n823), .B2(new_n962), .ZN(G57));
endmodule


