//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT72), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n208), .A2(new_n209), .A3(G134gat), .A4(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G127gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT70), .B1(new_n212), .B2(G134gat), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n212), .A2(KEYINPUT70), .A3(G134gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n209), .B1(new_n218), .B2(G134gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n207), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n206), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NOR4_X1   g026(.A1(KEYINPUT69), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(new_n227), .B2(new_n226), .ZN(new_n230));
  OAI221_X1 g029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT27), .B(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G183gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT27), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT27), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G183gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n239), .A3(new_n234), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n240), .A2(new_n241), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n231), .A2(new_n235), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT24), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(G183gat), .A3(G190gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(new_n227), .B2(KEYINPUT23), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT23), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n252), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n227), .A2(KEYINPUT23), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(G169gat), .A3(G176gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n249), .A2(new_n254), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT25), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n255), .A2(new_n225), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n263), .A2(new_n254), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n263), .B2(new_n254), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n267));
  INV_X1    g066(.A(new_n248), .ZN(new_n268));
  OR3_X1    g067(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n267), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n265), .A2(new_n266), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n224), .B1(new_n262), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G227gat), .ZN(new_n275));
  INV_X1    g074(.A(G233gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n225), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(new_n251), .B2(new_n253), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n264), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n254), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT66), .ZN(new_n282));
  INV_X1    g081(.A(new_n270), .ZN(new_n283));
  NOR3_X1   g082(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT25), .B1(new_n285), .B2(new_n248), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n287), .A2(new_n223), .A3(new_n261), .A4(new_n243), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n274), .A2(new_n277), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT32), .ZN(new_n290));
  XOR2_X1   g089(.A(G15gat), .B(G43gat), .Z(new_n291));
  XNOR2_X1  g090(.A(G71gat), .B(G99gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT34), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n274), .A2(new_n288), .ZN(new_n298));
  INV_X1    g097(.A(new_n277), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI211_X1 g099(.A(KEYINPUT34), .B(new_n277), .C1(new_n274), .C2(new_n288), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n296), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n296), .A2(new_n300), .A3(new_n301), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n290), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n300), .A2(new_n301), .ZN(new_n306));
  INV_X1    g105(.A(new_n296), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n290), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n302), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT36), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n305), .A2(KEYINPUT36), .A3(new_n310), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT5), .ZN(new_n316));
  NAND2_X1  g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT2), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT78), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n320), .A3(KEYINPUT2), .ZN(new_n321));
  AND2_X1   g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  OR2_X1    g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G141gat), .ZN(new_n332));
  INV_X1    g131(.A(G148gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n318), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n328), .A2(new_n317), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n325), .A2(new_n331), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n220), .A2(new_n338), .A3(new_n222), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT80), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n220), .A2(new_n338), .A3(new_n341), .A4(new_n222), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n331), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(new_n337), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n223), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n340), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n316), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(KEYINPUT3), .A2(new_n345), .B1(new_n220), .B2(new_n222), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n338), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT79), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n335), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n320), .B1(new_n317), .B2(KEYINPUT2), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n330), .B1(new_n357), .B2(new_n321), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n336), .A2(new_n337), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT3), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AND4_X1   g159(.A1(KEYINPUT79), .A2(new_n360), .A3(new_n223), .A4(new_n353), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n348), .B1(new_n354), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n339), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n340), .A2(new_n342), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n364), .B1(new_n365), .B2(KEYINPUT4), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n350), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n339), .A2(new_n363), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n365), .B2(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n360), .A2(new_n223), .A3(new_n353), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n351), .A2(KEYINPUT79), .A3(new_n353), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n369), .A2(new_n316), .A3(new_n374), .A4(new_n348), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT0), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  AOI21_X1  g179(.A(KEYINPUT6), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n367), .A2(new_n375), .ZN(new_n382));
  INV_X1    g181(.A(new_n380), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT6), .ZN(new_n386));
  AOI211_X1 g185(.A(new_n386), .B(new_n380), .C1(new_n367), .C2(new_n375), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G211gat), .B(G218gat), .ZN(new_n393));
  INV_X1    g192(.A(G197gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT73), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G197gat), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n395), .A2(new_n397), .A3(G204gat), .ZN(new_n398));
  AOI21_X1  g197(.A(G204gat), .B1(new_n395), .B2(new_n397), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n402));
  OAI21_X1  g201(.A(G211gat), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT22), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n393), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n395), .A2(new_n397), .A3(G204gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n395), .A2(new_n397), .ZN(new_n408));
  INV_X1    g207(.A(G204gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND4_X1   g209(.A1(new_n405), .A2(new_n407), .A3(new_n410), .A4(new_n393), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G226gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(new_n276), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n286), .B1(new_n279), .B2(new_n264), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n243), .B(new_n261), .C1(new_n415), .C2(new_n265), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT75), .B(KEYINPUT29), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n414), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n242), .A2(new_n235), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n421), .A2(new_n231), .B1(KEYINPUT25), .B2(new_n260), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n422), .B2(new_n287), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n412), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n407), .A3(new_n410), .ZN(new_n425));
  INV_X1    g224(.A(new_n393), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n400), .A2(new_n405), .A3(new_n393), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n416), .A2(new_n414), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT29), .B1(new_n422), .B2(new_n287), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n429), .B(new_n430), .C1(new_n431), .C2(new_n414), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n424), .A2(new_n432), .A3(KEYINPUT76), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT76), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(new_n412), .C1(new_n419), .C2(new_n423), .ZN(new_n435));
  AOI211_X1 g234(.A(KEYINPUT30), .B(new_n392), .C1(new_n433), .C2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n433), .A2(new_n435), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n391), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n433), .A2(new_n435), .A3(new_n392), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(KEYINPUT30), .A3(new_n440), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n385), .A2(new_n388), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT31), .B(G50gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G228gat), .A2(G233gat), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n418), .B1(new_n406), .B2(new_n411), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n338), .B1(new_n449), .B2(new_n352), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n417), .B1(new_n338), .B2(new_n352), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n429), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n448), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G22gat), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT29), .B1(new_n427), .B2(new_n428), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n345), .B1(new_n455), .B2(KEYINPUT3), .ZN(new_n456));
  INV_X1    g255(.A(new_n451), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n412), .ZN(new_n458));
  INV_X1    g257(.A(new_n448), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n453), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n454), .B1(new_n453), .B2(new_n460), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n447), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n417), .B1(new_n427), .B2(new_n428), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n345), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n459), .B1(new_n466), .B2(new_n458), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT29), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n406), .B2(new_n411), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n338), .B1(new_n469), .B2(new_n352), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n459), .B1(new_n451), .B2(new_n429), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(G22gat), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(KEYINPUT82), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n447), .B1(new_n473), .B2(new_n461), .ZN(new_n475));
  OAI22_X1  g274(.A1(new_n464), .A2(new_n474), .B1(new_n475), .B2(KEYINPUT81), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n467), .A2(new_n472), .A3(G22gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n446), .B1(new_n477), .B2(new_n462), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT81), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n443), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n479), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n462), .A2(new_n463), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n473), .A2(KEYINPUT82), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n447), .A4(new_n461), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n475), .A2(KEYINPUT81), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n482), .A2(new_n485), .A3(KEYINPUT83), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n315), .B1(new_n442), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n382), .A2(KEYINPUT85), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n367), .A2(new_n491), .A3(new_n375), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n383), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(KEYINPUT40), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n347), .A2(new_n349), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT39), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n369), .A2(new_n374), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(new_n349), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT39), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n500), .A3(new_n349), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n380), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n495), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n498), .A2(new_n349), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n504), .A2(KEYINPUT39), .A3(new_n496), .ZN(new_n505));
  INV_X1    g304(.A(new_n495), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n505), .A2(new_n380), .A3(new_n506), .A4(new_n501), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n493), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n441), .A2(new_n437), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT86), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n387), .B1(new_n493), .B2(new_n381), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n512));
  AOI21_X1  g311(.A(new_n391), .B1(new_n438), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n433), .A2(KEYINPUT37), .A3(new_n435), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT38), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n392), .B1(new_n433), .B2(new_n435), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT37), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n431), .A2(new_n414), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n423), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n518), .B1(new_n520), .B2(new_n412), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n429), .B1(new_n419), .B2(new_n423), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT38), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n517), .B1(new_n513), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n511), .A2(new_n516), .A3(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n510), .A2(new_n525), .A3(new_n488), .ZN(new_n526));
  OR3_X1    g325(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT86), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n489), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n529));
  INV_X1    g328(.A(new_n311), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n488), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g330(.A(KEYINPUT89), .B(new_n311), .C1(new_n481), .C2(new_n487), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n442), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT35), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT35), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n440), .A2(KEYINPUT30), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n536), .A2(new_n517), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n537), .B2(new_n436), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(new_n511), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n311), .B1(new_n481), .B2(new_n487), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT88), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT88), .B1(new_n539), .B2(new_n540), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n528), .B1(new_n534), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G15gat), .B(G22gat), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G1gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547));
  INV_X1    g346(.A(G1gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(KEYINPUT16), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G8gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT90), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n546), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n550), .A2(KEYINPUT90), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n552), .B(new_n553), .Z(new_n554));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n552), .B(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT91), .ZN(new_n558));
  INV_X1    g357(.A(G36gat), .ZN(new_n559));
  AND2_X1   g358(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G29gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n565), .A2(KEYINPUT15), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(KEYINPUT15), .ZN(new_n567));
  XNOR2_X1  g366(.A(G43gat), .B(G50gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT17), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(new_n569), .B2(new_n570), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n556), .B(new_n558), .C1(new_n572), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n571), .A2(new_n557), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT18), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n576), .B(KEYINPUT13), .Z(new_n582));
  NOR2_X1   g381(.A1(new_n571), .A2(new_n557), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT92), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n571), .B(new_n557), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n582), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n575), .A2(KEYINPUT18), .A3(new_n576), .A4(new_n578), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n581), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(G197gat), .ZN(new_n593));
  XOR2_X1   g392(.A(KEYINPUT11), .B(G169gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT12), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n579), .A2(new_n580), .B1(new_n585), .B2(new_n588), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n596), .B1(new_n599), .B2(new_n590), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n544), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT7), .ZN(new_n604));
  NAND2_X1  g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605));
  INV_X1    g404(.A(G85gat), .ZN(new_n606));
  INV_X1    g405(.A(G92gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(KEYINPUT8), .A2(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G99gat), .B(G106gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n571), .A2(new_n611), .B1(KEYINPUT41), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n572), .A2(new_n574), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n611), .B(KEYINPUT97), .Z(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n619), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT95), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT96), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n618), .A2(new_n621), .A3(new_n627), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G57gat), .B(G64gat), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G71gat), .B(G78gat), .Z(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT21), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT20), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n554), .B1(new_n639), .B2(new_n638), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT94), .ZN(new_n647));
  XOR2_X1   g446(.A(G127gat), .B(G155gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G183gat), .B(G211gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n645), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n638), .B(new_n611), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n611), .A2(KEYINPUT10), .A3(new_n637), .A4(new_n636), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G230gat), .A2(G233gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT99), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  OAI211_X1 g464(.A(new_n662), .B(new_n665), .C1(new_n654), .C2(new_n661), .ZN(new_n666));
  INV_X1    g465(.A(new_n665), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n660), .B1(new_n656), .B2(new_n657), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n654), .A2(new_n661), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n666), .A2(KEYINPUT100), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n672), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n631), .A2(new_n653), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n602), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n385), .A2(new_n388), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(new_n548), .ZN(G1324gat));
  NOR2_X1   g479(.A1(new_n677), .A2(new_n509), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n550), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT101), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT101), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT16), .B(G8gat), .Z(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n681), .B2(new_n686), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n681), .A2(new_n685), .A3(new_n686), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n683), .B(new_n684), .C1(new_n687), .C2(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(G15gat), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n677), .A2(new_n690), .A3(new_n315), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n677), .A2(new_n311), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(G15gat), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT102), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(KEYINPUT102), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n691), .B1(new_n694), .B2(new_n695), .ZN(G1326gat));
  NOR2_X1   g495(.A1(new_n677), .A2(new_n488), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n653), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n675), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n630), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n623), .B2(new_n628), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n602), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n678), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n563), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n706), .A2(KEYINPUT103), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT103), .B1(new_n706), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n442), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n488), .A2(new_n530), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT89), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n540), .A2(new_n529), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n543), .B1(new_n718), .B2(new_n535), .ZN(new_n719));
  INV_X1    g518(.A(new_n528), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n704), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(KEYINPUT105), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(KEYINPUT105), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n544), .B2(new_n704), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n591), .A2(new_n597), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n599), .A2(new_n596), .A3(new_n590), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n730), .A2(KEYINPUT104), .A3(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n702), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G29gat), .B1(new_n739), .B2(new_n678), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n709), .A2(KEYINPUT45), .A3(new_n710), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n713), .A2(new_n740), .A3(new_n741), .ZN(G1328gat));
  INV_X1    g541(.A(new_n706), .ZN(new_n743));
  INV_X1    g542(.A(new_n509), .ZN(new_n744));
  AOI21_X1  g543(.A(G36gat), .B1(KEYINPUT106), .B2(KEYINPUT46), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G36gat), .B1(new_n739), .B2(new_n509), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(new_n315), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n729), .A2(G43gat), .A3(new_n751), .A4(new_n738), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  INV_X1    g552(.A(G43gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n706), .B2(new_n311), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n752), .A2(KEYINPUT107), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n752), .A2(KEYINPUT107), .A3(new_n755), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(new_n753), .ZN(G1330gat));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759));
  INV_X1    g558(.A(new_n738), .ZN(new_n760));
  AOI211_X1 g559(.A(new_n488), .B(new_n760), .C1(new_n725), .C2(new_n728), .ZN(new_n761));
  INV_X1    g560(.A(G50gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n488), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n743), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n761), .B2(new_n762), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n763), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  OAI221_X1 g567(.A(new_n765), .B1(new_n759), .B2(KEYINPUT48), .C1(new_n761), .C2(new_n762), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(G1331gat));
  NAND3_X1  g569(.A1(new_n700), .A2(new_n704), .A3(new_n675), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n544), .A2(new_n736), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n707), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n744), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT49), .B(G64gat), .Z(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(G1333gat));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n530), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n780));
  AOI21_X1  g579(.A(G71gat), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n772), .A2(KEYINPUT109), .A3(new_n530), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n772), .A2(G71gat), .A3(new_n751), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT50), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(G1334gat));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n764), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g590(.A1(new_n737), .A2(KEYINPUT110), .A3(new_n653), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n700), .B2(new_n736), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT88), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n386), .B1(new_n382), .B2(new_n383), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n380), .B1(new_n382), .B2(KEYINPUT85), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n492), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n509), .B(new_n535), .C1(new_n799), .C2(new_n387), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n796), .B1(new_n715), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT88), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(KEYINPUT35), .B2(new_n533), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n631), .B(new_n795), .C1(new_n804), .C2(new_n528), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n721), .A2(KEYINPUT51), .A3(new_n795), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n809), .A2(new_n606), .A3(new_n707), .A4(new_n675), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n675), .ZN(new_n811));
  AOI211_X1 g610(.A(new_n678), .B(new_n811), .C1(new_n725), .C2(new_n728), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n812), .B2(new_n606), .ZN(G1336gat));
  NOR2_X1   g612(.A1(new_n509), .A2(G92gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n809), .A2(new_n675), .A3(new_n814), .ZN(new_n815));
  AOI211_X1 g614(.A(new_n509), .B(new_n811), .C1(new_n725), .C2(new_n728), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n815), .B(KEYINPUT111), .C1(new_n816), .C2(new_n607), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT52), .ZN(new_n818));
  INV_X1    g617(.A(new_n811), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n729), .A2(new_n744), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G92gat), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n821), .A2(KEYINPUT111), .A3(new_n822), .A4(new_n815), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n818), .A2(new_n823), .ZN(G1337gat));
  INV_X1    g623(.A(G99gat), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n825), .A3(new_n530), .A4(new_n675), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n315), .B(new_n811), .C1(new_n725), .C2(new_n728), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n827), .B2(new_n825), .ZN(G1338gat));
  NOR2_X1   g627(.A1(new_n488), .A2(G106gat), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT51), .B1(new_n721), .B2(new_n795), .ZN(new_n830));
  INV_X1    g629(.A(new_n795), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n544), .A2(new_n806), .A3(new_n704), .A4(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n675), .B(new_n829), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT112), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n809), .A2(new_n835), .A3(new_n675), .A4(new_n829), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n719), .A2(new_n720), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n837), .A2(new_n631), .B1(new_n726), .B2(new_n724), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n544), .A2(new_n704), .A3(new_n723), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n764), .B(new_n819), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G106gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n834), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT53), .ZN(new_n843));
  XNOR2_X1  g642(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n833), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1339gat));
  NOR4_X1   g645(.A1(new_n631), .A2(new_n736), .A3(new_n653), .A4(new_n675), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n576), .B1(new_n575), .B2(new_n578), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n586), .A2(new_n582), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n595), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n731), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n656), .A2(new_n657), .A3(new_n660), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n662), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n665), .B1(new_n668), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n854), .A2(KEYINPUT55), .A3(new_n856), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n859), .A2(new_n666), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n631), .A2(new_n852), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n674), .A2(new_n851), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n863), .B1(new_n736), .B2(new_n861), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n864), .B2(new_n631), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n847), .B1(new_n865), .B2(new_n653), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n764), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n678), .A2(new_n744), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n530), .A3(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n869), .A2(new_n204), .A3(new_n601), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n531), .A2(new_n532), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n866), .A2(new_n678), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n509), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n736), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n870), .B1(new_n875), .B2(new_n204), .ZN(G1340gat));
  NOR3_X1   g675(.A1(new_n869), .A2(new_n202), .A3(new_n674), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n675), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n202), .ZN(G1341gat));
  NAND3_X1  g678(.A1(new_n874), .A2(new_n218), .A3(new_n700), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n869), .A2(new_n653), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n218), .B2(new_n881), .ZN(G1342gat));
  NAND2_X1  g681(.A1(new_n631), .A2(new_n509), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT114), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(G134gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n872), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n887));
  OAI21_X1  g686(.A(G134gat), .B1(new_n869), .B2(new_n704), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G1343gat));
  NAND2_X1  g689(.A1(new_n868), .A2(new_n315), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n488), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n859), .A2(new_n666), .A3(new_n860), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n601), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n704), .B1(new_n896), .B2(new_n863), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n862), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n653), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n676), .A2(new_n737), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n894), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n892), .B1(new_n866), .B2(new_n488), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT115), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT115), .B(new_n892), .C1(new_n866), .C2(new_n488), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n891), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n332), .B1(new_n906), .B2(new_n736), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n866), .A2(new_n678), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n764), .A2(new_n315), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT116), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n601), .A2(G141gat), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n908), .A2(new_n509), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT58), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n735), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT104), .B1(new_n730), .B2(new_n731), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n861), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n863), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n631), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n704), .A2(new_n851), .A3(new_n895), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n653), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n488), .B1(new_n921), .B2(new_n900), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n903), .B1(new_n922), .B2(KEYINPUT57), .ZN(new_n923));
  INV_X1    g722(.A(new_n901), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n905), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n891), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n732), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G141gat), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT117), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n921), .A2(new_n900), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(new_n707), .A3(new_n910), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n933), .A2(KEYINPUT117), .A3(new_n509), .A4(new_n911), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT58), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n928), .A2(new_n929), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n929), .B1(new_n928), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n914), .B1(new_n936), .B2(new_n937), .ZN(G1344gat));
  INV_X1    g737(.A(new_n933), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n744), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n333), .A3(new_n675), .ZN(new_n941));
  AOI211_X1 g740(.A(KEYINPUT59), .B(new_n333), .C1(new_n906), .C2(new_n675), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT59), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n676), .A2(new_n601), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n488), .B1(new_n899), .B2(new_n944), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n945), .A2(KEYINPUT57), .B1(new_n866), .B2(new_n894), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(new_n675), .A3(new_n926), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n943), .B1(new_n947), .B2(G148gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n941), .B1(new_n942), .B2(new_n948), .ZN(G1345gat));
  AOI21_X1  g748(.A(G155gat), .B1(new_n940), .B2(new_n700), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n700), .A2(G155gat), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT119), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n906), .B2(new_n952), .ZN(G1346gat));
  NOR3_X1   g752(.A1(new_n939), .A2(G162gat), .A3(new_n884), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT120), .Z(new_n955));
  NAND2_X1  g754(.A1(new_n906), .A2(new_n631), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G162gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1347gat));
  NOR2_X1   g757(.A1(new_n707), .A2(new_n509), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n960), .A2(new_n311), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n867), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(G169gat), .A3(new_n732), .ZN(new_n964));
  NOR4_X1   g763(.A1(new_n866), .A2(new_n707), .A3(new_n509), .A4(new_n871), .ZN(new_n965));
  AOI21_X1  g764(.A(G169gat), .B1(new_n965), .B2(new_n736), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n964), .A2(new_n966), .ZN(G1348gat));
  OAI21_X1  g766(.A(G176gat), .B1(new_n962), .B2(new_n674), .ZN(new_n968));
  INV_X1    g767(.A(G176gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n965), .A2(new_n969), .A3(new_n675), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(G1349gat));
  OR3_X1    g770(.A1(new_n962), .A2(KEYINPUT121), .A3(new_n653), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT121), .B1(new_n962), .B2(new_n653), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n972), .A2(G183gat), .A3(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n975), .A2(KEYINPUT60), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n700), .A2(new_n233), .ZN(new_n977));
  AOI22_X1  g776(.A1(new_n965), .A2(new_n977), .B1(new_n975), .B2(KEYINPUT60), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n974), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n976), .B1(new_n974), .B2(new_n978), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n979), .A2(new_n980), .ZN(G1350gat));
  OAI21_X1  g780(.A(G190gat), .B1(new_n962), .B2(new_n704), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT61), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n234), .A3(new_n631), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1351gat));
  NOR2_X1   g784(.A1(new_n866), .A2(new_n707), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n909), .A2(new_n509), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g787(.A(KEYINPUT123), .B(G197gat), .Z(new_n989));
  NOR3_X1   g788(.A1(new_n988), .A2(new_n737), .A3(new_n989), .ZN(new_n990));
  XOR2_X1   g789(.A(new_n990), .B(KEYINPUT124), .Z(new_n991));
  NOR2_X1   g790(.A1(new_n960), .A2(new_n751), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n946), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(new_n732), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(new_n989), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n991), .A2(new_n995), .ZN(G1352gat));
  NOR2_X1   g795(.A1(new_n674), .A2(G204gat), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n986), .A2(new_n987), .A3(new_n997), .ZN(new_n998));
  XOR2_X1   g797(.A(new_n998), .B(KEYINPUT62), .Z(new_n999));
  NAND3_X1  g798(.A1(new_n946), .A2(new_n675), .A3(new_n992), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n946), .A2(KEYINPUT125), .A3(new_n675), .A4(new_n992), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1002), .A2(G204gat), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(KEYINPUT126), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n999), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1006), .A2(new_n1008), .ZN(G1353gat));
  OR3_X1    g808(.A1(new_n988), .A2(G211gat), .A3(new_n653), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n700), .ZN(new_n1011));
  AND3_X1   g810(.A1(new_n1011), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1012));
  AOI21_X1  g811(.A(KEYINPUT63), .B1(new_n1011), .B2(G211gat), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(G1354gat));
  OAI211_X1 g813(.A(new_n993), .B(new_n631), .C1(new_n402), .C2(new_n401), .ZN(new_n1015));
  INV_X1    g814(.A(G218gat), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1016), .B1(new_n988), .B2(new_n704), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


