//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1267, new_n1268,
    new_n1269;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI211_X1 g034(.A(G137), .B(new_n457), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT66), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n460), .A2(KEYINPUT66), .A3(new_n463), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT65), .B1(new_n469), .B2(new_n457), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n458), .A2(new_n459), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G2105), .ZN(new_n475));
  AOI211_X1 g050(.A(new_n464), .B(new_n465), .C1(new_n470), .C2(new_n475), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT68), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n471), .A2(new_n457), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(G124), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  OR3_X1    g058(.A1(new_n471), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT67), .B1(new_n471), .B2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n482), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n487), .B(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n458), .C2(new_n459), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n458), .B2(new_n459), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n468), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G543), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n503), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n503), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(G651), .B1(G50), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n516), .B(new_n504), .C1(new_n507), .C2(new_n508), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT70), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n505), .A2(new_n506), .A3(G543), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n519), .A2(new_n520), .B1(KEYINPUT5), .B2(new_n503), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(new_n516), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n518), .A2(G88), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n515), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(G166));
  AND3_X1   g101(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n514), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n518), .A2(new_n523), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(G89), .ZN(G168));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n509), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n535), .B1(new_n538), .B2(KEYINPUT72), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n539), .B1(KEYINPUT72), .B2(new_n538), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n518), .A2(G90), .A3(new_n523), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n514), .A2(G52), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND2_X1  g122(.A1(new_n533), .A2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n509), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G651), .B1(G43), .B2(new_n514), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  OAI211_X1 g134(.A(G65), .B(new_n504), .C1(new_n507), .C2(new_n508), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n535), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(KEYINPUT6), .A2(G651), .ZN(new_n563));
  NOR2_X1   g138(.A1(KEYINPUT6), .A2(G651), .ZN(new_n564));
  OAI211_X1 g139(.A(G53), .B(G543), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT75), .B1(new_n566), .B2(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n518), .A2(G91), .A3(new_n523), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n572), .A2(KEYINPUT76), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT76), .B1(new_n572), .B2(new_n573), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(new_n532), .ZN(new_n577));
  INV_X1    g152(.A(G89), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n518), .A2(new_n523), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(G286));
  AND3_X1   g155(.A1(new_n518), .A2(G88), .A3(new_n523), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n514), .A2(G50), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(new_n535), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT77), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n515), .A2(new_n586), .A3(new_n524), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n585), .A2(new_n587), .ZN(G303));
  INV_X1    g163(.A(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n509), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n514), .A2(KEYINPUT78), .A3(G49), .ZN(new_n594));
  AOI22_X1  g169(.A1(G651), .A2(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n518), .A2(G87), .A3(new_n523), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n595), .A2(KEYINPUT79), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT79), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(G288));
  NAND2_X1  g174(.A1(new_n514), .A2(G48), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI211_X1 g176(.A(G61), .B(new_n504), .C1(new_n507), .C2(new_n508), .ZN(new_n602));
  NAND2_X1  g177(.A1(G73), .A2(G543), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n601), .B1(new_n604), .B2(G651), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n518), .A2(G86), .A3(new_n523), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G305));
  NAND2_X1  g182(.A1(new_n533), .A2(G85), .ZN(new_n608));
  NAND2_X1  g183(.A1(G72), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G60), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n509), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(KEYINPUT80), .B(G47), .Z(new_n612));
  AOI22_X1  g187(.A1(new_n611), .A2(G651), .B1(new_n514), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(G290));
  XOR2_X1   g189(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n579), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n518), .A2(new_n523), .A3(G92), .A4(new_n615), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT82), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n509), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n623), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G171), .B2(new_n626), .ZN(G284));
  OAI21_X1  g203(.A(new_n627), .B1(G171), .B2(new_n626), .ZN(G321));
  NAND2_X1  g204(.A1(G299), .A2(new_n626), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n626), .B2(G168), .ZN(G297));
  OAI21_X1  g206(.A(new_n630), .B1(new_n626), .B2(G168), .ZN(G280));
  INV_X1    g207(.A(new_n625), .ZN(new_n633));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G860), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT83), .Z(G148));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n468), .A2(new_n462), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT12), .Z(new_n642));
  XOR2_X1   g217(.A(KEYINPUT84), .B(KEYINPUT13), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n645), .A2(G2100), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT85), .Z(new_n647));
  INV_X1    g222(.A(G2096), .ZN(new_n648));
  INV_X1    g223(.A(new_n486), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G135), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n651));
  INV_X1    g226(.A(G111), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(G2105), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n481), .B2(G123), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  AOI22_X1  g231(.A1(new_n645), .A2(G2100), .B1(new_n648), .B2(new_n656), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n647), .B(new_n657), .C1(new_n648), .C2(new_n656), .ZN(G156));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT86), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT14), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2427), .B(G2438), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2430), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT15), .B(G2435), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n667), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n663), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(G14), .B1(new_n670), .B2(new_n672), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(G401));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT87), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(G2072), .A2(G2078), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n442), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n677), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT18), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(KEYINPUT17), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(new_n677), .A3(new_n678), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n678), .B1(new_n677), .B2(new_n681), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(new_n677), .B2(new_n684), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n683), .B(new_n685), .C1(new_n688), .C2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G2096), .B(G2100), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G227));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1971), .B(G1976), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT19), .ZN(new_n697));
  XOR2_X1   g272(.A(G1956), .B(G2474), .Z(new_n698));
  XOR2_X1   g273(.A(G1961), .B(G1966), .Z(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n698), .A2(new_n699), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(new_n705), .B(new_n704), .S(new_n697), .Z(new_n706));
  OR3_X1    g281(.A1(new_n703), .A2(new_n706), .A3(KEYINPUT89), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n708));
  OAI21_X1  g283(.A(KEYINPUT89), .B1(new_n703), .B2(new_n706), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(new_n714));
  OR3_X1    g289(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n713), .B1(new_n711), .B2(new_n714), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1991), .B(G1996), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT91), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n715), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n719), .B1(new_n715), .B2(new_n716), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n695), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n722), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n724), .A2(new_n694), .A3(new_n720), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n725), .ZN(G229));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n633), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G4), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G1348), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(KEYINPUT92), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(KEYINPUT92), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(G35), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n736), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT29), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI211_X1 g315(.A(KEYINPUT29), .B(new_n737), .C1(G162), .C2(new_n736), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G2090), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n731), .B(new_n732), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G32), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n649), .A2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n481), .A2(G129), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT99), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT26), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n753), .A2(new_n754), .B1(G105), .B2(new_n462), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n747), .A2(new_n750), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n746), .B1(new_n756), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT100), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n758), .B(new_n759), .Z(new_n760));
  NOR2_X1   g335(.A1(G168), .A2(new_n727), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n727), .B2(G21), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT102), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n457), .A2(G103), .A3(G2104), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT25), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n770));
  INV_X1    g345(.A(G139), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n769), .B1(new_n457), .B2(new_n770), .C1(new_n486), .C2(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G33), .B(new_n772), .S(G29), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2072), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n498), .A2(new_n500), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n490), .A2(new_n493), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(new_n736), .ZN(new_n778));
  INV_X1    g353(.A(new_n736), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G27), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G2078), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT31), .B(G11), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT30), .B(G28), .Z(new_n786));
  OAI221_X1 g361(.A(new_n785), .B1(G29), .B2(new_n786), .C1(new_n655), .C2(new_n779), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n774), .A2(new_n783), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(G34), .ZN(new_n790));
  OR3_X1    g365(.A1(new_n790), .A2(KEYINPUT98), .A3(new_n736), .ZN(new_n791));
  OAI21_X1  g366(.A(KEYINPUT98), .B1(new_n790), .B2(new_n736), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n789), .A2(G34), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G160), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n733), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2084), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n760), .A2(new_n766), .A3(new_n788), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n762), .A2(new_n763), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT101), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n743), .B1(new_n740), .B2(new_n741), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n744), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n649), .A2(G131), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT93), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  INV_X1    g382(.A(G107), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G2105), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n481), .B2(G119), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(new_n736), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n779), .A2(G25), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G24), .B(G290), .S(G16), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1986), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n813), .B1(new_n812), .B2(new_n814), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n816), .A2(new_n818), .A3(new_n819), .A4(KEYINPUT95), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n727), .A2(G22), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G166), .B2(new_n727), .ZN(new_n822));
  INV_X1    g397(.A(G1971), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n596), .ZN(new_n825));
  MUX2_X1   g400(.A(G23), .B(new_n825), .S(G16), .Z(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT33), .B(G1976), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT94), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(G6), .A2(G16), .ZN(new_n830));
  INV_X1    g405(.A(G305), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(G16), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT32), .B(G1981), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n824), .A2(new_n829), .A3(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n820), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(G16), .A2(G19), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n554), .B2(G16), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(G1341), .Z(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n765), .B2(new_n764), .ZN(new_n844));
  NAND2_X1  g419(.A1(G299), .A2(G16), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n727), .A2(G20), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT23), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G1956), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n727), .A2(G5), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(G171), .B2(new_n727), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G1961), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n779), .A2(G26), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT28), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n855));
  INV_X1    g430(.A(G116), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n856), .B2(G2105), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(new_n481), .B2(G128), .ZN(new_n858));
  INV_X1    g433(.A(G140), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n486), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT96), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n854), .B1(new_n861), .B2(new_n733), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G2067), .ZN(new_n863));
  NOR4_X1   g438(.A1(new_n844), .A2(new_n849), .A3(new_n852), .A4(new_n863), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n820), .A2(KEYINPUT36), .A3(new_n836), .A4(new_n837), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n803), .A2(new_n840), .A3(new_n864), .A4(new_n865), .ZN(G150));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n867));
  XNOR2_X1  g442(.A(G150), .B(new_n867), .ZN(G311));
  NAND3_X1  g443(.A1(new_n518), .A2(G93), .A3(new_n523), .ZN(new_n869));
  NAND2_X1  g444(.A1(G80), .A2(G543), .ZN(new_n870));
  INV_X1    g445(.A(G67), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n509), .B2(new_n871), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n872), .A2(G651), .B1(G55), .B2(new_n514), .ZN(new_n873));
  AND4_X1   g448(.A1(new_n548), .A2(new_n552), .A3(new_n869), .A4(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n869), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n514), .A2(G55), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(new_n535), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT104), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n873), .A2(new_n880), .A3(new_n869), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n874), .B1(new_n882), .B2(new_n553), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT38), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n625), .A2(new_n634), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n887));
  AOI21_X1  g462(.A(G860), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n887), .B2(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n882), .A2(G860), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT105), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n892), .ZN(G145));
  NAND2_X1  g468(.A1(G162), .A2(new_n656), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(G162), .A2(new_n656), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n795), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n894), .A3(G160), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n811), .A2(new_n642), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n756), .B(new_n772), .ZN(new_n902));
  INV_X1    g477(.A(new_n642), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n806), .A2(new_n903), .A3(new_n810), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n902), .B1(new_n901), .B2(new_n904), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n860), .B(KEYINPUT96), .Z(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n777), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n861), .A2(G164), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n649), .A2(G142), .ZN(new_n911));
  OAI21_X1  g486(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n912));
  INV_X1    g487(.A(G118), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(G2105), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n914), .B1(new_n481), .B2(G130), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n909), .B2(new_n910), .ZN(new_n919));
  OAI22_X1  g494(.A1(new_n906), .A2(new_n907), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n907), .ZN(new_n921));
  INV_X1    g496(.A(new_n919), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n917), .A4(new_n905), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n900), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n900), .A3(new_n920), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT106), .B1(new_n930), .B2(new_n924), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(G395));
  XNOR2_X1  g509(.A(G166), .B(G290), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n825), .B(G305), .Z(new_n936));
  XNOR2_X1  g511(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT42), .ZN(new_n938));
  XNOR2_X1  g513(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n938), .B(KEYINPUT109), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  OR3_X1    g515(.A1(new_n937), .A2(KEYINPUT109), .A3(new_n939), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n881), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n880), .B1(new_n873), .B2(new_n869), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n553), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n548), .A2(new_n552), .A3(new_n869), .A4(new_n873), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(new_n637), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n624), .A2(new_n619), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n618), .B(new_n949), .C1(new_n574), .C2(new_n575), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n572), .A2(new_n573), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT76), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n572), .A2(KEYINPUT76), .A3(new_n573), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n625), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT41), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n950), .B2(new_n955), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n950), .A2(new_n955), .A3(new_n958), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n942), .B(new_n957), .C1(new_n962), .C2(new_n948), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n957), .B1(new_n962), .B2(new_n948), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n940), .A2(new_n941), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n626), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n882), .A2(new_n626), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT110), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n942), .B(new_n964), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n970), .B(new_n967), .C1(new_n971), .C2(new_n626), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n969), .A2(new_n972), .ZN(G295));
  OAI21_X1  g548(.A(new_n967), .B1(new_n971), .B2(new_n626), .ZN(G331));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n975));
  NAND2_X1  g550(.A1(G301), .A2(G286), .ZN(new_n976));
  OAI211_X1 g551(.A(G168), .B(new_n540), .C1(new_n544), .C2(new_n545), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n883), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n947), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n950), .A2(new_n955), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n979), .A2(KEYINPUT111), .A3(new_n947), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT111), .B1(new_n979), .B2(new_n947), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n979), .A2(new_n947), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n959), .B1(new_n988), .B2(new_n961), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n956), .A2(new_n988), .A3(KEYINPUT41), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n983), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n937), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n975), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n980), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n979), .A2(new_n947), .A3(KEYINPUT111), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n978), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n961), .A2(new_n988), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n960), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n990), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n982), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1003), .A2(KEYINPUT114), .A3(new_n937), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n995), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n978), .A2(new_n980), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n962), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n984), .A2(new_n985), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n976), .A2(new_n977), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n956), .B1(new_n1010), .B2(new_n883), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1008), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AND4_X1   g587(.A1(new_n1008), .A2(new_n1011), .A3(new_n997), .A4(new_n998), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n937), .B(new_n1007), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n927), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT43), .B1(new_n1005), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1011), .A2(new_n997), .A3(new_n998), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT112), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1009), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1020), .A2(new_n1021), .B1(new_n962), .B2(new_n1006), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1018), .B1(new_n1022), .B2(new_n937), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1017), .B1(new_n1023), .B2(new_n1015), .ZN(new_n1024));
  AOI21_X1  g599(.A(G37), .B1(new_n1022), .B2(new_n937), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1007), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n994), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1025), .A2(KEYINPUT115), .A3(new_n1018), .A4(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1016), .A2(new_n1024), .A3(new_n1028), .A4(KEYINPUT44), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1018), .B1(new_n1005), .B2(new_n1015), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1025), .A2(KEYINPUT43), .A3(new_n1027), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1029), .A2(new_n1033), .ZN(G397));
  NAND2_X1  g609(.A1(new_n470), .A2(new_n475), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n465), .A2(new_n464), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(G40), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT116), .B(G1384), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(G164), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G2067), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n861), .B(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1041), .B1(new_n1043), .B2(new_n756), .ZN(new_n1044));
  INV_X1    g619(.A(G1996), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT46), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT47), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1043), .A2(new_n1041), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT117), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n756), .B(G1996), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n1041), .B2(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n806), .A2(new_n813), .A3(new_n810), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n813), .B1(new_n806), .B2(new_n810), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1041), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(G290), .A2(G1986), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1041), .ZN(new_n1059));
  XOR2_X1   g634(.A(new_n1059), .B(KEYINPUT48), .Z(new_n1060));
  OAI21_X1  g635(.A(new_n1049), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1041), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n861), .A2(new_n1042), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1058), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G290), .A2(G1986), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1062), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1053), .A2(new_n1070), .A3(new_n1056), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1384), .B1(new_n775), .B2(new_n776), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1072), .A2(new_n1035), .A3(G40), .A4(new_n1036), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G8), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G305), .A2(G1981), .ZN(new_n1075));
  INV_X1    g650(.A(G1981), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n605), .A2(new_n606), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1074), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n605), .A2(new_n1076), .A3(new_n606), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1076), .B1(new_n605), .B2(new_n606), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1081), .B1(new_n1084), .B2(KEYINPUT49), .ZN(new_n1085));
  NOR4_X1   g660(.A1(new_n1082), .A2(new_n1083), .A3(KEYINPUT120), .A4(new_n1079), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1080), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G288), .A2(G1976), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1077), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1074), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n595), .A2(G1976), .A3(new_n596), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1073), .A2(new_n1092), .A3(G8), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT52), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n597), .A2(new_n598), .A3(G1976), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1073), .A2(new_n1092), .A3(new_n1096), .A4(G8), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1094), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT120), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1084), .A2(new_n1081), .A3(KEYINPUT49), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1101), .B2(new_n1080), .ZN(new_n1102));
  INV_X1    g677(.A(G8), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT119), .B1(new_n1072), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1384), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n777), .A2(new_n1104), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AND4_X1   g687(.A1(G40), .A2(new_n1035), .A3(new_n743), .A4(new_n1036), .ZN(new_n1113));
  AOI211_X1 g688(.A(KEYINPUT50), .B(G1384), .C1(new_n775), .C2(new_n776), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT118), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1108), .A2(new_n1112), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1038), .B1(G164), .B2(G1384), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1039), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n777), .A2(KEYINPUT45), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n823), .B1(new_n1120), .B2(new_n1037), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1103), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n585), .A2(G8), .A3(new_n587), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT55), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n585), .A2(new_n587), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1090), .A2(new_n1091), .B1(new_n1102), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(G160), .A2(G40), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1072), .A2(new_n1104), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(new_n1114), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1131), .A2(new_n823), .B1(new_n1133), .B2(new_n1113), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1125), .B(new_n1126), .C1(new_n1134), .C2(new_n1103), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1098), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1128), .A2(new_n1135), .A3(new_n1087), .A4(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1035), .A2(G40), .A3(new_n1036), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1108), .A2(new_n1138), .A3(new_n1112), .A4(new_n1115), .ZN(new_n1139));
  INV_X1    g714(.A(G1961), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1120), .A2(G2078), .A3(new_n1037), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1072), .A2(KEYINPUT45), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1138), .A2(new_n1117), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(G2078), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1142), .A2(KEYINPUT53), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(G171), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1137), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G2084), .ZN(new_n1151));
  AND4_X1   g726(.A1(G40), .A2(new_n1035), .A3(new_n1151), .A4(new_n1036), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1108), .A2(new_n1112), .A3(new_n1152), .A4(new_n1115), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1143), .A2(new_n1117), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n763), .B1(new_n1154), .B2(new_n1037), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1153), .A2(G168), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT51), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(G8), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(G168), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1161), .A2(G8), .A3(new_n1156), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1159), .B1(new_n1162), .B2(KEYINPUT51), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1150), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1156), .A2(G8), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT51), .B1(new_n1166), .B2(new_n1160), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1158), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(KEYINPUT62), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1130), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1103), .B(G286), .C1(new_n1153), .C2(new_n1155), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1128), .A2(new_n1171), .A3(KEYINPUT63), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(new_n1122), .B2(KEYINPUT121), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1175), .B(new_n1103), .C1(new_n1116), .C2(new_n1121), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1102), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1172), .B1(new_n1177), .B2(KEYINPUT122), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1179), .B(new_n1102), .C1(new_n1174), .C2(new_n1176), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1102), .A2(new_n1171), .A3(new_n1128), .A4(new_n1135), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1178), .A2(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1170), .A2(new_n1183), .ZN(new_n1184));
  AND4_X1   g759(.A1(new_n1087), .A2(new_n1128), .A3(new_n1136), .A4(new_n1135), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1138), .A2(new_n782), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1072), .A2(KEYINPUT45), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1038), .B(G1384), .C1(new_n775), .C2(new_n776), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1037), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1145), .A2(new_n1186), .B1(new_n1189), .B2(new_n1146), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1190), .A2(G301), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1146), .A2(G40), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1193), .B1(new_n473), .B2(G2105), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1040), .A2(new_n1036), .A3(new_n1194), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1186), .A2(new_n1145), .B1(new_n1195), .B2(new_n1119), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g772(.A(KEYINPUT54), .B(new_n1192), .C1(new_n1197), .C2(G301), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT54), .ZN(new_n1199));
  AND3_X1   g774(.A1(new_n1191), .A2(new_n1196), .A3(G301), .ZN(new_n1200));
  AOI21_X1  g775(.A(G301), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1168), .A2(new_n1185), .A3(new_n1198), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(KEYINPUT126), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1191), .A2(new_n1196), .A3(G301), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1149), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1137), .B1(new_n1199), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1207), .A2(new_n1208), .A3(new_n1168), .A4(new_n1198), .ZN(new_n1209));
  INV_X1    g784(.A(G1956), .ZN(new_n1210));
  OAI21_X1  g785(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1211), .A2(new_n1110), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1210), .B1(new_n1212), .B2(new_n1037), .ZN(new_n1213));
  XNOR2_X1  g788(.A(KEYINPUT56), .B(G2072), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1138), .A2(new_n1117), .A3(new_n1119), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n951), .A2(KEYINPUT57), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT57), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n572), .A2(new_n1217), .A3(new_n573), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1213), .A2(new_n1215), .A3(new_n1216), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1219), .A2(KEYINPUT123), .ZN(new_n1220));
  AND2_X1   g795(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT123), .ZN(new_n1222));
  NAND4_X1  g797(.A1(new_n1221), .A2(new_n1222), .A3(new_n1213), .A4(new_n1215), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1139), .A2(new_n730), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1138), .A2(new_n1042), .A3(new_n1072), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n625), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI22_X1  g802(.A1(new_n1213), .A2(new_n1215), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1224), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g804(.A(KEYINPUT125), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1219), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  NAND4_X1  g806(.A1(new_n1221), .A2(KEYINPUT125), .A3(new_n1213), .A4(new_n1215), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1231), .A2(KEYINPUT61), .A3(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g808(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n1234));
  NAND4_X1  g809(.A1(new_n1138), .A2(new_n1045), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1235));
  XOR2_X1   g810(.A(KEYINPUT58), .B(G1341), .Z(new_n1236));
  NAND2_X1  g811(.A1(new_n1073), .A2(new_n1236), .ZN(new_n1237));
  AOI211_X1 g812(.A(new_n553), .B(new_n1234), .C1(new_n1235), .C2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1239), .A2(new_n554), .ZN(new_n1240));
  NOR2_X1   g815(.A1(KEYINPUT124), .A2(KEYINPUT59), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1238), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g817(.A(new_n1228), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1243));
  OAI211_X1 g818(.A(new_n1233), .B(new_n1242), .C1(KEYINPUT61), .C2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1245));
  INV_X1    g820(.A(KEYINPUT60), .ZN(new_n1246));
  OAI21_X1  g821(.A(new_n633), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g822(.A1(new_n1225), .A2(KEYINPUT60), .A3(new_n625), .A4(new_n1226), .ZN(new_n1248));
  AOI22_X1  g823(.A1(new_n1247), .A2(new_n1248), .B1(new_n1246), .B2(new_n1245), .ZN(new_n1249));
  OAI21_X1  g824(.A(new_n1229), .B1(new_n1244), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g825(.A1(new_n1204), .A2(new_n1209), .A3(new_n1250), .ZN(new_n1251));
  AOI211_X1 g826(.A(KEYINPUT127), .B(new_n1071), .C1(new_n1184), .C2(new_n1251), .ZN(new_n1252));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1182), .A2(new_n1181), .ZN(new_n1255));
  NAND2_X1  g830(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g831(.A(new_n1130), .ZN(new_n1257));
  INV_X1    g832(.A(new_n1169), .ZN(new_n1258));
  NAND4_X1  g833(.A1(new_n1102), .A2(new_n1201), .A3(new_n1128), .A4(new_n1135), .ZN(new_n1259));
  AOI21_X1  g834(.A(new_n1259), .B1(new_n1168), .B2(KEYINPUT62), .ZN(new_n1260));
  AOI21_X1  g835(.A(new_n1257), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g836(.A1(new_n1251), .A2(new_n1256), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g837(.A(new_n1071), .ZN(new_n1263));
  AOI21_X1  g838(.A(new_n1253), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g839(.A(new_n1066), .B1(new_n1252), .B2(new_n1264), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g840(.A(G319), .B1(new_n673), .B2(new_n674), .ZN(new_n1267));
  NOR2_X1   g841(.A1(new_n1267), .A2(G227), .ZN(new_n1268));
  AND3_X1   g842(.A1(new_n723), .A2(new_n725), .A3(new_n1268), .ZN(new_n1269));
  NAND4_X1  g843(.A1(new_n1030), .A2(new_n1269), .A3(new_n932), .A4(new_n1032), .ZN(G225));
  INV_X1    g844(.A(G225), .ZN(G308));
endmodule


