//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n190), .B(new_n192), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT0), .B(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT64), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n193), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n203), .A2(new_n205), .A3(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n200), .B1(new_n210), .B2(new_n199), .ZN(new_n211));
  INV_X1    g025(.A(G953), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G224), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n211), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT4), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G107), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT3), .A3(G104), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT75), .B1(new_n219), .B2(G104), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT75), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n217), .A3(G107), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n215), .B(G101), .C1(new_n221), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G119), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G116), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT66), .B(G119), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G116), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G119), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n236), .A3(G116), .ZN(new_n237));
  INV_X1    g051(.A(new_n228), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(new_n231), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n226), .B1(new_n233), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n218), .A2(new_n220), .ZN(new_n242));
  INV_X1    g056(.A(G101), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(new_n243), .A3(new_n222), .A4(new_n224), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT4), .ZN(new_n245));
  INV_X1    g059(.A(new_n225), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n243), .B1(new_n246), .B2(new_n242), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT80), .B1(new_n241), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(G101), .B1(new_n221), .B2(new_n225), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n230), .A2(new_n232), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n239), .A2(new_n231), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n251), .A2(new_n254), .A3(new_n255), .A4(new_n226), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n249), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n237), .A2(KEYINPUT5), .A3(new_n238), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n234), .A2(new_n236), .A3(new_n260), .A4(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G113), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n252), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n217), .A2(G107), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n219), .A2(G104), .ZN(new_n265));
  OAI21_X1  g079(.A(G101), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n244), .A2(new_n266), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n263), .A2(KEYINPUT81), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT81), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n261), .A2(G113), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n270), .A2(new_n258), .B1(new_n230), .B2(new_n232), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n244), .A2(new_n266), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G122), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n257), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT6), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n257), .A2(new_n274), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n275), .B(KEYINPUT82), .Z(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n279), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n214), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OR3_X1    g097(.A1(new_n263), .A2(KEYINPUT83), .A3(new_n267), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT83), .B1(new_n263), .B2(new_n267), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n284), .B(new_n285), .C1(new_n272), .C2(new_n271), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n275), .B(KEYINPUT8), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n213), .A2(KEYINPUT7), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n211), .B(new_n289), .Z(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n276), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n188), .B1(new_n283), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n214), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n276), .A2(KEYINPUT6), .B1(new_n278), .B2(new_n279), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n279), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n290), .A2(new_n276), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n299), .B2(new_n288), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n300), .A3(new_n187), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n294), .A2(KEYINPUT84), .A3(new_n301), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n283), .A2(new_n188), .A3(new_n293), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT84), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G217), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(G234), .B2(new_n292), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT22), .B(G137), .ZN(new_n313));
  INV_X1    g127(.A(G221), .ZN(new_n314));
  INV_X1    g128(.A(G234), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n314), .A2(new_n315), .A3(G953), .ZN(new_n316));
  XOR2_X1   g130(.A(new_n313), .B(new_n316), .Z(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n322), .A2(KEYINPUT16), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(new_n189), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n189), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n229), .A2(G128), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT72), .B1(new_n196), .B2(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n229), .A2(KEYINPUT72), .A3(G128), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT24), .B(G110), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n328), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G110), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n234), .A2(new_n236), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n196), .ZN(new_n340));
  AOI22_X1  g154(.A1(KEYINPUT73), .A2(new_n340), .B1(new_n329), .B2(KEYINPUT23), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n340), .A2(KEYINPUT73), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n199), .A2(G140), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n322), .A2(new_n347), .A3(new_n189), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n325), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT74), .B(G110), .Z(new_n351));
  NAND3_X1  g165(.A1(new_n343), .A2(new_n344), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n331), .A2(new_n334), .A3(new_n332), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n318), .B1(new_n346), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n343), .A2(new_n344), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n328), .B(new_n336), .C1(new_n356), .C2(new_n338), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n353), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n349), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n359), .A3(new_n317), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(new_n360), .A3(new_n292), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n355), .A2(new_n360), .A3(KEYINPUT25), .A4(new_n292), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n312), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n355), .A2(new_n360), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n311), .A2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n203), .A2(new_n205), .A3(new_n209), .ZN(new_n373));
  INV_X1    g187(.A(G137), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT11), .A3(G134), .ZN(new_n375));
  INV_X1    g189(.A(G134), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G137), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT65), .ZN(new_n379));
  INV_X1    g193(.A(G131), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT11), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n376), .B2(G137), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n378), .A2(new_n379), .A3(new_n380), .A4(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n375), .A3(new_n380), .A4(new_n377), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT65), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n375), .A3(new_n377), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G131), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n373), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n377), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n376), .A2(G137), .ZN(new_n391));
  OAI21_X1  g205(.A(G131), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n195), .A2(new_n392), .A3(new_n197), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n393), .B1(new_n383), .B2(new_n385), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT70), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n198), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n386), .A2(new_n396), .A3(new_n392), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT70), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n383), .A2(new_n385), .B1(G131), .B2(new_n387), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(new_n373), .ZN(new_n400));
  INV_X1    g214(.A(new_n254), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n395), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT28), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n386), .A2(new_n388), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n210), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n401), .B1(new_n406), .B2(new_n397), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n384), .B(new_n379), .ZN(new_n408));
  OAI22_X1  g222(.A1(new_n399), .A2(new_n373), .B1(new_n408), .B2(new_n393), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(new_n254), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT28), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G237), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT67), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT67), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G237), .ZN(new_n415));
  AOI21_X1  g229(.A(G953), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g230(.A(KEYINPUT26), .B(G101), .Z(new_n417));
  AND3_X1   g231(.A1(new_n416), .A2(new_n417), .A3(G210), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n417), .B1(G210), .B2(new_n416), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OR3_X1    g235(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(new_n418), .B2(new_n419), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n404), .A2(new_n411), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n292), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n406), .A2(new_n430), .A3(new_n397), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n409), .A2(KEYINPUT30), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n254), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n406), .A2(new_n401), .A3(new_n397), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT29), .B1(new_n436), .B2(new_n425), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT69), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT69), .B1(new_n422), .B2(new_n423), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n404), .A2(new_n411), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n429), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G472), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT71), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n428), .A2(new_n292), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n401), .B1(new_n431), .B2(new_n432), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n425), .B1(new_n446), .B2(new_n410), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n441), .A2(new_n426), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(G472), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT31), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n434), .A2(new_n453), .A3(new_n424), .A4(new_n435), .ZN(new_n454));
  INV_X1    g268(.A(new_n440), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n254), .B1(new_n409), .B2(KEYINPUT70), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT28), .B1(new_n456), .B2(new_n400), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n409), .A2(new_n254), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n403), .B1(new_n435), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n455), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n446), .A2(new_n410), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n453), .B1(new_n462), .B2(new_n424), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n443), .B(new_n292), .C1(new_n461), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT32), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n434), .A2(new_n424), .A3(new_n435), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT31), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n460), .A3(new_n454), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT32), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n443), .A4(new_n292), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n372), .B1(new_n452), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT9), .B(G234), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n314), .B1(new_n474), .B2(new_n292), .ZN(new_n475));
  INV_X1    g289(.A(G469), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n292), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n251), .A2(new_n210), .A3(new_n226), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT10), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n267), .B2(new_n198), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n272), .A2(KEYINPUT10), .A3(new_n396), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT78), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n399), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n478), .A2(new_n481), .A3(KEYINPUT78), .A4(new_n480), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n478), .A2(new_n481), .A3(new_n399), .A4(new_n480), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G110), .B(G140), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n212), .A2(G227), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n491), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT79), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n487), .A2(KEYINPUT79), .A3(new_n493), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n267), .A2(new_n198), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n244), .A2(new_n266), .B1(new_n195), .B2(new_n197), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n405), .B(KEYINPUT76), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT12), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(KEYINPUT77), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT77), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n405), .B(new_n503), .C1(new_n498), .C2(new_n499), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n501), .B1(new_n500), .B2(KEYINPUT77), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n496), .B(new_n497), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n492), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n477), .B1(new_n508), .B2(new_n476), .ZN(new_n509));
  INV_X1    g323(.A(new_n494), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n486), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n505), .A2(new_n506), .ZN(new_n512));
  INV_X1    g326(.A(new_n487), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(G469), .B(new_n511), .C1(new_n514), .C2(new_n493), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n475), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT15), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G478), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT93), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT92), .B1(new_n196), .B2(G143), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n191), .A3(G128), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n196), .A2(G143), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n376), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n376), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G122), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G116), .ZN(new_n530));
  INV_X1    g344(.A(G116), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G122), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n219), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n532), .A3(G107), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n530), .A2(KEYINPUT14), .A3(G107), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n530), .A2(new_n532), .A3(KEYINPUT14), .A4(G107), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n519), .B1(new_n528), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n527), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n525), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n542), .A2(KEYINPUT93), .A3(new_n537), .A4(new_n538), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n523), .A2(new_n545), .B1(new_n196), .B2(G143), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n545), .B2(new_n523), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G134), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n548), .A2(new_n525), .A3(new_n534), .A4(new_n535), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n473), .A2(new_n310), .A3(G953), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n544), .A2(new_n549), .A3(new_n551), .ZN(new_n554));
  AOI21_X1  g368(.A(G902), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT94), .ZN(new_n556));
  INV_X1    g370(.A(new_n554), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n551), .B1(new_n544), .B2(new_n549), .ZN(new_n558));
  OAI211_X1 g372(.A(KEYINPUT94), .B(new_n292), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n518), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G952), .ZN(new_n562));
  AOI211_X1 g376(.A(G953), .B(new_n562), .C1(G234), .C2(G237), .ZN(new_n563));
  OAI211_X1 g377(.A(G902), .B(G953), .C1(new_n315), .C2(new_n412), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n564), .B(KEYINPUT95), .Z(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT21), .B(G898), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n559), .A2(new_n517), .A3(G478), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n561), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT20), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n413), .A2(new_n415), .ZN(new_n572));
  NAND2_X1  g386(.A1(KEYINPUT85), .A2(G143), .ZN(new_n573));
  OAI21_X1  g387(.A(G214), .B1(KEYINPUT85), .B2(G143), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AND4_X1   g389(.A1(new_n212), .A2(new_n572), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n573), .B1(new_n416), .B2(new_n575), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT88), .B1(new_n578), .B2(G131), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n572), .A2(new_n212), .A3(new_n575), .ZN(new_n580));
  INV_X1    g394(.A(new_n573), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n416), .A2(new_n573), .A3(new_n575), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n582), .A2(KEYINPUT88), .A3(G131), .A4(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT17), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n328), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n582), .A2(G131), .A3(new_n583), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT88), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n582), .A2(new_n583), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n380), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n590), .A2(new_n592), .A3(new_n593), .A4(new_n584), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(new_n587), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n189), .B1(new_n322), .B2(new_n347), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n319), .A2(new_n189), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT87), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT87), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n348), .B2(new_n596), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT18), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n380), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n602), .B1(new_n591), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT86), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n578), .B2(new_n604), .ZN(new_n608));
  NOR4_X1   g422(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT86), .A4(new_n605), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(G113), .B(G122), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n217), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT90), .Z(new_n613));
  NAND3_X1  g427(.A1(new_n595), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n590), .A2(new_n584), .A3(new_n592), .ZN(new_n615));
  NOR2_X1   g429(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n617));
  MUX2_X1   g431(.A(new_n616), .B(new_n617), .S(new_n319), .Z(new_n618));
  AOI21_X1  g432(.A(new_n325), .B1(new_n618), .B2(new_n189), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n610), .ZN(new_n621));
  INV_X1    g435(.A(new_n612), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n614), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(G475), .A2(G902), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n571), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n625), .ZN(new_n627));
  AOI211_X1 g441(.A(KEYINPUT20), .B(new_n627), .C1(new_n614), .C2(new_n623), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n595), .A2(new_n610), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n622), .ZN(new_n630));
  AOI21_X1  g444(.A(G902), .B1(new_n630), .B2(new_n614), .ZN(new_n631));
  INV_X1    g445(.A(G475), .ZN(new_n632));
  OAI22_X1  g446(.A1(new_n626), .A2(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT91), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n612), .B1(new_n620), .B2(new_n610), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n605), .B1(new_n576), .B2(new_n577), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n601), .A3(new_n599), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n578), .A2(new_n607), .A3(new_n604), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT86), .B1(new_n591), .B2(new_n605), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n590), .A2(new_n584), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n328), .B1(new_n641), .B2(KEYINPUT17), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n640), .B1(new_n642), .B2(new_n594), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n635), .B1(new_n643), .B2(new_n613), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT20), .B1(new_n644), .B2(new_n627), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n624), .A2(new_n571), .A3(new_n625), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT91), .ZN(new_n648));
  INV_X1    g462(.A(new_n614), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n612), .B1(new_n595), .B2(new_n610), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n292), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(G475), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n647), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n570), .B1(new_n634), .B2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n309), .A2(new_n472), .A3(new_n516), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G101), .ZN(G3));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n513), .B1(new_n484), .B2(new_n485), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n507), .B1(new_n493), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n476), .A3(new_n292), .ZN(new_n660));
  INV_X1    g474(.A(new_n477), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n515), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n292), .B1(new_n461), .B2(new_n463), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(KEYINPUT96), .A3(G472), .ZN(new_n664));
  INV_X1    g478(.A(new_n475), .ZN(new_n665));
  NAND2_X1  g479(.A1(KEYINPUT96), .A2(G472), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n468), .A2(new_n292), .A3(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n662), .A2(new_n664), .A3(new_n665), .A4(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n657), .B1(new_n668), .B2(new_n372), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n664), .A2(new_n667), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(new_n516), .A3(KEYINPUT97), .A4(new_n371), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n557), .A2(new_n558), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT33), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n557), .A2(KEYINPUT33), .A3(new_n558), .ZN(new_n676));
  OAI211_X1 g490(.A(G478), .B(new_n292), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT98), .B(G478), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n678), .B1(new_n673), .B2(G902), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n634), .A2(new_n653), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n187), .B1(new_n298), .B2(new_n300), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n307), .B1(new_n303), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n567), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n672), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT34), .B(G104), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G6));
  XNOR2_X1  g502(.A(new_n567), .B(KEYINPUT99), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n307), .B(new_n689), .C1(new_n303), .C2(new_n683), .ZN(new_n690));
  INV_X1    g504(.A(new_n633), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n561), .A2(new_n569), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n672), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT100), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT35), .B(G107), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  NAND2_X1  g512(.A1(new_n357), .A2(new_n359), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n318), .A2(KEYINPUT36), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n369), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n365), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n668), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n309), .A3(new_n654), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT101), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n705), .B(new_n707), .ZN(G12));
  AOI21_X1  g522(.A(new_n703), .B1(new_n452), .B2(new_n471), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT102), .B(G900), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n563), .B1(new_n565), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT103), .B1(new_n693), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  INV_X1    g527(.A(new_n711), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n691), .A2(new_n713), .A3(new_n692), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n662), .A2(new_n665), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n684), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n709), .A2(new_n712), .A3(new_n715), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  AND3_X1   g533(.A1(new_n647), .A2(new_n648), .A3(new_n652), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n648), .B1(new_n647), .B2(new_n652), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n306), .B(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n308), .B1(new_n561), .B2(new_n569), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n722), .A2(new_n725), .A3(new_n703), .A4(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n711), .B(KEYINPUT39), .Z(new_n728));
  NAND2_X1  g542(.A1(new_n516), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(KEYINPUT40), .Z(new_n730));
  OAI21_X1  g544(.A(new_n455), .B1(new_n410), .B2(new_n407), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n466), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n292), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G472), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n471), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n727), .A2(new_n730), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G143), .ZN(G45));
  NAND4_X1  g551(.A1(new_n634), .A2(new_n680), .A3(new_n653), .A4(new_n714), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n709), .A2(new_n739), .A3(new_n717), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G146), .ZN(G48));
  NAND2_X1  g555(.A1(new_n659), .A2(new_n292), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n665), .A3(new_n660), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n472), .A2(new_n682), .A3(new_n685), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NAND3_X1  g562(.A1(new_n472), .A2(new_n694), .A3(new_n745), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT105), .B(G116), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G18));
  NOR2_X1   g565(.A1(new_n684), .A2(new_n744), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n709), .A2(new_n654), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  NAND2_X1  g568(.A1(new_n294), .A2(new_n301), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n634), .A2(new_n755), .A3(new_n726), .A4(new_n653), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n663), .A2(G472), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n371), .A2(new_n758), .A3(new_n464), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n743), .A2(new_n665), .A3(new_n660), .A4(new_n689), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NAND4_X1  g577(.A1(new_n722), .A2(KEYINPUT106), .A3(new_n680), .A4(new_n714), .ZN(new_n764));
  INV_X1    g578(.A(new_n703), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n765), .A2(new_n464), .A3(new_n758), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT106), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n738), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(new_n752), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  NAND2_X1  g584(.A1(new_n452), .A2(new_n471), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n308), .B1(new_n302), .B2(new_n305), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n771), .A2(new_n772), .A3(new_n371), .A4(new_n516), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n738), .B(KEYINPUT106), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(KEYINPUT42), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT42), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n764), .A2(new_n768), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n777), .B1(new_n778), .B2(new_n773), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  NAND2_X1  g595(.A1(new_n712), .A2(new_n715), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n773), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n376), .ZN(G36));
  INV_X1    g598(.A(new_n772), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n634), .A2(new_n653), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n680), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT43), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n670), .A2(new_n703), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n785), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n512), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n487), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n797), .A2(new_n491), .B1(new_n486), .B2(new_n510), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT45), .ZN(new_n799));
  OAI21_X1  g613(.A(G469), .B1(new_n798), .B2(KEYINPUT45), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n661), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n801), .A2(new_n802), .B1(new_n476), .B2(new_n508), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n665), .A3(new_n728), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT107), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n795), .B(new_n806), .C1(new_n794), .C2(new_n793), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G137), .ZN(G39));
  NAND2_X1  g622(.A1(new_n804), .A2(new_n665), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n665), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n785), .A2(new_n771), .A3(new_n738), .A4(new_n371), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g629(.A(KEYINPUT109), .B(G140), .Z(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(G42));
  NAND2_X1  g631(.A1(new_n772), .A2(new_n516), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n764), .A2(new_n766), .A3(new_n768), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n692), .A2(new_n633), .A3(new_n711), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n709), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n822), .A2(new_n823), .A3(new_n783), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n746), .A2(new_n749), .A3(new_n753), .A4(new_n762), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n779), .B2(new_n776), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n307), .A2(new_n302), .A3(new_n305), .A4(new_n689), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n681), .A2(KEYINPUT111), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT111), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n634), .A2(new_n680), .A3(new_n653), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n827), .A2(new_n828), .A3(KEYINPUT112), .A4(new_n830), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n672), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n655), .A2(new_n705), .ZN(new_n836));
  INV_X1    g650(.A(new_n827), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n786), .A2(new_n692), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n786), .A2(KEYINPUT113), .A3(new_n692), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n836), .B1(new_n842), .B2(new_n672), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n824), .A2(new_n826), .A3(new_n835), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n662), .A2(new_n703), .A3(new_n665), .A4(new_n714), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n465), .A2(new_n470), .B1(G472), .B2(new_n733), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n756), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n769), .A2(new_n718), .A3(new_n740), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n756), .A2(new_n845), .A3(new_n846), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n717), .A2(new_n771), .A3(new_n765), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n852), .B2(new_n739), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT52), .A3(new_n718), .A4(new_n769), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT114), .B1(new_n844), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n822), .A2(new_n783), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n826), .A2(new_n857), .A3(new_n835), .A4(new_n843), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n823), .B1(new_n858), .B2(new_n855), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n746), .A2(new_n749), .A3(new_n753), .A4(new_n762), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT42), .B1(new_n774), .B2(new_n775), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n778), .A2(new_n773), .A3(new_n777), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n840), .A2(new_n841), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n672), .A2(new_n827), .A3(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n655), .A2(new_n705), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n835), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n850), .A2(new_n854), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n824), .ZN(new_n871));
  XOR2_X1   g685(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n872));
  NAND4_X1  g686(.A1(new_n856), .A2(new_n859), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT53), .B1(new_n858), .B2(new_n855), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n868), .A2(new_n823), .A3(new_n870), .A4(new_n857), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT54), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n873), .A2(KEYINPUT116), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n772), .A2(new_n745), .ZN(new_n881));
  INV_X1    g695(.A(new_n563), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n881), .A2(new_n372), .A3(new_n882), .A4(new_n735), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT119), .ZN(new_n884));
  OAI211_X1 g698(.A(G952), .B(new_n212), .C1(new_n884), .C2(new_n681), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n788), .A2(new_n882), .A3(new_n759), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n752), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n887), .A2(KEYINPUT120), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT120), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n725), .A2(new_n307), .A3(new_n744), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT50), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n886), .A2(new_n892), .A3(KEYINPUT50), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n887), .A2(new_n785), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n743), .A2(new_n660), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n665), .B1(new_n899), .B2(KEYINPUT117), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(KEYINPUT117), .B2(new_n899), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n811), .A2(new_n812), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n883), .B(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n722), .A2(new_n680), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n788), .A2(new_n882), .A3(new_n881), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n905), .A2(new_n906), .B1(new_n766), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n897), .A2(new_n903), .A3(new_n908), .A4(KEYINPUT51), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n472), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT48), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n891), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n907), .A2(new_n766), .ZN(new_n913));
  INV_X1    g727(.A(new_n906), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n884), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n895), .B2(new_n896), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n901), .B(KEYINPUT118), .Z(new_n917));
  OAI21_X1  g731(.A(new_n898), .B1(new_n813), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT51), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n879), .A2(new_n880), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT121), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n879), .A2(new_n920), .A3(new_n923), .A4(new_n880), .ZN(new_n924));
  NOR2_X1   g738(.A1(G952), .A2(G953), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT122), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n899), .B(KEYINPUT49), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n371), .A2(new_n665), .A3(new_n307), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT110), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  OR4_X1    g745(.A1(new_n735), .A2(new_n725), .A3(new_n931), .A4(new_n787), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n927), .A2(new_n932), .ZN(G75));
  NOR2_X1   g747(.A1(new_n212), .A2(G952), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n856), .A2(new_n859), .A3(new_n871), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(G902), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT56), .B1(new_n938), .B2(G210), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n296), .A2(new_n297), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n295), .ZN(new_n941));
  XOR2_X1   g755(.A(KEYINPUT123), .B(KEYINPUT55), .Z(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT124), .Z(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n935), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n939), .B2(new_n945), .ZN(G51));
  INV_X1    g761(.A(new_n872), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n936), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n949), .A2(new_n873), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n477), .B(KEYINPUT57), .Z(new_n951));
  OAI21_X1  g765(.A(new_n659), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n937), .A2(new_n799), .A3(new_n800), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n934), .B1(new_n952), .B2(new_n953), .ZN(G54));
  INV_X1    g768(.A(KEYINPUT58), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n937), .A2(new_n955), .A3(new_n632), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n935), .B1(new_n956), .B2(new_n624), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n624), .B2(new_n956), .ZN(G60));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n675), .A2(new_n676), .ZN(new_n960));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT59), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n959), .B(new_n935), .C1(new_n950), .C2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n949), .B2(new_n873), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT125), .B1(new_n965), .B2(new_n934), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n879), .A2(new_n880), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n960), .B1(new_n968), .B2(new_n962), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT60), .Z(new_n972));
  NAND2_X1  g786(.A1(new_n936), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n934), .B1(new_n973), .B2(new_n367), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n701), .B2(new_n973), .ZN(new_n975));
  XNOR2_X1  g789(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G66));
  INV_X1    g792(.A(new_n566), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n212), .B1(new_n979), .B2(G224), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n867), .A2(new_n825), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT127), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n982), .B2(new_n212), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n940), .B1(G898), .B2(new_n212), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n983), .B(new_n984), .Z(G69));
  AND2_X1   g799(.A1(new_n769), .A2(new_n718), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n736), .A2(new_n740), .A3(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n828), .A2(new_n830), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n990), .A2(new_n840), .A3(new_n841), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n774), .A2(new_n728), .ZN(new_n992));
  AOI22_X1  g806(.A1(new_n813), .A2(new_n814), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n988), .A2(new_n807), .A3(new_n989), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n212), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n433), .B(new_n618), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(G900), .B2(G953), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n783), .B1(new_n776), .B2(new_n779), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n986), .A2(new_n740), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n472), .A2(new_n757), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n806), .B2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n807), .A2(new_n815), .A3(new_n1000), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n999), .B1(new_n1004), .B2(G953), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n212), .B1(G227), .B2(G900), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(G72));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  OAI21_X1  g824(.A(new_n1010), .B1(new_n994), .B2(new_n982), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(new_n424), .A3(new_n436), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1010), .B1(new_n1004), .B2(new_n982), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1013), .A2(new_n425), .A3(new_n462), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n466), .A2(new_n447), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n874), .A2(new_n875), .A3(new_n1010), .A4(new_n1015), .ZN(new_n1016));
  AND4_X1   g830(.A1(new_n935), .A2(new_n1012), .A3(new_n1014), .A4(new_n1016), .ZN(G57));
endmodule


