

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U324 ( .A(n571), .B(n295), .ZN(G1351GAT) );
  XNOR2_X1 U325 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n295) );
  NOR2_X1 U326 ( .A1(n300), .A2(n539), .ZN(n570) );
  XNOR2_X1 U327 ( .A(n439), .B(n292), .ZN(n300) );
  XNOR2_X1 U328 ( .A(n438), .B(n293), .ZN(n292) );
  INV_X1 U329 ( .A(KEYINPUT55), .ZN(n293) );
  XNOR2_X1 U330 ( .A(n347), .B(n297), .ZN(n296) );
  INV_X1 U331 ( .A(n348), .ZN(n297) );
  XNOR2_X1 U332 ( .A(n369), .B(n346), .ZN(n558) );
  XNOR2_X1 U333 ( .A(n294), .B(n334), .ZN(n345) );
  XNOR2_X1 U334 ( .A(n338), .B(n335), .ZN(n294) );
  NOR2_X1 U335 ( .A1(n296), .A2(n581), .ZN(n364) );
  XNOR2_X1 U336 ( .A(n419), .B(KEYINPUT65), .ZN(n573) );
  NOR2_X1 U337 ( .A1(n374), .A2(n373), .ZN(n377) );
  XOR2_X1 U338 ( .A(KEYINPUT74), .B(n565), .Z(n298) );
  XOR2_X1 U339 ( .A(KEYINPUT74), .B(n565), .Z(n569) );
  XNOR2_X1 U340 ( .A(n363), .B(n362), .ZN(n565) );
  XNOR2_X1 U341 ( .A(n351), .B(KEYINPUT11), .ZN(n352) );
  AND2_X1 U342 ( .A1(G230GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n375), .B(KEYINPUT115), .ZN(n376) );
  XNOR2_X1 U344 ( .A(n385), .B(n299), .ZN(n338) );
  XOR2_X1 U345 ( .A(G71GAT), .B(KEYINPUT13), .Z(n331) );
  XNOR2_X1 U346 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U347 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT47), .B(KEYINPUT113), .Z(n366) );
  XOR2_X1 U349 ( .A(G64GAT), .B(G57GAT), .Z(n302) );
  XNOR2_X1 U350 ( .A(G183GAT), .B(G127GAT), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U352 ( .A(KEYINPUT15), .B(KEYINPUT75), .Z(n304) );
  XNOR2_X1 U353 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U355 ( .A(n306), .B(n305), .ZN(n314) );
  XOR2_X1 U356 ( .A(G22GAT), .B(G155GAT), .Z(n425) );
  XNOR2_X1 U357 ( .A(G15GAT), .B(G1GAT), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n307), .B(G8GAT), .ZN(n326) );
  XOR2_X1 U359 ( .A(n425), .B(n326), .Z(n309) );
  NAND2_X1 U360 ( .A1(G231GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U362 ( .A(n331), .B(n310), .Z(n312) );
  XNOR2_X1 U363 ( .A(G211GAT), .B(G78GAT), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n581) );
  XNOR2_X1 U366 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n348) );
  XOR2_X1 U367 ( .A(G29GAT), .B(G43GAT), .Z(n316) );
  XNOR2_X1 U368 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n359) );
  XOR2_X1 U370 ( .A(n359), .B(KEYINPUT29), .Z(n318) );
  NAND2_X1 U371 ( .A1(G229GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U373 ( .A(KEYINPUT30), .B(G113GAT), .Z(n320) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(G197GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U376 ( .A(n322), .B(n321), .Z(n328) );
  XOR2_X1 U377 ( .A(G22GAT), .B(G141GAT), .Z(n324) );
  XNOR2_X1 U378 ( .A(G36GAT), .B(G50GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n575) );
  XOR2_X1 U382 ( .A(KEYINPUT69), .B(KEYINPUT71), .Z(n330) );
  XNOR2_X1 U383 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n329) );
  XOR2_X1 U384 ( .A(n330), .B(n329), .Z(n335) );
  XOR2_X1 U385 ( .A(KEYINPUT32), .B(n331), .Z(n333) );
  XOR2_X1 U386 ( .A(G120GAT), .B(G57GAT), .Z(n407) );
  XNOR2_X1 U387 ( .A(n407), .B(G92GAT), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U389 ( .A(G64GAT), .B(KEYINPUT70), .Z(n337) );
  XNOR2_X1 U390 ( .A(G176GAT), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n385) );
  XNOR2_X1 U392 ( .A(G78GAT), .B(KEYINPUT66), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n340), .B(G148GAT), .ZN(n431) );
  XOR2_X1 U394 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n342) );
  XNOR2_X1 U395 ( .A(G106GAT), .B(G85GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U397 ( .A(G99GAT), .B(n343), .Z(n363) );
  XNOR2_X1 U398 ( .A(n431), .B(n363), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n369) );
  XOR2_X1 U400 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n346) );
  NAND2_X1 U401 ( .A1(n575), .A2(n558), .ZN(n347) );
  XNOR2_X1 U402 ( .A(G36GAT), .B(G190GAT), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n350), .B(G92GAT), .ZN(n386) );
  AND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n386), .B(n352), .ZN(n356) );
  XOR2_X1 U406 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n354) );
  XNOR2_X1 U407 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U409 ( .A(n356), .B(n355), .Z(n361) );
  XOR2_X1 U410 ( .A(G162GAT), .B(KEYINPUT72), .Z(n358) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(G218GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n433) );
  XNOR2_X1 U413 ( .A(n359), .B(n433), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n362) );
  NAND2_X1 U415 ( .A1(n364), .A2(n565), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n366), .B(n365), .ZN(n374) );
  INV_X1 U417 ( .A(n581), .ZN(n494) );
  INV_X1 U418 ( .A(KEYINPUT36), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n367), .B(n569), .ZN(n492) );
  NOR2_X1 U420 ( .A1(n494), .A2(n492), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n368), .B(KEYINPUT45), .ZN(n371) );
  NOR2_X1 U422 ( .A1(n575), .A2(n369), .ZN(n370) );
  NAND2_X1 U423 ( .A1(n371), .A2(n370), .ZN(n372) );
  XOR2_X1 U424 ( .A(n372), .B(KEYINPUT114), .Z(n373) );
  INV_X1 U425 ( .A(KEYINPUT48), .ZN(n375) );
  XNOR2_X1 U426 ( .A(n377), .B(n376), .ZN(n536) );
  XOR2_X1 U427 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n379) );
  XNOR2_X1 U428 ( .A(KEYINPUT78), .B(KEYINPUT18), .ZN(n378) );
  XNOR2_X1 U429 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U430 ( .A(n380), .B(KEYINPUT77), .Z(n382) );
  XNOR2_X1 U431 ( .A(G169GAT), .B(G183GAT), .ZN(n381) );
  XNOR2_X1 U432 ( .A(n382), .B(n381), .ZN(n453) );
  XOR2_X1 U433 ( .A(G211GAT), .B(KEYINPUT83), .Z(n384) );
  XNOR2_X1 U434 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n383) );
  XNOR2_X1 U435 ( .A(n384), .B(n383), .ZN(n430) );
  XNOR2_X1 U436 ( .A(n430), .B(n385), .ZN(n393) );
  XOR2_X1 U437 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n391) );
  XOR2_X1 U438 ( .A(G218GAT), .B(G8GAT), .Z(n388) );
  NAND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U441 ( .A(n386), .B(n389), .ZN(n390) );
  XNOR2_X1 U442 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U443 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U444 ( .A(n453), .B(n394), .ZN(n526) );
  NOR2_X1 U445 ( .A1(n536), .A2(n526), .ZN(n395) );
  XNOR2_X1 U446 ( .A(n395), .B(KEYINPUT54), .ZN(n418) );
  XOR2_X1 U447 ( .A(KEYINPUT4), .B(KEYINPUT86), .Z(n397) );
  XNOR2_X1 U448 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n397), .B(n396), .ZN(n417) );
  XOR2_X1 U450 ( .A(KEYINPUT88), .B(G85GAT), .Z(n399) );
  XNOR2_X1 U451 ( .A(G148GAT), .B(G155GAT), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U453 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n401) );
  XNOR2_X1 U454 ( .A(KEYINPUT87), .B(KEYINPUT85), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U456 ( .A(n403), .B(n402), .Z(n415) );
  XNOR2_X1 U457 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n404), .B(KEYINPUT2), .ZN(n432) );
  XOR2_X1 U459 ( .A(n432), .B(G1GAT), .Z(n406) );
  NAND2_X1 U460 ( .A1(G225GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n413) );
  XOR2_X1 U462 ( .A(n407), .B(G162GAT), .Z(n411) );
  XOR2_X1 U463 ( .A(G127GAT), .B(KEYINPUT0), .Z(n409) );
  XNOR2_X1 U464 ( .A(G113GAT), .B(G134GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n441) );
  XNOR2_X1 U466 ( .A(G29GAT), .B(n441), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n524) );
  NAND2_X1 U471 ( .A1(n418), .A2(n524), .ZN(n419) );
  XOR2_X1 U472 ( .A(KEYINPUT24), .B(KEYINPUT82), .Z(n421) );
  XNOR2_X1 U473 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n420) );
  XNOR2_X1 U474 ( .A(n421), .B(n420), .ZN(n429) );
  XOR2_X1 U475 ( .A(KEYINPUT81), .B(G204GAT), .Z(n423) );
  XNOR2_X1 U476 ( .A(G106GAT), .B(KEYINPUT84), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U478 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n437) );
  XOR2_X1 U482 ( .A(n431), .B(n430), .Z(n435) );
  XNOR2_X1 U483 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U484 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U485 ( .A(n437), .B(n436), .ZN(n473) );
  NAND2_X1 U486 ( .A1(n573), .A2(n473), .ZN(n439) );
  XOR2_X1 U487 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n438) );
  XOR2_X1 U488 ( .A(G190GAT), .B(n441), .Z(n443) );
  XNOR2_X1 U489 ( .A(G43GAT), .B(KEYINPUT79), .ZN(n442) );
  XNOR2_X1 U490 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U491 ( .A(n444), .B(G99GAT), .Z(n449) );
  XOR2_X1 U492 ( .A(KEYINPUT76), .B(KEYINPUT20), .Z(n446) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U494 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U495 ( .A(G71GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U496 ( .A(n449), .B(n448), .ZN(n455) );
  XOR2_X1 U497 ( .A(G176GAT), .B(G120GAT), .Z(n451) );
  XNOR2_X1 U498 ( .A(G15GAT), .B(KEYINPUT80), .ZN(n450) );
  XNOR2_X1 U499 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U500 ( .A(n453), .B(n452), .Z(n454) );
  XNOR2_X1 U501 ( .A(n455), .B(n454), .ZN(n539) );
  NAND2_X1 U502 ( .A1(n570), .A2(n558), .ZN(n459) );
  XOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n457) );
  XNOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n456) );
  INV_X1 U505 ( .A(n575), .ZN(n510) );
  NOR2_X1 U506 ( .A1(n369), .A2(n510), .ZN(n498) );
  NOR2_X1 U507 ( .A1(n494), .A2(n298), .ZN(n460) );
  XNOR2_X1 U508 ( .A(n460), .B(KEYINPUT16), .ZN(n480) );
  INV_X1 U509 ( .A(n524), .ZN(n471) );
  NOR2_X1 U510 ( .A1(n539), .A2(n526), .ZN(n461) );
  XNOR2_X1 U511 ( .A(KEYINPUT95), .B(n461), .ZN(n462) );
  NAND2_X1 U512 ( .A1(n462), .A2(n473), .ZN(n463) );
  XNOR2_X1 U513 ( .A(n463), .B(KEYINPUT25), .ZN(n464) );
  XNOR2_X1 U514 ( .A(KEYINPUT96), .B(n464), .ZN(n469) );
  XNOR2_X1 U515 ( .A(KEYINPUT27), .B(n526), .ZN(n474) );
  XNOR2_X1 U516 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n467) );
  INV_X1 U517 ( .A(n539), .ZN(n465) );
  NOR2_X1 U518 ( .A1(n465), .A2(n473), .ZN(n466) );
  XNOR2_X1 U519 ( .A(n467), .B(n466), .ZN(n574) );
  INV_X1 U520 ( .A(n574), .ZN(n554) );
  NOR2_X1 U521 ( .A1(n474), .A2(n554), .ZN(n468) );
  NOR2_X1 U522 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U523 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U524 ( .A(KEYINPUT97), .B(n472), .ZN(n479) );
  XOR2_X1 U525 ( .A(n473), .B(KEYINPUT28), .Z(n542) );
  NOR2_X1 U526 ( .A1(n474), .A2(n524), .ZN(n475) );
  XOR2_X1 U527 ( .A(KEYINPUT92), .B(n475), .Z(n537) );
  NOR2_X1 U528 ( .A1(n542), .A2(n537), .ZN(n476) );
  NAND2_X1 U529 ( .A1(n476), .A2(n539), .ZN(n477) );
  XOR2_X1 U530 ( .A(KEYINPUT93), .B(n477), .Z(n478) );
  NAND2_X1 U531 ( .A1(n479), .A2(n478), .ZN(n493) );
  NAND2_X1 U532 ( .A1(n480), .A2(n493), .ZN(n481) );
  XOR2_X1 U533 ( .A(KEYINPUT98), .B(n481), .Z(n511) );
  NAND2_X1 U534 ( .A1(n498), .A2(n511), .ZN(n490) );
  NOR2_X1 U535 ( .A1(n524), .A2(n490), .ZN(n483) );
  XNOR2_X1 U536 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n482) );
  XNOR2_X1 U537 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NOR2_X1 U539 ( .A1(n526), .A2(n490), .ZN(n485) );
  XOR2_X1 U540 ( .A(KEYINPUT100), .B(n485), .Z(n486) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U542 ( .A1(n539), .A2(n490), .ZN(n488) );
  XNOR2_X1 U543 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U544 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U545 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  INV_X1 U546 ( .A(n542), .ZN(n532) );
  NOR2_X1 U547 ( .A1(n532), .A2(n490), .ZN(n491) );
  XOR2_X1 U548 ( .A(G22GAT), .B(n491), .Z(G1327GAT) );
  XNOR2_X1 U549 ( .A(KEYINPUT103), .B(KEYINPUT38), .ZN(n500) );
  NAND2_X1 U550 ( .A1(n494), .A2(n493), .ZN(n495) );
  NOR2_X1 U551 ( .A1(n492), .A2(n495), .ZN(n497) );
  XOR2_X1 U552 ( .A(KEYINPUT37), .B(KEYINPUT102), .Z(n496) );
  XNOR2_X1 U553 ( .A(n497), .B(n496), .ZN(n522) );
  NAND2_X1 U554 ( .A1(n522), .A2(n498), .ZN(n499) );
  XOR2_X1 U555 ( .A(n500), .B(n499), .Z(n507) );
  NOR2_X1 U556 ( .A1(n507), .A2(n524), .ZN(n501) );
  XNOR2_X1 U557 ( .A(n501), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n507), .A2(n526), .ZN(n503) );
  XOR2_X1 U560 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  NOR2_X1 U561 ( .A1(n507), .A2(n539), .ZN(n505) );
  XNOR2_X1 U562 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U564 ( .A(G43GAT), .B(n506), .Z(G1330GAT) );
  NOR2_X1 U565 ( .A1(n507), .A2(n532), .ZN(n509) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n508) );
  XNOR2_X1 U567 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  XNOR2_X1 U568 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n515) );
  AND2_X1 U569 ( .A1(n510), .A2(n558), .ZN(n523) );
  NAND2_X1 U570 ( .A1(n523), .A2(n511), .ZN(n519) );
  NOR2_X1 U571 ( .A1(n524), .A2(n519), .ZN(n513) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n512) );
  XNOR2_X1 U573 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U574 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n526), .A2(n519), .ZN(n516) );
  XOR2_X1 U576 ( .A(KEYINPUT108), .B(n516), .Z(n517) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n517), .ZN(G1333GAT) );
  NOR2_X1 U578 ( .A1(n539), .A2(n519), .ZN(n518) );
  XOR2_X1 U579 ( .A(G71GAT), .B(n518), .Z(G1334GAT) );
  NOR2_X1 U580 ( .A1(n532), .A2(n519), .ZN(n521) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n520) );
  XNOR2_X1 U582 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n523), .A2(n522), .ZN(n531) );
  NOR2_X1 U584 ( .A1(n524), .A2(n531), .ZN(n525) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n525), .Z(G1336GAT) );
  NOR2_X1 U586 ( .A1(n526), .A2(n531), .ZN(n528) );
  XNOR2_X1 U587 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n527) );
  XNOR2_X1 U588 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NOR2_X1 U590 ( .A1(n539), .A2(n531), .ZN(n530) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n530), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U593 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U594 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U597 ( .A(KEYINPUT116), .B(n538), .Z(n555) );
  NOR2_X1 U598 ( .A1(n555), .A2(n539), .ZN(n540) );
  XNOR2_X1 U599 ( .A(n540), .B(KEYINPUT117), .ZN(n541) );
  NOR2_X1 U600 ( .A1(n542), .A2(n541), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n551), .A2(n575), .ZN(n543) );
  XNOR2_X1 U602 ( .A(n543), .B(KEYINPUT118), .ZN(n544) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n544), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT120), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U605 ( .A1(n551), .A2(n558), .ZN(n545) );
  XNOR2_X1 U606 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT119), .Z(n547) );
  XNOR2_X1 U608 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  NAND2_X1 U609 ( .A1(n551), .A2(n581), .ZN(n549) );
  XNOR2_X1 U610 ( .A(n549), .B(KEYINPUT50), .ZN(n550) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U613 ( .A1(n551), .A2(n298), .ZN(n552) );
  XNOR2_X1 U614 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NOR2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U616 ( .A(KEYINPUT121), .B(n556), .Z(n563) );
  NAND2_X1 U617 ( .A1(n563), .A2(n575), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n557), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n560) );
  NAND2_X1 U620 ( .A1(n563), .A2(n558), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n563), .A2(n581), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n562), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U625 ( .A(n563), .ZN(n564) );
  NOR2_X1 U626 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n566), .Z(G1347GAT) );
  NAND2_X1 U628 ( .A1(n570), .A2(n575), .ZN(n567) );
  XNOR2_X1 U629 ( .A(n567), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n570), .A2(n581), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n570), .A2(n298), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n577) );
  NAND2_X1 U634 ( .A1(n573), .A2(n574), .ZN(n587) );
  INV_X1 U635 ( .A(n587), .ZN(n582) );
  NAND2_X1 U636 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U637 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U640 ( .A1(n582), .A2(n369), .ZN(n579) );
  XNOR2_X1 U641 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT125), .Z(n584) );
  NAND2_X1 U643 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U644 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n586) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U647 ( .A(n586), .B(n585), .ZN(n589) );
  NOR2_X1 U648 ( .A1(n492), .A2(n587), .ZN(n588) );
  XOR2_X1 U649 ( .A(n589), .B(n588), .Z(G1355GAT) );
endmodule

