

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773;

  NAND2_X1 U374 ( .A1(n354), .A2(n643), .ZN(n644) );
  INV_X1 U375 ( .A(n641), .ZN(n355) );
  NOR2_X1 U376 ( .A1(n742), .A2(n765), .ZN(n686) );
  AND2_X1 U377 ( .A1(n650), .A2(KEYINPUT86), .ZN(n598) );
  AND2_X1 U378 ( .A1(n587), .A2(n698), .ZN(n616) );
  INV_X1 U379 ( .A(n535), .ZN(n681) );
  XNOR2_X1 U380 ( .A(n463), .B(n462), .ZN(n582) );
  OR2_X1 U381 ( .A1(n737), .A2(G902), .ZN(n497) );
  XNOR2_X2 U382 ( .A(n642), .B(n355), .ZN(n354) );
  INV_X2 U383 ( .A(G953), .ZN(n766) );
  NOR2_X2 U384 ( .A1(n659), .A2(n741), .ZN(n660) );
  INV_X2 U385 ( .A(n742), .ZN(n385) );
  XNOR2_X2 U386 ( .A(n628), .B(n627), .ZN(n742) );
  XNOR2_X2 U387 ( .A(n441), .B(KEYINPUT4), .ZN(n482) );
  NAND2_X1 U388 ( .A1(n770), .A2(n646), .ZN(n538) );
  XNOR2_X2 U389 ( .A(n635), .B(KEYINPUT65), .ZN(n661) );
  NOR2_X1 U390 ( .A1(n765), .A2(n391), .ZN(n384) );
  NAND2_X1 U391 ( .A1(n367), .A2(n362), .ZN(n765) );
  OR2_X1 U392 ( .A1(n640), .A2(G902), .ZN(n417) );
  XNOR2_X1 U393 ( .A(G116), .B(G113), .ZN(n412) );
  XNOR2_X1 U394 ( .A(G101), .B(KEYINPUT74), .ZN(n411) );
  XNOR2_X2 U395 ( .A(n635), .B(KEYINPUT65), .ZN(n356) );
  NAND2_X2 U396 ( .A1(n388), .A2(n690), .ZN(n635) );
  XNOR2_X2 U397 ( .A(n597), .B(n596), .ZN(n650) );
  XNOR2_X1 U398 ( .A(n546), .B(KEYINPUT38), .ZN(n708) );
  XNOR2_X1 U399 ( .A(n528), .B(n527), .ZN(n565) );
  AND2_X1 U400 ( .A1(n539), .A2(n540), .ZN(n368) );
  INV_X1 U401 ( .A(n395), .ZN(n391) );
  NOR2_X1 U402 ( .A1(G237), .A2(G902), .ZN(n485) );
  NOR2_X1 U403 ( .A1(n618), .A2(n398), .ZN(n397) );
  NAND2_X1 U404 ( .A1(n708), .A2(n399), .ZN(n398) );
  INV_X1 U405 ( .A(G902), .ZN(n550) );
  XNOR2_X1 U406 ( .A(n368), .B(n541), .ZN(n367) );
  INV_X1 U407 ( .A(KEYINPUT71), .ZN(n405) );
  INV_X1 U408 ( .A(G122), .ZN(n425) );
  XNOR2_X1 U409 ( .A(G140), .B(G143), .ZN(n421) );
  XOR2_X1 U410 ( .A(KEYINPUT99), .B(G113), .Z(n422) );
  XNOR2_X1 U411 ( .A(G101), .B(G104), .ZN(n492) );
  XNOR2_X1 U412 ( .A(G146), .B(G125), .ZN(n479) );
  NAND2_X1 U413 ( .A1(n376), .A2(n373), .ZN(n727) );
  NAND2_X1 U414 ( .A1(n375), .A2(n374), .ZN(n373) );
  NOR2_X1 U415 ( .A1(n711), .A2(n379), .ZN(n374) );
  XNOR2_X1 U416 ( .A(n488), .B(n364), .ZN(n561) );
  NOR2_X1 U417 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U418 ( .A(n524), .B(KEYINPUT110), .ZN(n712) );
  NOR2_X1 U419 ( .A1(G953), .A2(G237), .ZN(n418) );
  INV_X1 U420 ( .A(G128), .ZN(n403) );
  NOR2_X1 U421 ( .A1(n765), .A2(n366), .ZN(n389) );
  NAND2_X1 U422 ( .A1(n395), .A2(n392), .ZN(n390) );
  INV_X1 U423 ( .A(KEYINPUT41), .ZN(n379) );
  NAND2_X1 U424 ( .A1(n711), .A2(n379), .ZN(n377) );
  XNOR2_X1 U425 ( .A(n448), .B(n447), .ZN(n526) );
  XNOR2_X1 U426 ( .A(KEYINPUT3), .B(G119), .ZN(n413) );
  XNOR2_X1 U427 ( .A(G128), .B(G110), .ZN(n455) );
  XNOR2_X1 U428 ( .A(G134), .B(G107), .ZN(n438) );
  INV_X1 U429 ( .A(KEYINPUT101), .ZN(n437) );
  XNOR2_X1 U430 ( .A(G116), .B(G122), .ZN(n435) );
  XNOR2_X1 U431 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n478) );
  XNOR2_X1 U432 ( .A(n400), .B(n534), .ZN(n549) );
  XNOR2_X1 U433 ( .A(n394), .B(KEYINPUT97), .ZN(n704) );
  AND2_X1 U434 ( .A1(n695), .A2(n698), .ZN(n393) );
  NAND2_X2 U435 ( .A1(n370), .A2(n369), .ZN(n546) );
  OR2_X1 U436 ( .A1(n663), .A2(n360), .ZN(n369) );
  NAND2_X1 U437 ( .A1(n486), .A2(n633), .ZN(n371) );
  BUF_X1 U438 ( .A(n579), .Z(n695) );
  NAND2_X1 U439 ( .A1(n561), .A2(n560), .ZN(n563) );
  AND2_X1 U440 ( .A1(n578), .A2(n577), .ZN(n606) );
  XNOR2_X1 U441 ( .A(n430), .B(n429), .ZN(n656) );
  XNOR2_X1 U442 ( .A(n428), .B(n460), .ZN(n429) );
  BUF_X1 U443 ( .A(n356), .Z(n734) );
  XNOR2_X1 U444 ( .A(n387), .B(n496), .ZN(n737) );
  NOR2_X1 U445 ( .A1(n727), .A2(n529), .ZN(n531) );
  XNOR2_X1 U446 ( .A(n536), .B(KEYINPUT40), .ZN(n646) );
  OR2_X1 U447 ( .A1(n549), .A2(n535), .ZN(n536) );
  XNOR2_X1 U448 ( .A(n386), .B(n581), .ZN(n583) );
  XOR2_X1 U449 ( .A(n426), .B(G134), .Z(n357) );
  XOR2_X1 U450 ( .A(n455), .B(KEYINPUT89), .Z(n358) );
  XOR2_X1 U451 ( .A(KEYINPUT23), .B(KEYINPUT75), .Z(n359) );
  OR2_X1 U452 ( .A1(n486), .A2(n633), .ZN(n360) );
  AND2_X1 U453 ( .A1(n648), .A2(n645), .ZN(n362) );
  AND2_X1 U454 ( .A1(n577), .A2(n580), .ZN(n363) );
  XOR2_X1 U455 ( .A(KEYINPUT68), .B(KEYINPUT19), .Z(n364) );
  NOR2_X1 U456 ( .A1(n401), .A2(n634), .ZN(n365) );
  XNOR2_X1 U457 ( .A(KEYINPUT15), .B(G902), .ZN(n484) );
  NAND2_X1 U458 ( .A1(n392), .A2(n633), .ZN(n366) );
  AND2_X1 U459 ( .A1(n372), .A2(n371), .ZN(n370) );
  NAND2_X1 U460 ( .A1(n663), .A2(n486), .ZN(n372) );
  XNOR2_X1 U461 ( .A(n483), .B(n751), .ZN(n663) );
  NAND2_X1 U462 ( .A1(n712), .A2(n379), .ZN(n378) );
  INV_X1 U463 ( .A(n712), .ZN(n375) );
  AND2_X1 U464 ( .A1(n378), .A2(n377), .ZN(n376) );
  INV_X1 U465 ( .A(n380), .ZN(n586) );
  NAND2_X1 U466 ( .A1(n649), .A2(n584), .ZN(n380) );
  NAND2_X1 U467 ( .A1(n380), .A2(n604), .ZN(n615) );
  NAND2_X1 U468 ( .A1(n382), .A2(n381), .ZN(n388) );
  NAND2_X1 U469 ( .A1(n389), .A2(n385), .ZN(n381) );
  NAND2_X1 U470 ( .A1(n383), .A2(n390), .ZN(n382) );
  NAND2_X1 U471 ( .A1(n385), .A2(n384), .ZN(n383) );
  NOR2_X2 U472 ( .A1(n546), .A2(n511), .ZN(n488) );
  NAND2_X1 U473 ( .A1(n578), .A2(n363), .ZN(n386) );
  XNOR2_X2 U474 ( .A(n569), .B(n568), .ZN(n578) );
  XNOR2_X1 U475 ( .A(n387), .B(n416), .ZN(n640) );
  XNOR2_X2 U476 ( .A(n758), .B(G146), .ZN(n387) );
  NAND2_X1 U477 ( .A1(n686), .A2(KEYINPUT2), .ZN(n690) );
  INV_X1 U478 ( .A(KEYINPUT81), .ZN(n392) );
  NAND2_X1 U479 ( .A1(n393), .A2(n587), .ZN(n394) );
  NAND2_X1 U480 ( .A1(n704), .A2(n590), .ZN(n617) );
  NOR2_X1 U481 ( .A1(n365), .A2(n631), .ZN(n395) );
  NOR2_X1 U482 ( .A1(n618), .A2(n516), .ZN(n396) );
  AND2_X1 U483 ( .A1(n517), .A2(n396), .ZN(n532) );
  NAND2_X1 U484 ( .A1(n517), .A2(n397), .ZN(n400) );
  INV_X1 U485 ( .A(n516), .ZN(n399) );
  XNOR2_X1 U486 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X1 U487 ( .A1(KEYINPUT81), .A2(KEYINPUT67), .ZN(n401) );
  AND2_X1 U488 ( .A1(n639), .A2(n643), .ZN(G63) );
  OR2_X1 U489 ( .A1(n522), .A2(n678), .ZN(n523) );
  INV_X1 U490 ( .A(KEYINPUT102), .ZN(n527) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n446) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n525) );
  INV_X1 U495 ( .A(n741), .ZN(n643) );
  XNOR2_X2 U496 ( .A(G143), .B(KEYINPUT64), .ZN(n404) );
  XNOR2_X2 U497 ( .A(n404), .B(n403), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n405), .B(G131), .ZN(n426) );
  XNOR2_X2 U499 ( .A(n482), .B(n357), .ZN(n758) );
  XOR2_X1 U500 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n407) );
  NAND2_X1 U501 ( .A1(n418), .A2(G210), .ZN(n406) );
  XNOR2_X1 U502 ( .A(n407), .B(n406), .ZN(n410) );
  XNOR2_X1 U503 ( .A(KEYINPUT96), .B(KEYINPUT5), .ZN(n408) );
  XNOR2_X1 U504 ( .A(n408), .B(G137), .ZN(n409) );
  XNOR2_X1 U505 ( .A(n410), .B(n409), .ZN(n415) );
  XNOR2_X1 U506 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X1 U507 ( .A(n414), .B(n413), .ZN(n476) );
  XNOR2_X1 U508 ( .A(n415), .B(n476), .ZN(n416) );
  XNOR2_X2 U509 ( .A(n417), .B(G472), .ZN(n579) );
  XNOR2_X1 U510 ( .A(n579), .B(KEYINPUT6), .ZN(n605) );
  XOR2_X1 U511 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n420) );
  NAND2_X1 U512 ( .A1(n418), .A2(G214), .ZN(n419) );
  XNOR2_X1 U513 ( .A(n420), .B(n419), .ZN(n424) );
  XNOR2_X1 U514 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U515 ( .A(n424), .B(n423), .Z(n430) );
  XNOR2_X1 U516 ( .A(n425), .B(G104), .ZN(n474) );
  XNOR2_X1 U517 ( .A(n426), .B(n474), .ZN(n428) );
  XNOR2_X1 U518 ( .A(KEYINPUT10), .B(KEYINPUT70), .ZN(n427) );
  XNOR2_X1 U519 ( .A(n427), .B(n479), .ZN(n460) );
  NOR2_X1 U520 ( .A1(G902), .A2(n656), .ZN(n434) );
  XNOR2_X1 U521 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n432) );
  INV_X1 U522 ( .A(G475), .ZN(n431) );
  XOR2_X1 U523 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n436) );
  XNOR2_X1 U524 ( .A(n436), .B(n435), .ZN(n440) );
  INV_X1 U525 ( .A(n441), .ZN(n444) );
  NAND2_X1 U526 ( .A1(G234), .A2(n766), .ZN(n442) );
  XOR2_X1 U527 ( .A(KEYINPUT8), .B(n442), .Z(n454) );
  NAND2_X1 U528 ( .A1(G217), .A2(n454), .ZN(n443) );
  XNOR2_X1 U529 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U530 ( .A(n446), .B(n445), .ZN(n636) );
  NAND2_X1 U531 ( .A1(n636), .A2(n550), .ZN(n448) );
  INV_X1 U532 ( .A(G478), .ZN(n447) );
  INV_X1 U533 ( .A(n526), .ZN(n508) );
  OR2_X1 U534 ( .A1(n525), .A2(n508), .ZN(n535) );
  XOR2_X1 U535 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n452) );
  NAND2_X1 U536 ( .A1(n484), .A2(G234), .ZN(n449) );
  XNOR2_X1 U537 ( .A(n449), .B(KEYINPUT20), .ZN(n450) );
  XNOR2_X1 U538 ( .A(KEYINPUT90), .B(n450), .ZN(n464) );
  NAND2_X1 U539 ( .A1(G217), .A2(n464), .ZN(n451) );
  XNOR2_X1 U540 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U541 ( .A(n453), .B(KEYINPUT91), .ZN(n463) );
  NAND2_X1 U542 ( .A1(G221), .A2(n454), .ZN(n459) );
  XNOR2_X1 U543 ( .A(G119), .B(KEYINPUT24), .ZN(n456) );
  XNOR2_X1 U544 ( .A(n359), .B(n456), .ZN(n457) );
  XNOR2_X1 U545 ( .A(n358), .B(n457), .ZN(n458) );
  XNOR2_X1 U546 ( .A(n459), .B(n458), .ZN(n461) );
  XOR2_X1 U547 ( .A(G137), .B(G140), .Z(n490) );
  XNOR2_X1 U548 ( .A(n490), .B(n460), .ZN(n757) );
  XNOR2_X1 U549 ( .A(n461), .B(n757), .ZN(n651) );
  NAND2_X1 U550 ( .A1(n651), .A2(n550), .ZN(n462) );
  NAND2_X1 U551 ( .A1(n464), .A2(G221), .ZN(n465) );
  XNOR2_X1 U552 ( .A(n465), .B(KEYINPUT21), .ZN(n691) );
  NAND2_X1 U553 ( .A1(G237), .A2(G234), .ZN(n466) );
  XNOR2_X1 U554 ( .A(n466), .B(KEYINPUT14), .ZN(n723) );
  NOR2_X1 U555 ( .A1(G900), .A2(n766), .ZN(n467) );
  NAND2_X1 U556 ( .A1(n467), .A2(G902), .ZN(n468) );
  NAND2_X1 U557 ( .A1(G952), .A2(n766), .ZN(n555) );
  NAND2_X1 U558 ( .A1(n468), .A2(n555), .ZN(n469) );
  NAND2_X1 U559 ( .A1(n723), .A2(n469), .ZN(n516) );
  NOR2_X1 U560 ( .A1(n691), .A2(n516), .ZN(n470) );
  XOR2_X1 U561 ( .A(n470), .B(KEYINPUT73), .Z(n471) );
  AND2_X1 U562 ( .A1(n582), .A2(n471), .ZN(n502) );
  NAND2_X1 U563 ( .A1(n681), .A2(n502), .ZN(n472) );
  NOR2_X1 U564 ( .A1(n605), .A2(n472), .ZN(n473) );
  XNOR2_X1 U565 ( .A(n473), .B(KEYINPUT106), .ZN(n542) );
  XNOR2_X2 U566 ( .A(G110), .B(G107), .ZN(n493) );
  XNOR2_X1 U567 ( .A(n493), .B(KEYINPUT16), .ZN(n475) );
  XNOR2_X1 U568 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X1 U569 ( .A(n477), .B(n476), .ZN(n751) );
  NAND2_X1 U570 ( .A1(n766), .A2(G224), .ZN(n745) );
  XNOR2_X1 U571 ( .A(n478), .B(n745), .ZN(n480) );
  XNOR2_X1 U572 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U573 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U574 ( .A(n484), .ZN(n633) );
  XNOR2_X1 U575 ( .A(n485), .B(KEYINPUT79), .ZN(n487) );
  NAND2_X1 U576 ( .A1(n487), .A2(G210), .ZN(n486) );
  AND2_X1 U577 ( .A1(n487), .A2(G214), .ZN(n511) );
  AND2_X1 U578 ( .A1(n542), .A2(n488), .ZN(n489) );
  XNOR2_X1 U579 ( .A(n489), .B(KEYINPUT36), .ZN(n499) );
  NAND2_X1 U580 ( .A1(n766), .A2(G227), .ZN(n491) );
  XNOR2_X1 U581 ( .A(n491), .B(n490), .ZN(n495) );
  XNOR2_X1 U582 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U583 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X2 U584 ( .A(n497), .B(G469), .ZN(n504) );
  XNOR2_X2 U585 ( .A(n504), .B(KEYINPUT1), .ZN(n587) );
  XNOR2_X1 U586 ( .A(n587), .B(KEYINPUT87), .ZN(n571) );
  INV_X1 U587 ( .A(n571), .ZN(n498) );
  NAND2_X1 U588 ( .A1(n499), .A2(n498), .ZN(n501) );
  INV_X1 U589 ( .A(KEYINPUT112), .ZN(n500) );
  XNOR2_X1 U590 ( .A(n501), .B(n500), .ZN(n772) );
  NAND2_X1 U591 ( .A1(n579), .A2(n502), .ZN(n503) );
  XNOR2_X1 U592 ( .A(n503), .B(KEYINPUT28), .ZN(n506) );
  INV_X1 U593 ( .A(n504), .ZN(n505) );
  OR2_X1 U594 ( .A1(n506), .A2(n505), .ZN(n529) );
  INV_X1 U595 ( .A(n561), .ZN(n507) );
  NOR2_X2 U596 ( .A1(n529), .A2(n507), .ZN(n679) );
  AND2_X1 U597 ( .A1(n525), .A2(n508), .ZN(n683) );
  INV_X1 U598 ( .A(n683), .ZN(n548) );
  AND2_X1 U599 ( .A1(n548), .A2(n535), .ZN(n713) );
  NOR2_X1 U600 ( .A1(n713), .A2(KEYINPUT69), .ZN(n509) );
  NAND2_X1 U601 ( .A1(n679), .A2(n509), .ZN(n510) );
  XNOR2_X1 U602 ( .A(n510), .B(KEYINPUT47), .ZN(n522) );
  INV_X1 U603 ( .A(n511), .ZN(n707) );
  NAND2_X1 U604 ( .A1(n579), .A2(n707), .ZN(n514) );
  INV_X1 U605 ( .A(KEYINPUT108), .ZN(n512) );
  XNOR2_X1 U606 ( .A(n512), .B(KEYINPUT30), .ZN(n513) );
  XNOR2_X1 U607 ( .A(n514), .B(n513), .ZN(n517) );
  INV_X1 U608 ( .A(n582), .ZN(n515) );
  XNOR2_X1 U609 ( .A(n691), .B(KEYINPUT93), .ZN(n564) );
  AND2_X1 U610 ( .A1(n515), .A2(n564), .ZN(n698) );
  NAND2_X1 U611 ( .A1(n504), .A2(n698), .ZN(n618) );
  INV_X1 U612 ( .A(n546), .ZN(n518) );
  NAND2_X1 U613 ( .A1(n532), .A2(n518), .ZN(n519) );
  XNOR2_X1 U614 ( .A(n519), .B(KEYINPUT109), .ZN(n521) );
  OR2_X1 U615 ( .A1(n525), .A2(n526), .ZN(n520) );
  XNOR2_X1 U616 ( .A(n520), .B(KEYINPUT105), .ZN(n593) );
  AND2_X1 U617 ( .A1(n521), .A2(n593), .ZN(n678) );
  NOR2_X1 U618 ( .A1(n772), .A2(n523), .ZN(n540) );
  NAND2_X1 U619 ( .A1(n708), .A2(n707), .ZN(n524) );
  NAND2_X1 U620 ( .A1(n526), .A2(n525), .ZN(n528) );
  INV_X1 U621 ( .A(n565), .ZN(n711) );
  XNOR2_X1 U622 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n530) );
  XNOR2_X1 U623 ( .A(n531), .B(n530), .ZN(n770) );
  XNOR2_X1 U624 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n533) );
  XNOR2_X1 U625 ( .A(n533), .B(KEYINPUT77), .ZN(n534) );
  XNOR2_X1 U626 ( .A(KEYINPUT83), .B(KEYINPUT46), .ZN(n537) );
  XNOR2_X1 U627 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U628 ( .A(KEYINPUT72), .B(KEYINPUT48), .ZN(n541) );
  NAND2_X1 U629 ( .A1(n542), .A2(n707), .ZN(n543) );
  XNOR2_X1 U630 ( .A(KEYINPUT107), .B(n543), .ZN(n544) );
  INV_X1 U631 ( .A(n587), .ZN(n577) );
  NAND2_X1 U632 ( .A1(n544), .A2(n577), .ZN(n545) );
  XNOR2_X1 U633 ( .A(n545), .B(KEYINPUT43), .ZN(n547) );
  NAND2_X1 U634 ( .A1(n547), .A2(n546), .ZN(n648) );
  OR2_X1 U635 ( .A1(n549), .A2(n548), .ZN(n645) );
  INV_X1 U636 ( .A(G898), .ZN(n748) );
  NAND2_X1 U637 ( .A1(G953), .A2(n748), .ZN(n752) );
  OR2_X1 U638 ( .A1(n550), .A2(n752), .ZN(n552) );
  NOR2_X1 U639 ( .A1(KEYINPUT88), .A2(n552), .ZN(n551) );
  NAND2_X1 U640 ( .A1(n723), .A2(n551), .ZN(n554) );
  NAND2_X1 U641 ( .A1(KEYINPUT88), .A2(n552), .ZN(n553) );
  NAND2_X1 U642 ( .A1(n554), .A2(n553), .ZN(n556) );
  NAND2_X1 U643 ( .A1(n556), .A2(n555), .ZN(n559) );
  INV_X1 U644 ( .A(KEYINPUT88), .ZN(n557) );
  OR2_X1 U645 ( .A1(n723), .A2(n557), .ZN(n558) );
  AND2_X1 U646 ( .A1(n559), .A2(n558), .ZN(n560) );
  INV_X1 U647 ( .A(KEYINPUT0), .ZN(n562) );
  XNOR2_X2 U648 ( .A(n563), .B(n562), .ZN(n590) );
  NAND2_X1 U649 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U650 ( .A(n566), .B(KEYINPUT103), .ZN(n567) );
  NAND2_X1 U651 ( .A1(n590), .A2(n567), .ZN(n569) );
  INV_X1 U652 ( .A(KEYINPUT22), .ZN(n568) );
  XNOR2_X1 U653 ( .A(n582), .B(KEYINPUT104), .ZN(n692) );
  NAND2_X1 U654 ( .A1(n605), .A2(n692), .ZN(n570) );
  OR2_X1 U655 ( .A1(n571), .A2(n570), .ZN(n573) );
  INV_X1 U656 ( .A(KEYINPUT80), .ZN(n572) );
  XNOR2_X1 U657 ( .A(n573), .B(n572), .ZN(n574) );
  NAND2_X1 U658 ( .A1(n578), .A2(n574), .ZN(n576) );
  INV_X1 U659 ( .A(KEYINPUT32), .ZN(n575) );
  XNOR2_X1 U660 ( .A(n576), .B(n575), .ZN(n771) );
  INV_X1 U661 ( .A(n771), .ZN(n584) );
  INV_X1 U662 ( .A(n695), .ZN(n580) );
  INV_X1 U663 ( .A(KEYINPUT66), .ZN(n581) );
  NAND2_X1 U664 ( .A1(n583), .A2(n582), .ZN(n649) );
  INV_X1 U665 ( .A(KEYINPUT44), .ZN(n610) );
  NAND2_X1 U666 ( .A1(n610), .A2(KEYINPUT76), .ZN(n604) );
  INV_X1 U667 ( .A(n604), .ZN(n585) );
  NAND2_X1 U668 ( .A1(n586), .A2(n585), .ZN(n599) );
  INV_X1 U669 ( .A(n605), .ZN(n588) );
  NAND2_X1 U670 ( .A1(n616), .A2(n588), .ZN(n589) );
  XNOR2_X2 U671 ( .A(n589), .B(KEYINPUT33), .ZN(n716) );
  NAND2_X1 U672 ( .A1(n716), .A2(n590), .ZN(n592) );
  XOR2_X1 U673 ( .A(KEYINPUT78), .B(KEYINPUT34), .Z(n591) );
  XNOR2_X1 U674 ( .A(n592), .B(n591), .ZN(n594) );
  NAND2_X1 U675 ( .A1(n594), .A2(n593), .ZN(n597) );
  INV_X1 U676 ( .A(KEYINPUT82), .ZN(n595) );
  XNOR2_X1 U677 ( .A(n595), .B(KEYINPUT35), .ZN(n596) );
  NAND2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U679 ( .A1(KEYINPUT86), .A2(KEYINPUT44), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n600), .A2(KEYINPUT76), .ZN(n601) );
  OR2_X1 U681 ( .A1(n650), .A2(n601), .ZN(n602) );
  NAND2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n626) );
  NAND2_X1 U683 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT85), .ZN(n609) );
  INV_X1 U685 ( .A(n692), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n668) );
  NAND2_X1 U687 ( .A1(n610), .A2(KEYINPUT86), .ZN(n612) );
  NAND2_X1 U688 ( .A1(KEYINPUT76), .A2(KEYINPUT44), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n613) );
  AND2_X1 U690 ( .A1(n668), .A2(n613), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n624) );
  XNOR2_X1 U692 ( .A(n617), .B(KEYINPUT31), .ZN(n684) );
  NOR2_X1 U693 ( .A1(n618), .A2(n695), .ZN(n619) );
  AND2_X1 U694 ( .A1(n590), .A2(n619), .ZN(n671) );
  OR2_X2 U695 ( .A1(n684), .A2(n671), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(KEYINPUT98), .ZN(n622) );
  INV_X1 U697 ( .A(n713), .ZN(n621) );
  AND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n628) );
  INV_X1 U700 ( .A(KEYINPUT45), .ZN(n627) );
  INV_X1 U701 ( .A(KEYINPUT67), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n629), .A2(KEYINPUT2), .ZN(n630) );
  NOR2_X1 U703 ( .A1(n484), .A2(n630), .ZN(n631) );
  INV_X1 U704 ( .A(KEYINPUT2), .ZN(n687) );
  NAND2_X1 U705 ( .A1(n687), .A2(KEYINPUT67), .ZN(n632) );
  AND2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n734), .A2(G478), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(n639) );
  INV_X1 U709 ( .A(G952), .ZN(n638) );
  AND2_X1 U710 ( .A1(n638), .A2(G953), .ZN(n741) );
  NAND2_X1 U711 ( .A1(n661), .A2(G472), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n640), .B(KEYINPUT62), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n644), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U714 ( .A(n645), .B(G134), .ZN(G36) );
  XNOR2_X1 U715 ( .A(n646), .B(G131), .ZN(G33) );
  XOR2_X1 U716 ( .A(G140), .B(KEYINPUT115), .Z(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(G42) );
  XNOR2_X1 U718 ( .A(n649), .B(G110), .ZN(G12) );
  XNOR2_X1 U719 ( .A(n650), .B(G122), .ZN(G24) );
  NAND2_X1 U720 ( .A1(n356), .A2(G217), .ZN(n653) );
  INV_X1 U721 ( .A(n651), .ZN(n652) );
  NOR2_X2 U722 ( .A1(n654), .A2(n741), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(KEYINPUT122), .ZN(G66) );
  NAND2_X1 U724 ( .A1(n661), .A2(G475), .ZN(n658) );
  XOR2_X1 U725 ( .A(KEYINPUT59), .B(n656), .Z(n657) );
  XNOR2_X1 U726 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U727 ( .A(n660), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U728 ( .A1(n356), .A2(G210), .ZN(n665) );
  XOR2_X1 U729 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n662) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X2 U732 ( .A1(n666), .A2(n741), .ZN(n667) );
  XNOR2_X1 U733 ( .A(n667), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U734 ( .A(G101), .B(n668), .ZN(G3) );
  XOR2_X1 U735 ( .A(G104), .B(KEYINPUT113), .Z(n670) );
  NAND2_X1 U736 ( .A1(n671), .A2(n681), .ZN(n669) );
  XNOR2_X1 U737 ( .A(n670), .B(n669), .ZN(G6) );
  XOR2_X1 U738 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n673) );
  NAND2_X1 U739 ( .A1(n671), .A2(n683), .ZN(n672) );
  XNOR2_X1 U740 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U741 ( .A(G107), .B(n674), .ZN(G9) );
  XOR2_X1 U742 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n676) );
  NAND2_X1 U743 ( .A1(n679), .A2(n683), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U745 ( .A(G128), .B(n677), .ZN(G30) );
  XOR2_X1 U746 ( .A(G143), .B(n678), .Z(G45) );
  NAND2_X1 U747 ( .A1(n679), .A2(n681), .ZN(n680) );
  XNOR2_X1 U748 ( .A(n680), .B(G146), .ZN(G48) );
  NAND2_X1 U749 ( .A1(n684), .A2(n681), .ZN(n682) );
  XNOR2_X1 U750 ( .A(n682), .B(G113), .ZN(G15) );
  NAND2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U752 ( .A(n685), .B(G116), .ZN(G18) );
  INV_X1 U753 ( .A(n686), .ZN(n688) );
  NAND2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n732) );
  NAND2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U757 ( .A(n693), .B(KEYINPUT49), .ZN(n694) );
  XNOR2_X1 U758 ( .A(n694), .B(KEYINPUT116), .ZN(n696) );
  NOR2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U760 ( .A(n697), .B(KEYINPUT117), .ZN(n701) );
  NOR2_X1 U761 ( .A1(n587), .A2(n698), .ZN(n699) );
  XNOR2_X1 U762 ( .A(n699), .B(KEYINPUT50), .ZN(n700) );
  NOR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U764 ( .A(n702), .B(KEYINPUT118), .ZN(n703) );
  NOR2_X1 U765 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U766 ( .A(KEYINPUT51), .B(n705), .Z(n706) );
  NOR2_X1 U767 ( .A1(n727), .A2(n706), .ZN(n720) );
  NOR2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U769 ( .A(KEYINPUT119), .B(n709), .Z(n710) );
  NOR2_X1 U770 ( .A1(n711), .A2(n710), .ZN(n715) );
  NOR2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U772 ( .A1(n715), .A2(n714), .ZN(n718) );
  INV_X1 U773 ( .A(n716), .ZN(n717) );
  NOR2_X1 U774 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U775 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U776 ( .A(n721), .B(KEYINPUT52), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n722), .B(KEYINPUT120), .ZN(n725) );
  NAND2_X1 U778 ( .A1(G952), .A2(n723), .ZN(n724) );
  NOR2_X1 U779 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U780 ( .A1(G953), .A2(n726), .ZN(n730) );
  INV_X1 U781 ( .A(n727), .ZN(n728) );
  NAND2_X1 U782 ( .A1(n728), .A2(n716), .ZN(n729) );
  NAND2_X1 U783 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U785 ( .A(KEYINPUT53), .B(n733), .ZN(G75) );
  NAND2_X1 U786 ( .A1(n734), .A2(G469), .ZN(n739) );
  XNOR2_X1 U787 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n735) );
  XNOR2_X1 U788 ( .A(n735), .B(KEYINPUT57), .ZN(n736) );
  XNOR2_X1 U789 ( .A(n737), .B(n736), .ZN(n738) );
  XNOR2_X1 U790 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U791 ( .A1(n741), .A2(n740), .ZN(G54) );
  AND2_X1 U792 ( .A1(KEYINPUT61), .A2(G898), .ZN(n743) );
  NOR2_X1 U793 ( .A1(n385), .A2(n743), .ZN(n744) );
  NOR2_X1 U794 ( .A1(n744), .A2(G953), .ZN(n750) );
  XOR2_X1 U795 ( .A(G224), .B(KEYINPUT61), .Z(n746) );
  NAND2_X1 U796 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U797 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U798 ( .A1(n750), .A2(n749), .ZN(n756) );
  XOR2_X1 U799 ( .A(KEYINPUT123), .B(n751), .Z(n753) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U801 ( .A(n754), .B(KEYINPUT124), .ZN(n755) );
  XNOR2_X1 U802 ( .A(n756), .B(n755), .ZN(G69) );
  XNOR2_X1 U803 ( .A(n758), .B(n757), .ZN(n764) );
  XOR2_X1 U804 ( .A(G227), .B(n764), .Z(n759) );
  XNOR2_X1 U805 ( .A(n759), .B(KEYINPUT125), .ZN(n760) );
  NAND2_X1 U806 ( .A1(n760), .A2(G900), .ZN(n761) );
  XOR2_X1 U807 ( .A(KEYINPUT126), .B(n761), .Z(n762) );
  NOR2_X1 U808 ( .A1(n766), .A2(n762), .ZN(n763) );
  XNOR2_X1 U809 ( .A(n763), .B(KEYINPUT127), .ZN(n769) );
  XNOR2_X1 U810 ( .A(n765), .B(n764), .ZN(n767) );
  NAND2_X1 U811 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U812 ( .A1(n769), .A2(n768), .ZN(G72) );
  XNOR2_X1 U813 ( .A(G137), .B(n770), .ZN(G39) );
  XOR2_X1 U814 ( .A(G119), .B(n771), .Z(G21) );
  XNOR2_X1 U815 ( .A(G125), .B(KEYINPUT37), .ZN(n773) );
  XNOR2_X1 U816 ( .A(n773), .B(n772), .ZN(G27) );
endmodule

