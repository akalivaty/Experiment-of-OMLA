

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U549 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U550 ( .A1(n529), .A2(n528), .ZN(G160) );
  BUF_X1 U551 ( .A(n707), .Z(n708) );
  OR2_X1 U552 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U553 ( .A(n660), .B(n659), .ZN(n666) );
  INV_X1 U554 ( .A(KEYINPUT32), .ZN(n681) );
  NOR2_X1 U555 ( .A1(n695), .A2(n694), .ZN(n705) );
  INV_X1 U556 ( .A(n629), .ZN(n645) );
  OR2_X1 U557 ( .A1(n636), .A2(n965), .ZN(n516) );
  OR2_X1 U558 ( .A1(n670), .A2(n693), .ZN(n517) );
  XNOR2_X1 U559 ( .A(KEYINPUT98), .B(KEYINPUT30), .ZN(n652) );
  XNOR2_X1 U560 ( .A(n653), .B(n652), .ZN(n654) );
  INV_X1 U561 ( .A(KEYINPUT31), .ZN(n658) );
  XNOR2_X1 U562 ( .A(n658), .B(KEYINPUT99), .ZN(n659) );
  OR2_X1 U563 ( .A1(n667), .A2(n666), .ZN(n669) );
  NAND2_X1 U564 ( .A1(n978), .A2(n517), .ZN(n694) );
  NOR2_X1 U565 ( .A1(n578), .A2(n542), .ZN(n788) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n789) );
  INV_X1 U567 ( .A(n772), .ZN(n964) );
  OR2_X1 U568 ( .A1(n535), .A2(n534), .ZN(n536) );
  INV_X1 U569 ( .A(G2104), .ZN(n519) );
  INV_X1 U570 ( .A(G2105), .ZN(n518) );
  NOR2_X2 U571 ( .A1(n519), .A2(n518), .ZN(n881) );
  NAND2_X1 U572 ( .A1(n881), .A2(G113), .ZN(n522) );
  NOR2_X1 U573 ( .A1(G2105), .A2(n519), .ZN(n706) );
  NAND2_X1 U574 ( .A1(G101), .A2(n706), .ZN(n520) );
  XOR2_X1 U575 ( .A(KEYINPUT23), .B(n520), .Z(n521) );
  NAND2_X1 U576 ( .A1(n522), .A2(n521), .ZN(n529) );
  XNOR2_X1 U577 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n524) );
  NOR2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XNOR2_X1 U579 ( .A(n524), .B(n523), .ZN(n707) );
  NAND2_X1 U580 ( .A1(n707), .A2(G137), .ZN(n527) );
  NOR2_X1 U581 ( .A1(n518), .A2(G2104), .ZN(n525) );
  XNOR2_X1 U582 ( .A(n525), .B(KEYINPUT66), .ZN(n711) );
  NAND2_X1 U583 ( .A1(G125), .A2(n711), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U585 ( .A1(G114), .A2(n881), .ZN(n531) );
  BUF_X1 U586 ( .A(n706), .Z(n888) );
  NAND2_X1 U587 ( .A1(G102), .A2(n888), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n707), .A2(G138), .ZN(n533) );
  NAND2_X1 U590 ( .A1(G126), .A2(n711), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U592 ( .A(n536), .B(KEYINPUT89), .ZN(G164) );
  INV_X1 U593 ( .A(G651), .ZN(n542) );
  NOR2_X1 U594 ( .A1(G543), .A2(n542), .ZN(n537) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n537), .Z(n792) );
  NAND2_X1 U596 ( .A1(G65), .A2(n792), .ZN(n540) );
  XOR2_X1 U597 ( .A(G543), .B(KEYINPUT0), .Z(n578) );
  NOR2_X1 U598 ( .A1(G651), .A2(n578), .ZN(n538) );
  XOR2_X2 U599 ( .A(KEYINPUT65), .B(n538), .Z(n793) );
  NAND2_X1 U600 ( .A1(G53), .A2(n793), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U602 ( .A(KEYINPUT70), .B(n541), .Z(n546) );
  NAND2_X1 U603 ( .A1(G78), .A2(n788), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G91), .A2(n789), .ZN(n543) );
  AND2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(G299) );
  NAND2_X1 U607 ( .A1(G64), .A2(n792), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G52), .A2(n793), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U610 ( .A(KEYINPUT69), .B(n549), .Z(n554) );
  NAND2_X1 U611 ( .A1(G77), .A2(n788), .ZN(n551) );
  NAND2_X1 U612 ( .A1(G90), .A2(n789), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U614 ( .A(KEYINPUT9), .B(n552), .Z(n553) );
  NOR2_X1 U615 ( .A1(n554), .A2(n553), .ZN(G171) );
  INV_X1 U616 ( .A(G171), .ZN(G301) );
  NAND2_X1 U617 ( .A1(n789), .A2(G89), .ZN(n555) );
  XNOR2_X1 U618 ( .A(KEYINPUT4), .B(n555), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n788), .A2(G76), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT75), .B(n556), .Z(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(KEYINPUT5), .ZN(n564) );
  NAND2_X1 U623 ( .A1(G63), .A2(n792), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G51), .A2(n793), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U626 ( .A(KEYINPUT6), .B(n562), .Z(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(n789), .A2(G88), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G62), .A2(n792), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G50), .A2(n793), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT82), .B(n568), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G75), .A2(n788), .ZN(n569) );
  XNOR2_X1 U636 ( .A(KEYINPUT83), .B(n569), .ZN(n570) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT84), .B(n574), .Z(G166) );
  XOR2_X1 U640 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  NAND2_X1 U641 ( .A1(G49), .A2(n793), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U644 ( .A1(n792), .A2(n577), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n578), .A2(G87), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(G288) );
  NAND2_X1 U647 ( .A1(G73), .A2(n788), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT2), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n789), .A2(G86), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n582), .B(KEYINPUT80), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G61), .A2(n792), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G48), .A2(n793), .ZN(n585) );
  XNOR2_X1 U654 ( .A(KEYINPUT81), .B(n585), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(G305) );
  NAND2_X1 U657 ( .A1(G72), .A2(n788), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G85), .A2(n789), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U660 ( .A(KEYINPUT68), .B(n592), .Z(n596) );
  NAND2_X1 U661 ( .A1(G60), .A2(n792), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G47), .A2(n793), .ZN(n593) );
  AND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n596), .A2(n595), .ZN(G290) );
  NAND2_X1 U665 ( .A1(G160), .A2(G40), .ZN(n726) );
  XNOR2_X1 U666 ( .A(KEYINPUT93), .B(n726), .ZN(n597) );
  NOR2_X1 U667 ( .A1(G164), .A2(G1384), .ZN(n725) );
  NAND2_X2 U668 ( .A1(n597), .A2(n725), .ZN(n629) );
  NOR2_X1 U669 ( .A1(G2084), .A2(n629), .ZN(n650) );
  NAND2_X1 U670 ( .A1(G8), .A2(n650), .ZN(n598) );
  XNOR2_X1 U671 ( .A(KEYINPUT94), .B(n598), .ZN(n664) );
  NAND2_X1 U672 ( .A1(G8), .A2(n629), .ZN(n670) );
  NOR2_X1 U673 ( .A1(G1966), .A2(n670), .ZN(n662) );
  INV_X1 U674 ( .A(G299), .ZN(n638) );
  INV_X1 U675 ( .A(KEYINPUT96), .ZN(n604) );
  INV_X1 U676 ( .A(G2072), .ZN(n992) );
  NOR2_X1 U677 ( .A1(n629), .A2(n992), .ZN(n600) );
  XOR2_X1 U678 ( .A(KEYINPUT95), .B(KEYINPUT27), .Z(n599) );
  XNOR2_X1 U679 ( .A(n600), .B(n599), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n629), .A2(G1956), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U682 ( .A(n604), .B(n603), .ZN(n637) );
  NOR2_X1 U683 ( .A1(n638), .A2(n637), .ZN(n605) );
  XOR2_X1 U684 ( .A(n605), .B(KEYINPUT28), .Z(n643) );
  AND2_X1 U685 ( .A1(n645), .A2(G1996), .ZN(n607) );
  XOR2_X1 U686 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n606) );
  XNOR2_X1 U687 ( .A(n607), .B(n606), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n629), .A2(G1341), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n635) );
  NAND2_X1 U690 ( .A1(n788), .A2(G68), .ZN(n610) );
  XNOR2_X1 U691 ( .A(KEYINPUT71), .B(n610), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n789), .A2(G81), .ZN(n611) );
  XOR2_X1 U693 ( .A(KEYINPUT12), .B(n611), .Z(n612) );
  NOR2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U695 ( .A(n614), .B(KEYINPUT13), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n792), .A2(G56), .ZN(n615) );
  XOR2_X1 U697 ( .A(KEYINPUT14), .B(n615), .Z(n616) );
  NOR2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U699 ( .A(KEYINPUT72), .B(n618), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G43), .A2(n793), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n772) );
  NAND2_X1 U702 ( .A1(G79), .A2(n788), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G92), .A2(n789), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G66), .A2(n792), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G54), .A2(n793), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U709 ( .A(KEYINPUT15), .B(n627), .Z(n628) );
  XNOR2_X2 U710 ( .A(KEYINPUT73), .B(n628), .ZN(n965) );
  NAND2_X1 U711 ( .A1(G1348), .A2(n629), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n645), .A2(G2067), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U714 ( .A(KEYINPUT97), .B(n632), .Z(n636) );
  NAND2_X1 U715 ( .A1(n965), .A2(n636), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n964), .A2(n633), .ZN(n634) );
  NOR2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n516), .A2(n639), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U721 ( .A(n644), .B(KEYINPUT29), .ZN(n649) );
  NAND2_X1 U722 ( .A1(G1961), .A2(n629), .ZN(n647) );
  XOR2_X1 U723 ( .A(G2078), .B(KEYINPUT25), .Z(n946) );
  NAND2_X1 U724 ( .A1(n645), .A2(n946), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n655) );
  NOR2_X1 U726 ( .A1(G301), .A2(n655), .ZN(n648) );
  NOR2_X1 U727 ( .A1(n649), .A2(n648), .ZN(n667) );
  NOR2_X1 U728 ( .A1(n662), .A2(n650), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n651), .A2(G8), .ZN(n653) );
  NOR2_X1 U730 ( .A1(G168), .A2(n654), .ZN(n657) );
  AND2_X1 U731 ( .A1(G301), .A2(n655), .ZN(n656) );
  NOR2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n660) );
  NOR2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n661) );
  NOR2_X1 U734 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n665), .B(KEYINPUT100), .ZN(n684) );
  AND2_X1 U737 ( .A1(G286), .A2(G8), .ZN(n668) );
  NAND2_X1 U738 ( .A1(n669), .A2(n668), .ZN(n680) );
  INV_X1 U739 ( .A(G8), .ZN(n678) );
  NOR2_X1 U740 ( .A1(G1971), .A2(n670), .ZN(n671) );
  XOR2_X1 U741 ( .A(KEYINPUT101), .B(n671), .Z(n673) );
  NOR2_X1 U742 ( .A1(G2090), .A2(n629), .ZN(n672) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n674), .B(KEYINPUT102), .ZN(n675) );
  NAND2_X1 U745 ( .A1(n675), .A2(G303), .ZN(n676) );
  XOR2_X1 U746 ( .A(KEYINPUT103), .B(n676), .Z(n677) );
  OR2_X1 U747 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U750 ( .A(n685), .B(KEYINPUT104), .ZN(n697) );
  NOR2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n692) );
  NOR2_X1 U752 ( .A1(G1971), .A2(G303), .ZN(n686) );
  NOR2_X1 U753 ( .A1(n692), .A2(n686), .ZN(n982) );
  AND2_X1 U754 ( .A1(n697), .A2(n982), .ZN(n689) );
  NAND2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n968) );
  INV_X1 U756 ( .A(n670), .ZN(n687) );
  NAND2_X1 U757 ( .A1(n968), .A2(n687), .ZN(n688) );
  NOR2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U759 ( .A1(KEYINPUT33), .A2(n690), .ZN(n695) );
  XNOR2_X1 U760 ( .A(G1981), .B(KEYINPUT105), .ZN(n691) );
  XNOR2_X1 U761 ( .A(n691), .B(G305), .ZN(n978) );
  NAND2_X1 U762 ( .A1(n692), .A2(KEYINPUT33), .ZN(n693) );
  NOR2_X1 U763 ( .A1(G2090), .A2(G303), .ZN(n696) );
  NAND2_X1 U764 ( .A1(G8), .A2(n696), .ZN(n698) );
  NAND2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n699), .A2(n670), .ZN(n703) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XOR2_X1 U768 ( .A(n700), .B(KEYINPUT24), .Z(n701) );
  OR2_X1 U769 ( .A1(n670), .A2(n701), .ZN(n702) );
  NAND2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U771 ( .A1(n705), .A2(n704), .ZN(n740) );
  NAND2_X1 U772 ( .A1(G95), .A2(n888), .ZN(n710) );
  NAND2_X1 U773 ( .A1(G131), .A2(n708), .ZN(n709) );
  NAND2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n715) );
  NAND2_X1 U775 ( .A1(G107), .A2(n881), .ZN(n713) );
  BUF_X1 U776 ( .A(n711), .Z(n882) );
  NAND2_X1 U777 ( .A1(G119), .A2(n882), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n870) );
  XOR2_X1 U780 ( .A(KEYINPUT92), .B(G1991), .Z(n945) );
  NOR2_X1 U781 ( .A1(n870), .A2(n945), .ZN(n724) );
  NAND2_X1 U782 ( .A1(G117), .A2(n881), .ZN(n717) );
  NAND2_X1 U783 ( .A1(G129), .A2(n882), .ZN(n716) );
  NAND2_X1 U784 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U785 ( .A1(n888), .A2(G105), .ZN(n718) );
  XOR2_X1 U786 ( .A(KEYINPUT38), .B(n718), .Z(n719) );
  NOR2_X1 U787 ( .A1(n720), .A2(n719), .ZN(n722) );
  NAND2_X1 U788 ( .A1(n708), .A2(G141), .ZN(n721) );
  NAND2_X1 U789 ( .A1(n722), .A2(n721), .ZN(n880) );
  AND2_X1 U790 ( .A1(G1996), .A2(n880), .ZN(n723) );
  NOR2_X1 U791 ( .A1(n724), .A2(n723), .ZN(n1010) );
  NOR2_X1 U792 ( .A1(n726), .A2(n725), .ZN(n755) );
  INV_X1 U793 ( .A(n755), .ZN(n727) );
  NOR2_X1 U794 ( .A1(n1010), .A2(n727), .ZN(n746) );
  INV_X1 U795 ( .A(n746), .ZN(n738) );
  XNOR2_X1 U796 ( .A(G2067), .B(KEYINPUT37), .ZN(n752) );
  NAND2_X1 U797 ( .A1(G104), .A2(n888), .ZN(n729) );
  NAND2_X1 U798 ( .A1(G140), .A2(n708), .ZN(n728) );
  NAND2_X1 U799 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U800 ( .A(KEYINPUT34), .B(n730), .ZN(n736) );
  NAND2_X1 U801 ( .A1(n881), .A2(G116), .ZN(n731) );
  XOR2_X1 U802 ( .A(KEYINPUT91), .B(n731), .Z(n733) );
  NAND2_X1 U803 ( .A1(G128), .A2(n882), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U805 ( .A(KEYINPUT35), .B(n734), .Z(n735) );
  NOR2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U807 ( .A(KEYINPUT36), .B(n737), .ZN(n899) );
  NOR2_X1 U808 ( .A1(n752), .A2(n899), .ZN(n1006) );
  NAND2_X1 U809 ( .A1(n755), .A2(n1006), .ZN(n750) );
  NAND2_X1 U810 ( .A1(n738), .A2(n750), .ZN(n739) );
  NOR2_X1 U811 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U812 ( .A(n741), .B(KEYINPUT106), .ZN(n743) );
  XNOR2_X1 U813 ( .A(G1986), .B(G290), .ZN(n967) );
  NAND2_X1 U814 ( .A1(n755), .A2(n967), .ZN(n742) );
  NAND2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n758) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n880), .ZN(n997) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n744) );
  AND2_X1 U818 ( .A1(n870), .A2(n945), .ZN(n1005) );
  NOR2_X1 U819 ( .A1(n744), .A2(n1005), .ZN(n745) );
  NOR2_X1 U820 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U821 ( .A(KEYINPUT107), .B(n747), .Z(n748) );
  NOR2_X1 U822 ( .A1(n997), .A2(n748), .ZN(n749) );
  XNOR2_X1 U823 ( .A(KEYINPUT39), .B(n749), .ZN(n751) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U825 ( .A1(n752), .A2(n899), .ZN(n1001) );
  NAND2_X1 U826 ( .A1(n753), .A2(n1001), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U828 ( .A(n756), .B(KEYINPUT108), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U830 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U831 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U832 ( .A(G57), .ZN(G237) );
  NAND2_X1 U833 ( .A1(G7), .A2(G661), .ZN(n760) );
  XNOR2_X1 U834 ( .A(n760), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U835 ( .A(G223), .ZN(n826) );
  NAND2_X1 U836 ( .A1(n826), .A2(G567), .ZN(n761) );
  XOR2_X1 U837 ( .A(KEYINPUT11), .B(n761), .Z(G234) );
  NAND2_X1 U838 ( .A1(n964), .A2(G860), .ZN(G153) );
  INV_X1 U839 ( .A(G868), .ZN(n808) );
  NAND2_X1 U840 ( .A1(n965), .A2(n808), .ZN(n762) );
  XNOR2_X1 U841 ( .A(n762), .B(KEYINPUT74), .ZN(n764) );
  NAND2_X1 U842 ( .A1(G868), .A2(G301), .ZN(n763) );
  NAND2_X1 U843 ( .A1(n764), .A2(n763), .ZN(G284) );
  NOR2_X1 U844 ( .A1(G868), .A2(G299), .ZN(n765) );
  XNOR2_X1 U845 ( .A(n765), .B(KEYINPUT76), .ZN(n767) );
  NOR2_X1 U846 ( .A1(n808), .A2(G286), .ZN(n766) );
  NOR2_X1 U847 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U848 ( .A(KEYINPUT77), .B(n768), .Z(G297) );
  INV_X1 U849 ( .A(G860), .ZN(n787) );
  NAND2_X1 U850 ( .A1(n787), .A2(G559), .ZN(n769) );
  INV_X1 U851 ( .A(n965), .ZN(n785) );
  NAND2_X1 U852 ( .A1(n769), .A2(n785), .ZN(n770) );
  XNOR2_X1 U853 ( .A(n770), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U854 ( .A1(n785), .A2(G868), .ZN(n771) );
  NOR2_X1 U855 ( .A1(G559), .A2(n771), .ZN(n774) );
  NOR2_X1 U856 ( .A1(G868), .A2(n772), .ZN(n773) );
  NOR2_X1 U857 ( .A1(n774), .A2(n773), .ZN(G282) );
  XNOR2_X1 U858 ( .A(G2100), .B(KEYINPUT79), .ZN(n784) );
  NAND2_X1 U859 ( .A1(G111), .A2(n881), .ZN(n776) );
  NAND2_X1 U860 ( .A1(G99), .A2(n888), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n781) );
  NAND2_X1 U862 ( .A1(G123), .A2(n882), .ZN(n777) );
  XNOR2_X1 U863 ( .A(n777), .B(KEYINPUT18), .ZN(n779) );
  NAND2_X1 U864 ( .A1(G135), .A2(n708), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n1004) );
  XNOR2_X1 U867 ( .A(n1004), .B(G2096), .ZN(n782) );
  XNOR2_X1 U868 ( .A(n782), .B(KEYINPUT78), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(G156) );
  NAND2_X1 U870 ( .A1(G559), .A2(n785), .ZN(n786) );
  XNOR2_X1 U871 ( .A(n786), .B(n964), .ZN(n805) );
  NAND2_X1 U872 ( .A1(n787), .A2(n805), .ZN(n798) );
  NAND2_X1 U873 ( .A1(G80), .A2(n788), .ZN(n791) );
  NAND2_X1 U874 ( .A1(G93), .A2(n789), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n797) );
  NAND2_X1 U876 ( .A1(G67), .A2(n792), .ZN(n795) );
  NAND2_X1 U877 ( .A1(G55), .A2(n793), .ZN(n794) );
  NAND2_X1 U878 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U879 ( .A1(n797), .A2(n796), .ZN(n807) );
  XOR2_X1 U880 ( .A(n798), .B(n807), .Z(G145) );
  XNOR2_X1 U881 ( .A(KEYINPUT85), .B(G305), .ZN(n799) );
  XNOR2_X1 U882 ( .A(n799), .B(G288), .ZN(n800) );
  XNOR2_X1 U883 ( .A(KEYINPUT19), .B(n800), .ZN(n802) );
  XNOR2_X1 U884 ( .A(G290), .B(n807), .ZN(n801) );
  XNOR2_X1 U885 ( .A(n802), .B(n801), .ZN(n803) );
  XNOR2_X1 U886 ( .A(n803), .B(G299), .ZN(n804) );
  XNOR2_X1 U887 ( .A(n804), .B(G166), .ZN(n906) );
  XOR2_X1 U888 ( .A(n906), .B(n805), .Z(n806) );
  NOR2_X1 U889 ( .A1(n808), .A2(n806), .ZN(n810) );
  AND2_X1 U890 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U891 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U892 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XOR2_X1 U893 ( .A(KEYINPUT20), .B(n811), .Z(n812) );
  NAND2_X1 U894 ( .A1(G2090), .A2(n812), .ZN(n813) );
  XNOR2_X1 U895 ( .A(KEYINPUT21), .B(n813), .ZN(n814) );
  NAND2_X1 U896 ( .A1(n814), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U897 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U898 ( .A1(G483), .A2(G661), .ZN(n824) );
  XOR2_X1 U899 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n816) );
  NAND2_X1 U900 ( .A1(G132), .A2(G82), .ZN(n815) );
  XNOR2_X1 U901 ( .A(n816), .B(n815), .ZN(n817) );
  NAND2_X1 U902 ( .A1(n817), .A2(G96), .ZN(n818) );
  NOR2_X1 U903 ( .A1(n818), .A2(G218), .ZN(n819) );
  XNOR2_X1 U904 ( .A(n819), .B(KEYINPUT87), .ZN(n830) );
  NAND2_X1 U905 ( .A1(n830), .A2(G2106), .ZN(n823) );
  NAND2_X1 U906 ( .A1(G108), .A2(G120), .ZN(n820) );
  NOR2_X1 U907 ( .A1(G237), .A2(n820), .ZN(n821) );
  NAND2_X1 U908 ( .A1(G69), .A2(n821), .ZN(n831) );
  NAND2_X1 U909 ( .A1(n831), .A2(G567), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n823), .A2(n822), .ZN(n915) );
  NOR2_X1 U911 ( .A1(n824), .A2(n915), .ZN(n825) );
  XNOR2_X1 U912 ( .A(n825), .B(KEYINPUT88), .ZN(n829) );
  NAND2_X1 U913 ( .A1(G36), .A2(n829), .ZN(G176) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U916 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n829), .A2(n828), .ZN(G188) );
  XOR2_X1 U919 ( .A(G120), .B(KEYINPUT110), .Z(G236) );
  INV_X1 U921 ( .A(G132), .ZN(G219) );
  INV_X1 U922 ( .A(G108), .ZN(G238) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G82), .ZN(G220) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U927 ( .A(G1341), .B(G2454), .ZN(n832) );
  XNOR2_X1 U928 ( .A(n832), .B(G2430), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n833), .B(G1348), .ZN(n839) );
  XOR2_X1 U930 ( .A(G2443), .B(G2427), .Z(n835) );
  XNOR2_X1 U931 ( .A(G2438), .B(G2446), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n837) );
  XOR2_X1 U933 ( .A(G2451), .B(G2435), .Z(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(n840) );
  NAND2_X1 U936 ( .A1(n840), .A2(G14), .ZN(n841) );
  XNOR2_X1 U937 ( .A(KEYINPUT109), .B(n841), .ZN(G401) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2084), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n842), .B(G2100), .ZN(n852) );
  XOR2_X1 U940 ( .A(KEYINPUT113), .B(G2678), .Z(n844) );
  XNOR2_X1 U941 ( .A(G2096), .B(KEYINPUT43), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U943 ( .A(KEYINPUT112), .B(G2072), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2090), .B(G2078), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U947 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U950 ( .A(G1976), .B(G1971), .Z(n854) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1966), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n855), .B(G2474), .Z(n857) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(KEYINPUT41), .B(G1981), .Z(n859) );
  XNOR2_X1 U957 ( .A(G1961), .B(G1956), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G112), .A2(n881), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G100), .A2(n888), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U963 ( .A1(G136), .A2(n708), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n864), .B(KEYINPUT114), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n882), .A2(G124), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n865), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n872) );
  XNOR2_X1 U970 ( .A(n870), .B(KEYINPUT116), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n898) );
  NAND2_X1 U972 ( .A1(G118), .A2(n881), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G130), .A2(n882), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G106), .A2(n888), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G142), .A2(n708), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n894) );
  XOR2_X1 U980 ( .A(n880), .B(n1004), .Z(n892) );
  NAND2_X1 U981 ( .A1(G115), .A2(n881), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n885), .B(KEYINPUT47), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G139), .A2(n708), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G103), .A2(n888), .ZN(n889) );
  XNOR2_X1 U988 ( .A(KEYINPUT115), .B(n889), .ZN(n890) );
  NOR2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n991) );
  XNOR2_X1 U990 ( .A(n892), .B(n991), .ZN(n893) );
  XOR2_X1 U991 ( .A(n894), .B(n893), .Z(n896) );
  XNOR2_X1 U992 ( .A(G164), .B(G160), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n899), .B(G162), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U997 ( .A1(G37), .A2(n902), .ZN(n903) );
  XOR2_X1 U998 ( .A(KEYINPUT117), .B(n903), .Z(G395) );
  XNOR2_X1 U999 ( .A(n965), .B(KEYINPUT118), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(G171), .B(n964), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n908) );
  XOR2_X1 U1002 ( .A(G286), .B(n906), .Z(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n909), .ZN(G397) );
  OR2_X1 U1005 ( .A1(n915), .A2(G401), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(n915), .ZN(G319) );
  INV_X1 U1013 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1014 ( .A(KEYINPUT125), .B(G1966), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n916), .B(G21), .ZN(n929) );
  XOR2_X1 U1016 ( .A(G1956), .B(G20), .Z(n921) );
  XNOR2_X1 U1017 ( .A(G1341), .B(G19), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(G1981), .B(G6), .ZN(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(KEYINPUT124), .B(n919), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n924) );
  XOR2_X1 U1022 ( .A(KEYINPUT59), .B(G1348), .Z(n922) );
  XNOR2_X1 U1023 ( .A(G4), .B(n922), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1025 ( .A(KEYINPUT60), .B(n925), .Z(n927) );
  XNOR2_X1 U1026 ( .A(G1961), .B(G5), .ZN(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(G1986), .B(G24), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(G1971), .B(G22), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n933) );
  XOR2_X1 U1032 ( .A(G1976), .B(G23), .Z(n932) );
  NAND2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(KEYINPUT58), .B(n934), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1036 ( .A(n937), .B(KEYINPUT126), .Z(n938) );
  XNOR2_X1 U1037 ( .A(KEYINPUT61), .B(n938), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(G16), .A2(n939), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(KEYINPUT127), .B(n940), .ZN(n990) );
  XOR2_X1 U1040 ( .A(G29), .B(KEYINPUT122), .Z(n961) );
  XOR2_X1 U1041 ( .A(G2084), .B(G34), .Z(n941) );
  XNOR2_X1 U1042 ( .A(KEYINPUT54), .B(n941), .ZN(n957) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n955) );
  XOR2_X1 U1044 ( .A(G2067), .B(G26), .Z(n942) );
  NAND2_X1 U1045 ( .A1(n942), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G1996), .B(G32), .ZN(n944) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1048 ( .A1(n944), .A2(n943), .ZN(n950) );
  XOR2_X1 U1049 ( .A(n945), .B(G25), .Z(n948) );
  XNOR2_X1 U1050 ( .A(G27), .B(n946), .ZN(n947) );
  NOR2_X1 U1051 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1052 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n953), .ZN(n954) );
  NOR2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1057 ( .A(n958), .B(KEYINPUT121), .ZN(n959) );
  XNOR2_X1 U1058 ( .A(n959), .B(KEYINPUT55), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n962), .ZN(n988) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n963) );
  XNOR2_X1 U1062 ( .A(n963), .B(KEYINPUT123), .ZN(n986) );
  XNOR2_X1 U1063 ( .A(n964), .B(G1341), .ZN(n977) );
  XNOR2_X1 U1064 ( .A(G1348), .B(n965), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n969) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(G301), .B(G1961), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(G299), .B(G1956), .ZN(n970) );
  NOR2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n973) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n972) );
  NAND2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G168), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(n980), .B(KEYINPUT57), .ZN(n981) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n1020) );
  XOR2_X1 U1082 ( .A(G164), .B(G2078), .Z(n994) );
  XNOR2_X1 U1083 ( .A(n992), .B(n991), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1085 ( .A(KEYINPUT50), .B(n995), .Z(n1000) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(KEYINPUT51), .B(n998), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1014) );
  XOR2_X1 U1091 ( .A(G2084), .B(G160), .Z(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1008) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(KEYINPUT119), .B(n1009), .ZN(n1011) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(KEYINPUT120), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(KEYINPUT52), .B(n1015), .Z(n1016) );
  NOR2_X1 U1100 ( .A1(KEYINPUT55), .A2(n1016), .ZN(n1018) );
  INV_X1 U1101 ( .A(G29), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1021), .ZN(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

