//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1310, new_n1311, new_n1312, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n212), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  INV_X1    g0030(.A(G264), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n206), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n209), .B(new_n220), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT65), .Z(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n239), .B(new_n244), .ZN(G358));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n222), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n230), .A2(G97), .ZN(new_n251));
  INV_X1    g0051(.A(G97), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G107), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n250), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n213), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n267), .A2(new_n202), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(new_n219), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT64), .B(G20), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(KEYINPUT67), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n270), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n278), .A2(new_n262), .B1(new_n202), .B2(new_n260), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n268), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n282), .B1(new_n214), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n288), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n290), .B1(G226), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT3), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G33), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT66), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT66), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(G223), .A3(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G222), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n304), .B1(new_n228), .B2(new_n303), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n294), .B1(new_n308), .B2(new_n291), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n281), .A2(KEYINPUT9), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n281), .A2(KEYINPUT9), .B1(new_n309), .B2(G190), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n309), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT9), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n316), .A2(new_n317), .B1(new_n318), .B2(new_n280), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT10), .B1(new_n319), .B2(new_n311), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n281), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G179), .B2(new_n316), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n303), .A2(G238), .A3(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n298), .A2(new_n302), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G107), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n327), .B(new_n329), .C1(new_n306), .C2(new_n241), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n291), .ZN(new_n331));
  INV_X1    g0131(.A(new_n290), .ZN(new_n332));
  INV_X1    g0132(.A(new_n292), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n229), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(G179), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n266), .A2(G77), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n263), .A2(new_n339), .B1(new_n228), .B2(new_n260), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n224), .A2(KEYINPUT15), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n224), .A2(KEYINPUT15), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT70), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT15), .B(G87), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT70), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n276), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n269), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n228), .A2(new_n274), .B1(new_n277), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n262), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n340), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n334), .B1(new_n330), .B2(new_n291), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(G169), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n337), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n336), .A2(G200), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(KEYINPUT69), .A3(G190), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(KEYINPUT71), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT71), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(new_n340), .C1(new_n351), .C2(new_n352), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n357), .A2(new_n358), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT69), .B1(new_n354), .B2(G190), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n326), .A2(new_n356), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n332), .B1(new_n333), .B2(new_n223), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n214), .A2(new_n283), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n298), .A2(G226), .A3(new_n305), .A4(new_n302), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n298), .A2(G232), .A3(G1698), .A4(new_n302), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G97), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT72), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n368), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT72), .A4(new_n371), .ZN(new_n375));
  AOI211_X1 g0175(.A(KEYINPUT13), .B(new_n367), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT13), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(new_n373), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(new_n375), .A3(new_n291), .ZN(new_n379));
  INV_X1    g0179(.A(new_n367), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n366), .B(G169), .C1(new_n376), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT13), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n379), .A2(new_n377), .A3(new_n380), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(G179), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(G169), .B1(new_n376), .B2(new_n381), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT73), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT14), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n389), .B2(KEYINPUT14), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n273), .A2(G77), .A3(new_n275), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n352), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n396), .A2(KEYINPUT11), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(KEYINPUT11), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n263), .A2(G68), .A3(new_n266), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT12), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n260), .B2(new_n222), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n259), .A2(KEYINPUT12), .A3(G68), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n397), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n393), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n376), .A2(new_n381), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G190), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n408), .B(new_n404), .C1(new_n310), .C2(new_n407), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT74), .B1(new_n272), .B2(KEYINPUT3), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT74), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(new_n295), .A3(G33), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n413), .A3(new_n299), .ZN(new_n414));
  OR2_X1    g0214(.A1(G223), .A2(G1698), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G226), .B2(new_n305), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n414), .A2(new_n416), .B1(new_n272), .B2(new_n224), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n291), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT75), .ZN(new_n419));
  INV_X1    g0219(.A(G179), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n292), .A2(G232), .B1(new_n284), .B2(new_n288), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n418), .A2(new_n419), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT75), .ZN(new_n424));
  AOI21_X1  g0224(.A(G169), .B1(new_n418), .B2(new_n421), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT76), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n428), .B(new_n422), .C1(new_n424), .C2(new_n425), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G58), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n222), .ZN(new_n432));
  OAI21_X1  g0232(.A(G20), .B1(new_n432), .B2(new_n201), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n269), .A2(G159), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n411), .A2(new_n413), .A3(new_n299), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT7), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n274), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(G68), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n414), .B2(new_n215), .ZN(new_n441));
  OAI211_X1 g0241(.A(KEYINPUT16), .B(new_n436), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n299), .A2(new_n300), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n438), .B1(new_n443), .B2(new_n274), .ZN(new_n444));
  NOR2_X1   g0244(.A1(KEYINPUT7), .A2(G20), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n444), .B1(new_n328), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n435), .B1(new_n446), .B2(G68), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n262), .B(new_n442), .C1(new_n447), .C2(KEYINPUT16), .ZN(new_n448));
  INV_X1    g0248(.A(new_n277), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n260), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n267), .B2(new_n449), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n430), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT18), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n427), .A2(new_n429), .B1(new_n452), .B2(new_n448), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n310), .B1(new_n418), .B2(new_n421), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n418), .A2(new_n421), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n459), .B1(G190), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n448), .A2(new_n461), .A3(new_n452), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT17), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n455), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n365), .A2(new_n410), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G116), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n352), .B1(G20), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT84), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n252), .B2(G33), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n274), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n219), .A2(new_n470), .A3(KEYINPUT84), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n467), .B(KEYINPUT20), .C1(new_n472), .C2(new_n473), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n258), .A2(G33), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n352), .A2(new_n259), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT83), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n259), .B2(G116), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n260), .A2(KEYINPUT83), .A3(new_n466), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n481), .A2(G116), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n411), .A2(new_n413), .A3(new_n305), .A4(new_n299), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(G303), .A2(new_n328), .B1(new_n489), .B2(G257), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n231), .A2(new_n305), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n411), .A2(new_n491), .A3(new_n413), .A4(new_n299), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT81), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n492), .B(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n368), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n286), .A2(KEYINPUT5), .ZN(new_n496));
  OR2_X1    g0296(.A1(new_n496), .A2(KEYINPUT77), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(KEYINPUT77), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n258), .B(G45), .C1(new_n286), .C2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n496), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n368), .B1(new_n502), .B2(new_n499), .ZN(new_n503));
  INV_X1    g0303(.A(G270), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n501), .A2(new_n285), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT82), .B1(new_n495), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n328), .A2(G303), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n437), .A2(new_n493), .A3(new_n491), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n437), .A2(G257), .A3(new_n305), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n492), .A2(KEYINPUT81), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n291), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  INV_X1    g0313(.A(new_n505), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n506), .A2(G200), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n506), .A2(new_n515), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n487), .B(new_n516), .C1(new_n517), .C2(new_n317), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n322), .B1(new_n478), .B2(new_n485), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(new_n506), .A3(KEYINPUT21), .A4(new_n515), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n495), .A2(new_n420), .A3(new_n505), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n486), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n519), .A2(new_n506), .A3(new_n515), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n518), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT80), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n343), .A2(new_n346), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(new_n481), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n347), .A2(new_n480), .A3(KEYINPUT80), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n347), .A2(new_n260), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n216), .B(new_n218), .C1(new_n534), .C2(new_n371), .ZN(new_n535));
  OR2_X1    g0335(.A1(KEYINPUT79), .A2(G87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(KEYINPUT79), .A2(G87), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n536), .A2(new_n252), .A3(new_n230), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n274), .A2(new_n299), .A3(new_n411), .A4(new_n413), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n540), .B2(new_n222), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n273), .A2(G97), .A3(new_n275), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n534), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n532), .B(new_n533), .C1(new_n543), .C2(new_n352), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G238), .A2(G1698), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n229), .B2(G1698), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(new_n299), .A3(new_n411), .A4(new_n413), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n368), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT78), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n287), .A2(G1), .A3(G274), .ZN(new_n551));
  AOI21_X1  g0351(.A(G250), .B1(new_n258), .B2(G45), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n291), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n229), .A2(G1698), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(G238), .B2(G1698), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n548), .B1(new_n414), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n553), .B1(new_n557), .B2(new_n291), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(KEYINPUT78), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n322), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n550), .B1(new_n549), .B2(new_n553), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(KEYINPUT78), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n420), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n544), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(G200), .B1(new_n554), .B2(new_n559), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n542), .A2(new_n534), .ZN(new_n566));
  INV_X1    g0366(.A(new_n541), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n262), .B1(new_n260), .B2(new_n347), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n561), .A2(new_n562), .A3(G190), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n481), .A2(G87), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n565), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G257), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G1698), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(G250), .B2(G1698), .ZN(new_n576));
  INV_X1    g0376(.A(G294), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n414), .A2(new_n576), .B1(new_n272), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT87), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n368), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI221_X1 g0380(.A(KEYINPUT87), .B1(new_n272), .B2(new_n577), .C1(new_n414), .C2(new_n576), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n501), .A2(new_n285), .ZN(new_n583));
  INV_X1    g0383(.A(new_n503), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G264), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n322), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n580), .A2(new_n581), .B1(G264), .B2(new_n584), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n420), .A3(new_n583), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT23), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n230), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT23), .B1(new_n215), .B2(G107), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n274), .A2(new_n591), .B1(KEYINPUT85), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n590), .B1(G20), .B2(new_n230), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT85), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n594), .A2(new_n595), .B1(G20), .B2(new_n548), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT86), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n219), .A2(new_n590), .A3(new_n230), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n548), .A2(G20), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(KEYINPUT85), .B2(new_n592), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT86), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n594), .A2(new_n595), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n598), .A2(new_n600), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n298), .A2(G87), .A3(new_n274), .A4(new_n302), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT22), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n414), .A2(new_n219), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n224), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n605), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT24), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT24), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n604), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n352), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT25), .B1(new_n260), .B2(new_n230), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n260), .A2(KEYINPUT25), .A3(new_n230), .ZN(new_n617));
  AOI22_X1  g0417(.A1(G107), .A2(new_n481), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n587), .B(new_n589), .C1(new_n614), .C2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n604), .A2(new_n609), .A3(new_n612), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n612), .B1(new_n604), .B2(new_n609), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n262), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n586), .A2(G200), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n588), .A2(G190), .A3(new_n583), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n623), .A2(new_n618), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n573), .A2(new_n620), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n445), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n298), .B2(new_n302), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n629), .A2(new_n230), .A3(new_n444), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT6), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n251), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(G97), .B(G107), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n632), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  OAI22_X1  g0434(.A1(new_n634), .A2(new_n274), .B1(new_n228), .B2(new_n349), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n262), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n259), .A2(G97), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n481), .B2(G97), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n501), .A2(new_n285), .B1(new_n503), .B2(new_n574), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT4), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n488), .B2(new_n229), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n229), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n298), .A2(new_n305), .A3(new_n302), .A4(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n298), .A2(G250), .A3(G1698), .A4(new_n302), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n642), .A2(new_n644), .A3(new_n645), .A4(new_n469), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n640), .B1(new_n646), .B2(new_n291), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G190), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n639), .B(new_n648), .C1(new_n310), .C2(new_n647), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n646), .A2(new_n291), .ZN(new_n650));
  INV_X1    g0450(.A(new_n640), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n322), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(new_n420), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n636), .A2(new_n638), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n527), .A2(new_n627), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n465), .A2(new_n658), .ZN(G372));
  INV_X1    g0459(.A(new_n324), .ZN(new_n660));
  INV_X1    g0460(.A(new_n409), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n406), .B1(new_n661), .B2(new_n356), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n463), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n455), .A2(new_n458), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n660), .B1(new_n666), .B2(new_n321), .ZN(new_n667));
  INV_X1    g0467(.A(new_n558), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n322), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n544), .A2(new_n563), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(G200), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n569), .A2(new_n570), .A3(new_n671), .A4(new_n571), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n652), .A2(new_n322), .B1(new_n636), .B2(new_n638), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT88), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n654), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n656), .A2(KEYINPUT88), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n673), .A2(new_n674), .A3(new_n677), .A4(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n670), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n564), .A2(new_n572), .A3(new_n654), .A4(new_n675), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(KEYINPUT26), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n620), .A2(new_n526), .A3(new_n522), .A4(new_n520), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n626), .A2(new_n670), .A3(new_n672), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n679), .B(new_n682), .C1(new_n685), .C2(new_n657), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n465), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n667), .A2(new_n687), .ZN(G369));
  NAND2_X1  g0488(.A1(new_n523), .A2(new_n526), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n274), .A2(new_n258), .A3(G13), .ZN(new_n690));
  OAI21_X1  g0490(.A(G213), .B1(new_n690), .B2(KEYINPUT27), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(KEYINPUT27), .B2(new_n690), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n487), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n689), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n527), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  INV_X1    g0500(.A(new_n620), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n695), .B1(new_n614), .B2(new_n619), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n626), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n620), .A2(new_n695), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n704), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n689), .A2(new_n696), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT90), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n707), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n207), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n258), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n538), .A2(G116), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n718), .A2(new_n719), .B1(new_n212), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT94), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n686), .A2(new_n696), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT92), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n649), .B2(new_n656), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n649), .A2(new_n726), .A3(new_n656), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT93), .B1(new_n730), .B2(new_n685), .ZN(new_n731));
  INV_X1    g0531(.A(new_n729), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n727), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT93), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n683), .A4(new_n684), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n670), .B1(new_n681), .B2(KEYINPUT26), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n673), .A2(new_n677), .A3(new_n678), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n736), .B1(KEYINPUT26), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n731), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n696), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n725), .B1(new_n740), .B2(KEYINPUT29), .ZN(new_n741));
  INV_X1    g0541(.A(G330), .ZN(new_n742));
  AOI211_X1 g0542(.A(G179), .B(new_n558), .C1(new_n588), .C2(new_n583), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(new_n506), .A3(new_n515), .A4(new_n652), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  INV_X1    g0545(.A(new_n521), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n647), .A2(new_n588), .A3(new_n561), .A4(new_n562), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n588), .A2(new_n561), .A3(new_n562), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(new_n521), .A3(KEYINPUT30), .A4(new_n647), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n744), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n695), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n658), .B2(new_n696), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n742), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n723), .B1(new_n741), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n741), .A2(new_n723), .A3(new_n758), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n722), .B1(new_n762), .B2(G1), .ZN(G364));
  NAND3_X1  g0563(.A1(new_n274), .A2(G13), .A3(G45), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n718), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n699), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n213), .B1(G20), .B2(new_n322), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n437), .A2(new_n716), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n287), .B2(new_n212), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n250), .B2(new_n287), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n328), .A2(new_n716), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G355), .B1(new_n466), .B2(new_n716), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n773), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n215), .A2(new_n317), .A3(new_n310), .A4(G179), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n328), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n317), .A2(G200), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n274), .B1(new_n420), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n784), .B1(G294), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n274), .A2(new_n420), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n790), .A2(G190), .A3(new_n310), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(KEYINPUT33), .B(G317), .Z(new_n793));
  INV_X1    g0593(.A(G326), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n790), .A2(new_n317), .A3(new_n310), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n788), .B1(new_n792), .B2(new_n793), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G179), .A2(G190), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n219), .A2(G200), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G283), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n789), .A2(new_n785), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n219), .A2(new_n310), .A3(new_n798), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n803), .A2(G322), .B1(G329), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n789), .A2(new_n317), .A3(new_n310), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT95), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n801), .B(new_n806), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G159), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n804), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT32), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n817), .B1(new_n792), .B2(new_n222), .C1(new_n202), .C2(new_n796), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n799), .A2(new_n230), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n536), .A2(new_n537), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n328), .B(new_n819), .C1(new_n820), .C2(new_n781), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n803), .A2(G58), .B1(new_n787), .B2(G97), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n821), .B(new_n822), .C1(new_n812), .C2(new_n228), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n797), .A2(new_n814), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n780), .B1(new_n824), .B2(new_n771), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n765), .B1(new_n770), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n765), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n699), .A2(G330), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(new_n828), .B2(new_n700), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT96), .ZN(G396));
  NOR3_X1   g0631(.A1(new_n337), .A2(new_n355), .A3(new_n695), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n695), .A2(new_n353), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n362), .B2(new_n363), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n832), .B1(new_n834), .B2(new_n356), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT99), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n835), .B(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n724), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n649), .A2(new_n656), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n683), .A2(new_n840), .A3(new_n684), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n682), .A2(new_n679), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n835), .B(new_n696), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT100), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n686), .A2(KEYINPUT100), .A3(new_n696), .A4(new_n835), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n839), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n848), .A2(new_n757), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n765), .B1(new_n848), .B2(new_n757), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n835), .A2(new_n767), .ZN(new_n851));
  INV_X1    g0651(.A(new_n771), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n791), .A2(G283), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n303), .B1(G107), .B2(new_n781), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(new_n252), .C2(new_n786), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n803), .A2(G294), .B1(G87), .B2(new_n800), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n856), .B1(new_n813), .B2(new_n804), .C1(new_n812), .C2(new_n466), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n855), .B(new_n857), .C1(G303), .C2(new_n795), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT97), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n795), .A2(G137), .B1(G143), .B2(new_n803), .ZN(new_n860));
  INV_X1    g0660(.A(G150), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n860), .B1(new_n861), .B2(new_n792), .C1(new_n812), .C2(new_n815), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(KEYINPUT34), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n863), .A2(KEYINPUT34), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n800), .A2(G68), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n866), .B(new_n437), .C1(new_n202), .C2(new_n782), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n786), .A2(new_n431), .B1(new_n804), .B2(new_n868), .ZN(new_n869));
  OR3_X1    g0669(.A1(new_n865), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n859), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT98), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n852), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n872), .B2(new_n871), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n771), .A2(new_n766), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n874), .B(new_n827), .C1(G77), .C2(new_n876), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n849), .A2(new_n850), .B1(new_n851), .B2(new_n877), .ZN(G384));
  INV_X1    g0678(.A(KEYINPUT89), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n692), .B(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n665), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n405), .B(new_n695), .C1(new_n393), .C2(new_n661), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n405), .A2(new_n695), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n322), .B1(new_n384), .B2(new_n385), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT73), .B1(new_n884), .B2(new_n366), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT14), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n387), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n409), .B(new_n883), .C1(new_n887), .C2(new_n404), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n832), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n847), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  INV_X1    g0693(.A(new_n442), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n414), .A2(new_n215), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT7), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n216), .A2(new_n218), .A3(new_n438), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n222), .B1(new_n897), .B2(new_n414), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n435), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n262), .B1(new_n899), .B2(KEYINPUT16), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n894), .B1(new_n900), .B2(KEYINPUT102), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT102), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n902), .B(new_n262), .C1(new_n899), .C2(KEYINPUT16), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n451), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n462), .B1(new_n904), .B2(new_n693), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n900), .A2(KEYINPUT102), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n442), .A3(new_n903), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n427), .A2(new_n429), .B1(new_n907), .B2(new_n452), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT103), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT104), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n453), .A2(new_n880), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n454), .A2(new_n912), .A3(new_n462), .A4(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT103), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n915), .B(KEYINPUT37), .C1(new_n905), .C2(new_n908), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n910), .A2(new_n911), .A3(new_n914), .A4(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n436), .B1(new_n440), .B2(new_n441), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT16), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n352), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n442), .B1(new_n920), .B2(new_n902), .ZN(new_n921));
  INV_X1    g0721(.A(new_n903), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n452), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n464), .A2(new_n880), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n913), .A2(new_n462), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n456), .A2(new_n926), .A3(KEYINPUT37), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n448), .A2(new_n461), .A3(new_n452), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n923), .B2(new_n880), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n430), .A2(new_n923), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n912), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n927), .B1(new_n931), .B2(new_n915), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n911), .B1(new_n932), .B2(new_n910), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n893), .B1(new_n925), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n916), .A2(new_n914), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n929), .A2(new_n930), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n915), .B1(new_n936), .B2(KEYINPUT37), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT104), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n938), .A2(new_n917), .A3(KEYINPUT38), .A4(new_n924), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n881), .B1(new_n892), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n913), .B1(new_n665), .B2(new_n463), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT37), .B1(new_n456), .B2(new_n926), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n914), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n893), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n934), .A2(KEYINPUT39), .A3(new_n939), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n406), .A2(new_n695), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n941), .A2(new_n951), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n365), .A2(new_n410), .A3(new_n464), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n741), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n664), .B1(new_n662), .B2(new_n463), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n315), .A2(new_n320), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n324), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n952), .B(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT105), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n752), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n751), .A2(KEYINPUT105), .A3(new_n695), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n753), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n627), .A2(new_n657), .ZN(new_n964));
  INV_X1    g0764(.A(new_n527), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n964), .A2(new_n965), .A3(new_n696), .ZN(new_n966));
  INV_X1    g0766(.A(new_n754), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n889), .A2(new_n835), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n946), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT40), .ZN(new_n971));
  AND4_X1   g0771(.A1(new_n971), .A2(new_n889), .A3(new_n835), .A4(new_n968), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n970), .A2(KEYINPUT40), .B1(new_n940), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n465), .A2(new_n968), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n742), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n975), .B2(new_n974), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n959), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n978), .A2(KEYINPUT106), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(KEYINPUT106), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n959), .A2(new_n977), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n258), .B1(new_n274), .B2(G13), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n979), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n634), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT35), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n274), .A2(new_n466), .A3(new_n213), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n984), .B2(KEYINPUT35), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT101), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n988), .B2(new_n987), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT36), .ZN(new_n991));
  OR3_X1    g0791(.A1(new_n211), .A2(new_n228), .A3(new_n432), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n258), .B(G13), .C1(new_n992), .C2(new_n246), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n983), .A2(new_n991), .A3(new_n993), .ZN(G367));
  AOI22_X1  g0794(.A1(new_n787), .A2(G68), .B1(new_n805), .B2(G137), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n861), .B2(new_n802), .ZN(new_n996));
  INV_X1    g0796(.A(new_n812), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(G50), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n799), .A2(new_n228), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n303), .B1(new_n431), .B2(new_n782), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(G143), .C2(new_n795), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n998), .B(new_n1001), .C1(new_n815), .C2(new_n792), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n997), .A2(G283), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n799), .A2(new_n252), .ZN(new_n1004));
  INV_X1    g0804(.A(G317), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n802), .A2(new_n783), .B1(new_n1005), .B2(new_n804), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(G107), .C2(new_n787), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n795), .A2(G311), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT46), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n782), .B2(new_n466), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n414), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G294), .B2(new_n791), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1003), .A2(new_n1007), .A3(new_n1008), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1002), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT47), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n771), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n773), .B1(new_n529), .B2(new_n716), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n238), .A2(new_n774), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n765), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n569), .A2(new_n571), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n695), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n673), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n680), .A2(new_n1021), .A3(new_n695), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(KEYINPUT107), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(KEYINPUT107), .B2(new_n1024), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1017), .B(new_n1020), .C1(new_n1027), .C2(new_n769), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n764), .A2(G1), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n696), .A2(new_n639), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n730), .A2(new_n1030), .B1(new_n656), .B2(new_n696), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n712), .A2(new_n713), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT44), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  AND3_X1   g0836(.A1(new_n714), .A2(KEYINPUT45), .A3(new_n1031), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT45), .B1(new_n714), .B2(new_n1031), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n1035), .A2(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n706), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n707), .B1(new_n1037), .B2(new_n1038), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n705), .B(new_n709), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(new_n700), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n762), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(KEYINPUT110), .B(KEYINPUT41), .Z(new_n1046));
  XNOR2_X1  g0846(.A(new_n717), .B(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1029), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1031), .B(KEYINPUT108), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT109), .B1(new_n707), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n707), .A2(new_n1049), .A3(KEYINPUT109), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1027), .A2(KEYINPUT43), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1053), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n656), .B1(new_n1049), .B2(new_n620), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n694), .B2(new_n693), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1032), .A2(new_n705), .A3(new_n709), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT42), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1027), .A2(KEYINPUT43), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1057), .B(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1028), .B1(new_n1048), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT111), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(KEYINPUT111), .B(new_n1028), .C1(new_n1048), .C2(new_n1065), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(G387));
  INV_X1    g0871(.A(new_n1044), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n762), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n760), .A2(new_n761), .A3(new_n1044), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n717), .A3(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n719), .B(KEYINPUT112), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n287), .B1(new_n222), .B2(new_n228), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n277), .A2(G50), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT50), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1076), .B(new_n1080), .C1(new_n1079), .C2(new_n1078), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1081), .B(new_n774), .C1(new_n244), .C2(new_n287), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n778), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1082), .B1(G107), .B2(new_n207), .C1(new_n719), .C2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n765), .B1(new_n1084), .B2(new_n772), .ZN(new_n1085));
  OR3_X1    g0885(.A1(new_n796), .A2(KEYINPUT113), .A3(new_n815), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT113), .B1(new_n796), .B2(new_n815), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n812), .C2(new_n222), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n347), .A2(new_n786), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n802), .A2(new_n202), .B1(new_n861), .B2(new_n804), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n414), .B(new_n1004), .C1(G77), .C2(new_n781), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n277), .B2(new_n792), .ZN(new_n1092));
  NOR4_X1   g0892(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n791), .A2(G311), .B1(G317), .B2(new_n803), .ZN(new_n1094));
  INV_X1    g0894(.A(G322), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1094), .B1(new_n1095), .B2(new_n796), .C1(new_n812), .C2(new_n783), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT48), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n787), .A2(G283), .B1(new_n781), .B2(G294), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT114), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT49), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n414), .B1(new_n799), .B2(new_n466), .C1(new_n794), .C2(new_n804), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT115), .Z(new_n1106));
  NOR2_X1   g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1093), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1085), .B1(new_n1109), .B2(new_n852), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n705), .B2(new_n768), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1072), .B2(new_n1029), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1075), .A2(new_n1112), .ZN(G393));
  INV_X1    g0913(.A(new_n1042), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1073), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1042), .A2(new_n1073), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n717), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1049), .A2(new_n768), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n787), .A2(G77), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n202), .B2(new_n792), .C1(new_n812), .C2(new_n277), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT116), .Z(new_n1122));
  OAI221_X1 g0922(.A(new_n437), .B1(new_n799), .B2(new_n224), .C1(new_n782), .C2(new_n222), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n795), .A2(G150), .B1(G159), .B2(new_n803), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT51), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(G143), .C2(new_n805), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n792), .A2(new_n783), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n303), .B(new_n819), .C1(G283), .C2(new_n781), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n466), .B2(new_n786), .C1(new_n1095), .C2(new_n804), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1127), .B(new_n1129), .C1(G294), .C2(new_n997), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n795), .A2(G317), .B1(G311), .B2(new_n803), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT52), .Z(new_n1132));
  AOI22_X1  g0932(.A1(new_n1122), .A2(new_n1126), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1133), .A2(new_n852), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n775), .A2(new_n256), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n773), .B(new_n1135), .C1(G97), .C2(new_n716), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1134), .A2(new_n765), .A3(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT117), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1114), .A2(new_n1029), .B1(new_n1119), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1118), .A2(new_n1139), .ZN(G390));
  AOI21_X1  g0940(.A(new_n767), .B1(new_n948), .B2(new_n949), .ZN(new_n1141));
  OR3_X1    g0941(.A1(new_n782), .A2(KEYINPUT53), .A3(new_n861), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT53), .B1(new_n782), .B2(new_n861), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n303), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n796), .A2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(G137), .C2(new_n791), .ZN(new_n1147));
  INV_X1    g0947(.A(G125), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n202), .A2(new_n799), .B1(new_n804), .B2(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n802), .A2(new_n868), .B1(new_n786), .B2(new_n815), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT54), .B(G143), .Z(new_n1151));
  AOI211_X1 g0951(.A(new_n1149), .B(new_n1150), .C1(new_n997), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n795), .A2(G283), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n303), .B1(G87), .B2(new_n781), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n866), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G107), .B2(new_n791), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1120), .B1(new_n577), .B2(new_n804), .C1(new_n802), .C2(new_n466), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n997), .B2(G97), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1147), .A2(new_n1152), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n827), .B1(new_n449), .B2(new_n876), .C1(new_n1159), .C2(new_n852), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1141), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT118), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n847), .A2(new_n891), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n889), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n950), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1164), .A2(new_n1165), .B1(new_n948), .B2(new_n949), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n757), .A2(new_n835), .A3(new_n889), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n946), .A2(new_n1165), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n834), .A2(new_n356), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n739), .A2(new_n696), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n890), .B1(new_n1170), .B2(new_n891), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1167), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1162), .B1(new_n1166), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n948), .A2(new_n949), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n832), .B1(new_n845), .B2(new_n846), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1165), .B1(new_n1175), .B2(new_n890), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1167), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1170), .A2(new_n891), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n889), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n950), .B1(new_n939), .B2(new_n945), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1177), .A2(new_n1182), .A3(KEYINPUT118), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1177), .A2(new_n1185), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n889), .A2(new_n835), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n742), .B1(new_n755), .B2(new_n963), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1173), .A2(new_n1183), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1161), .B1(new_n1190), .B2(new_n1029), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n465), .A2(new_n1188), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n667), .B(new_n1192), .C1(new_n953), .C2(new_n741), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n967), .A2(new_n966), .A3(new_n756), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(G330), .A3(new_n835), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1187), .A2(new_n1188), .B1(new_n890), .B2(new_n1195), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(new_n1175), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n837), .A2(G330), .A3(new_n968), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n890), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1199), .A2(new_n1167), .A3(new_n891), .A4(new_n1170), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1193), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n717), .B1(new_n1190), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1189), .B1(new_n1166), .B2(new_n1184), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1166), .A2(new_n1162), .A3(new_n1172), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT118), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1201), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1191), .B1(new_n1202), .B2(new_n1207), .ZN(G378));
  OAI21_X1  g1008(.A(new_n827), .B1(G50), .B2(new_n876), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n281), .A2(new_n693), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n325), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n325), .A2(new_n1210), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OR3_X1    g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(new_n767), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n800), .A2(G58), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT119), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n414), .B(new_n286), .C1(new_n782), .C2(new_n228), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G283), .B2(new_n805), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT120), .Z(new_n1224));
  OAI22_X1  g1024(.A1(new_n796), .A2(new_n466), .B1(new_n222), .B2(new_n786), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT121), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n802), .B2(new_n230), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n803), .A2(KEYINPUT121), .A3(G107), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n792), .C2(new_n252), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1225), .B(new_n1229), .C1(new_n529), .C2(new_n997), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n414), .A2(new_n286), .ZN(new_n1232));
  AOI21_X1  g1032(.A(G50), .B1(new_n272), .B2(new_n286), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1231), .A2(KEYINPUT58), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G125), .A2(new_n795), .B1(new_n791), .B2(G132), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n787), .A2(G150), .B1(new_n781), .B2(new_n1151), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n1145), .C2(new_n802), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G137), .B2(new_n997), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n800), .A2(G159), .ZN(new_n1242));
  AOI211_X1 g1042(.A(G33), .B(G41), .C1(new_n805), .C2(G124), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1234), .B1(KEYINPUT58), .B2(new_n1231), .C1(new_n1240), .C2(new_n1244), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1209), .B(new_n1218), .C1(new_n771), .C2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1217), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n973), .B2(new_n742), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n971), .B1(new_n969), .B2(new_n946), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n889), .A2(new_n968), .A3(new_n971), .A4(new_n835), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n939), .B2(new_n934), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G330), .B(new_n1217), .C1(new_n1249), .C2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n952), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1248), .A2(new_n952), .A3(new_n1252), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1246), .B1(new_n1257), .B2(new_n1029), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1193), .B1(new_n1190), .B2(new_n1201), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1248), .A2(new_n952), .A3(new_n1252), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n952), .B1(new_n1248), .B2(new_n1252), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT57), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n717), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1193), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1206), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT57), .B1(new_n1265), .B2(new_n1257), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1258), .B1(new_n1263), .B2(new_n1266), .ZN(G375));
  INV_X1    g1067(.A(new_n1201), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1197), .A2(new_n1193), .A3(new_n1200), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1047), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1200), .B1(new_n1175), .B2(new_n1196), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n890), .A2(new_n766), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n827), .B1(G68), .B2(new_n876), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n997), .A2(G107), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n795), .A2(G294), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n328), .B1(new_n782), .B2(new_n252), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n999), .B(new_n1276), .C1(new_n791), .C2(G116), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n804), .A2(new_n783), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1278), .B(new_n1089), .C1(G283), .C2(new_n803), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1274), .A2(new_n1275), .A3(new_n1277), .A4(new_n1279), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n812), .A2(new_n861), .B1(new_n202), .B2(new_n786), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT123), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n795), .A2(G132), .ZN(new_n1283));
  XOR2_X1   g1083(.A(new_n1283), .B(KEYINPUT122), .Z(new_n1284));
  NOR2_X1   g1084(.A1(new_n804), .A2(new_n1145), .ZN(new_n1285));
  INV_X1    g1085(.A(G137), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n437), .B1(new_n782), .B2(new_n815), .C1(new_n802), .C2(new_n1286), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1285), .B(new_n1287), .C1(new_n791), .C2(new_n1151), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1284), .A2(new_n1220), .A3(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1280), .B1(new_n1282), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1273), .B1(new_n1290), .B2(new_n771), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1271), .A2(new_n1029), .B1(new_n1272), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1270), .A2(new_n1292), .ZN(new_n1293));
  XOR2_X1   g1093(.A(new_n1293), .B(KEYINPUT124), .Z(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(G381));
  INV_X1    g1095(.A(KEYINPUT125), .ZN(new_n1296));
  NOR4_X1   g1096(.A1(G393), .A2(new_n1296), .A3(G396), .A4(G384), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(G393), .A2(G396), .ZN(new_n1298));
  INV_X1    g1098(.A(G384), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT125), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NOR4_X1   g1100(.A1(G381), .A2(new_n1297), .A3(G390), .A4(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1029), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n1302), .A2(new_n1303), .B1(new_n1141), .B2(new_n1160), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n717), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1302), .B2(new_n1268), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1304), .B1(new_n1306), .B2(new_n1206), .ZN(new_n1307));
  INV_X1    g1107(.A(G375), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1301), .A2(new_n1070), .A3(new_n1307), .A4(new_n1308), .ZN(G407));
  NAND2_X1  g1109(.A1(new_n694), .A2(G213), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1308), .A2(new_n1307), .A3(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(G407), .A2(G213), .A3(new_n1312), .ZN(G409));
  OAI211_X1 g1113(.A(G378), .B(new_n1258), .C1(new_n1263), .C2(new_n1266), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1265), .A2(new_n1047), .A3(new_n1257), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1258), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1307), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1310), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1311), .A2(G2897), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT126), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT60), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1323), .B1(new_n1264), .B2(new_n1271), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1264), .A2(new_n1271), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1322), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(KEYINPUT126), .B(new_n1269), .C1(new_n1201), .C2(new_n1323), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1305), .B1(new_n1325), .B2(KEYINPUT60), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1326), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1329), .A2(G384), .A3(new_n1292), .ZN(new_n1330));
  AOI21_X1  g1130(.A(G384), .B1(new_n1329), .B2(new_n1292), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1321), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1329), .A2(new_n1292), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1299), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1329), .A2(G384), .A3(new_n1292), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n1335), .A3(new_n1320), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1332), .A2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT61), .B1(new_n1319), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT63), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1339), .B1(new_n1319), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1066), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(G390), .ZN(new_n1344));
  INV_X1    g1144(.A(G390), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1066), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(G396), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(G393), .B(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT127), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1349), .B(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1347), .A2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1068), .A2(new_n1069), .A3(new_n1345), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1349), .B1(new_n1343), .B2(G390), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1352), .A2(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1311), .B1(new_n1314), .B2(new_n1317), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1357), .A2(KEYINPUT63), .A3(new_n1340), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1338), .A2(new_n1342), .A3(new_n1356), .A4(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT62), .ZN(new_n1360));
  AND3_X1   g1160(.A1(new_n1357), .A2(new_n1360), .A3(new_n1340), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT61), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1332), .A2(new_n1336), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1362), .B1(new_n1357), .B2(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1360), .B1(new_n1357), .B2(new_n1340), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1361), .A2(new_n1364), .A3(new_n1365), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1359), .B1(new_n1366), .B2(new_n1356), .ZN(G405));
  NAND2_X1  g1167(.A1(G375), .A2(new_n1307), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1368), .A2(new_n1314), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1369), .A2(new_n1340), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1341), .A2(new_n1368), .A3(new_n1314), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  AOI22_X1  g1172(.A1(new_n1347), .A2(new_n1351), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1373));
  XNOR2_X1  g1173(.A(new_n1372), .B(new_n1373), .ZN(G402));
endmodule


