//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n202));
  INV_X1    g001(.A(G134gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G127gat), .ZN(new_n204));
  INV_X1    g003(.A(G127gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G134gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G113gat), .ZN(new_n211));
  INV_X1    g010(.A(G113gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G120gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G134gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n209), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G169gat), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT23), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT24), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n229), .B2(new_n226), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n225), .B(new_n230), .C1(KEYINPUT65), .C2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n221), .A2(new_n223), .A3(KEYINPUT65), .A4(new_n224), .ZN(new_n233));
  AND3_X1   g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n226), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(new_n228), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n237));
  OAI211_X1 g036(.A(KEYINPUT25), .B(new_n233), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT26), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(new_n224), .ZN(new_n242));
  NOR3_X1   g041(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n235), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  NAND2_X1  g044(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n246), .A2(KEYINPUT27), .ZN(new_n247));
  INV_X1    g046(.A(G190gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n246), .B2(KEYINPUT27), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n245), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT27), .B(G183gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT28), .A3(new_n248), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n244), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n218), .B1(new_n239), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n244), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n252), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n209), .A2(new_n217), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n232), .A4(new_n238), .ZN(new_n259));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT64), .Z(new_n261));
  NAND3_X1  g060(.A1(new_n254), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT67), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n254), .A2(new_n259), .A3(new_n264), .A4(new_n261), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n202), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT33), .ZN(new_n267));
  XNOR2_X1  g066(.A(G15gat), .B(G43gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(G71gat), .B(G99gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n270), .B(KEYINPUT69), .Z(new_n271));
  OAI21_X1  g070(.A(new_n266), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT33), .B1(new_n263), .B2(new_n265), .ZN(new_n273));
  NOR4_X1   g072(.A1(new_n273), .A2(new_n266), .A3(KEYINPUT68), .A4(new_n270), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n263), .A2(new_n265), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n270), .B1(new_n276), .B2(KEYINPUT32), .ZN(new_n277));
  INV_X1    g076(.A(new_n273), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n272), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n254), .A2(new_n259), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n260), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT34), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n261), .A2(KEYINPUT34), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G22gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT2), .ZN(new_n291));
  OR2_X1    g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT75), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n295), .A3(new_n293), .ZN(new_n296));
  INV_X1    g095(.A(new_n290), .ZN(new_n297));
  NOR2_X1   g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n294), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G155gat), .B(G162gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n303), .B(new_n291), .C1(new_n304), .C2(new_n295), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n310));
  NAND2_X1  g109(.A1(G211gat), .A2(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT22), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G204gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G197gat), .ZN(new_n315));
  INV_X1    g114(.A(G197gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G204gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n311), .ZN(new_n319));
  NOR2_X1   g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n310), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G211gat), .B(G218gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(G197gat), .B(G204gat), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT70), .A4(new_n313), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(new_n321), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n322), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G228gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n322), .A2(new_n325), .A3(new_n326), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT3), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n300), .A2(new_n305), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n328), .B(new_n330), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT3), .B1(new_n331), .B2(new_n308), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n328), .B1(new_n337), .B2(new_n334), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n335), .A2(new_n336), .B1(new_n338), .B2(new_n329), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n329), .B1(new_n309), .B2(new_n327), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n340), .B(KEYINPUT79), .C1(new_n334), .C2(new_n333), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n289), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n328), .A2(new_n330), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n331), .A2(new_n332), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n334), .B1(new_n344), .B2(new_n306), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n336), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n308), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n334), .B1(new_n347), .B2(new_n306), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n331), .B1(new_n307), .B2(new_n308), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n329), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n346), .A2(new_n341), .A3(new_n350), .A4(new_n289), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT31), .B(G50gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n342), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n351), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n339), .A2(KEYINPUT80), .A3(new_n289), .A4(new_n341), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n341), .A3(new_n350), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n363), .A2(new_n364), .A3(G22gat), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n363), .B2(G22gat), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n358), .B1(new_n367), .B2(new_n355), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n272), .B(new_n286), .C1(new_n274), .C2(new_n279), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n288), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT71), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n239), .B2(new_n253), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n257), .A2(KEYINPUT71), .A3(new_n232), .A4(new_n238), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n308), .ZN(new_n377));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(KEYINPUT73), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n257), .A2(new_n232), .A3(new_n238), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(G226gat), .A3(G233gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT73), .B1(new_n377), .B2(new_n378), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n327), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n380), .A2(new_n332), .A3(new_n378), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n375), .A2(new_n376), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(new_n378), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n331), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n384), .A2(KEYINPUT74), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT74), .B1(new_n384), .B2(new_n388), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n373), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n373), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n384), .A2(new_n392), .A3(new_n388), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT30), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT30), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n384), .A2(new_n395), .A3(new_n392), .A4(new_n388), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT0), .ZN(new_n399));
  XNOR2_X1  g198(.A(G57gat), .B(G85gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n300), .A2(new_n305), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n218), .B1(KEYINPUT3), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n404), .B1(new_n406), .B2(new_n307), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT77), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n334), .A2(new_n408), .A3(new_n218), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT77), .B1(new_n405), .B2(new_n258), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT4), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n405), .A2(new_n258), .ZN(new_n412));
  XOR2_X1   g211(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n407), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n405), .A2(new_n258), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n409), .A2(new_n410), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(new_n404), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n409), .A2(KEYINPUT4), .A3(new_n410), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n412), .A2(new_n413), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT78), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n406), .A2(new_n307), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n404), .A2(KEYINPUT5), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n421), .A2(new_n422), .B1(new_n307), .B2(new_n406), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n424), .B1(new_n429), .B2(new_n426), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n402), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n423), .A2(new_n425), .A3(new_n426), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT78), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n434), .A2(new_n401), .A3(new_n427), .A4(new_n420), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(KEYINPUT6), .B(new_n402), .C1(new_n428), .C2(new_n430), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n391), .A2(new_n397), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n370), .B(new_n440), .C1(KEYINPUT88), .C2(KEYINPUT35), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n288), .A2(new_n368), .A3(KEYINPUT88), .A4(new_n369), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT35), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n288), .A2(new_n368), .A3(new_n369), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n442), .B(new_n443), .C1(new_n444), .C2(new_n439), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n436), .A2(new_n437), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n392), .A2(KEYINPUT38), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n331), .B1(new_n382), .B2(new_n383), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT37), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n387), .B2(new_n327), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n454));
  NAND3_X1  g253(.A1(new_n384), .A2(new_n388), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n447), .A2(new_n448), .A3(new_n456), .A4(new_n393), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n437), .A3(new_n393), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n453), .A2(new_n455), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT86), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n384), .A2(new_n388), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT74), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n384), .A2(KEYINPUT74), .A3(new_n388), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n451), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n462), .B1(new_n467), .B2(new_n392), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT37), .B1(new_n389), .B2(new_n390), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(KEYINPUT87), .A3(new_n373), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(new_n455), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n461), .B1(new_n471), .B2(KEYINPUT38), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n429), .A2(new_n403), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n473), .A2(KEYINPUT39), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n473), .B(KEYINPUT39), .C1(new_n404), .C2(new_n418), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n474), .A2(new_n475), .A3(new_n401), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT40), .A4(new_n401), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  OAI221_X1 g279(.A(new_n431), .B1(KEYINPUT40), .B2(new_n476), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n391), .A2(new_n397), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n368), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n472), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n365), .A2(new_n366), .ZN(new_n485));
  INV_X1    g284(.A(new_n362), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n355), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT82), .B1(new_n487), .B2(new_n357), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT82), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(new_n358), .C1(new_n367), .C2(new_n355), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n439), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n288), .A2(new_n369), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT36), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n288), .A2(new_n494), .A3(new_n369), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT83), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n491), .A2(new_n493), .A3(new_n498), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n446), .B1(new_n484), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G113gat), .B(G141gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT11), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(new_n219), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(G197gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT12), .Z(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G43gat), .B(G50gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(KEYINPUT90), .ZN(new_n514));
  OR3_X1    g313(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n515));
  MUX2_X1   g314(.A(KEYINPUT90), .B(new_n514), .S(new_n515), .Z(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  INV_X1    g316(.A(G36gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(KEYINPUT15), .B(new_n511), .C1(new_n516), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n515), .B1(new_n513), .B2(KEYINPUT91), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(KEYINPUT91), .B2(new_n515), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n509), .A2(KEYINPUT15), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(new_n519), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G8gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT16), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(G1gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(G1gat), .B2(new_n529), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n527), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n527), .B(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n508), .B(new_n538), .C1(new_n540), .C2(new_n537), .ZN(new_n541));
  NOR2_X1   g340(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n527), .B(new_n537), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n508), .B(KEYINPUT13), .Z(new_n544));
  AOI22_X1  g343(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n527), .B(KEYINPUT17), .ZN(new_n546));
  INV_X1    g345(.A(new_n537), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n542), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n548), .A2(new_n508), .A3(new_n538), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n507), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n545), .A2(new_n550), .A3(new_n507), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n501), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT100), .ZN(new_n557));
  XOR2_X1   g356(.A(G99gat), .B(G106gat), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT98), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G99gat), .ZN(new_n562));
  INV_X1    g361(.A(G106gat), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT8), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(KEYINPUT97), .B(G85gat), .Z(new_n565));
  OAI221_X1 g364(.A(new_n564), .B1(new_n565), .B2(G92gat), .C1(new_n559), .C2(KEYINPUT98), .ZN(new_n566));
  NOR2_X1   g365(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(G85gat), .B(G92gat), .C1(KEYINPUT96), .C2(KEYINPUT7), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n570), .A2(new_n571), .B1(KEYINPUT96), .B2(KEYINPUT7), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n561), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n566), .A2(new_n572), .A3(new_n561), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT99), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n578), .A3(new_n573), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n576), .A2(new_n579), .B1(new_n520), .B2(new_n526), .ZN(new_n580));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT41), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n557), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NOR3_X1   g383(.A1(new_n574), .A2(KEYINPUT99), .A3(new_n575), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n578), .B1(new_n577), .B2(new_n573), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n527), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n583), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(KEYINPUT100), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n546), .A2(new_n576), .A3(new_n579), .ZN(new_n591));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n590), .B2(new_n591), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT101), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n599), .A3(new_n594), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n582), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  OAI211_X1 g404(.A(KEYINPUT101), .B(new_n605), .C1(new_n595), .C2(new_n596), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G57gat), .B(G64gat), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT9), .ZN(new_n609));
  XNOR2_X1  g408(.A(G71gat), .B(G78gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n613), .A2(KEYINPUT94), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(KEYINPUT94), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n610), .B(new_n608), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G127gat), .B(G155gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G183gat), .B(G211gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n617), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n537), .B1(new_n628), .B2(KEYINPUT21), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT95), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n627), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n607), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT102), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n628), .B1(new_n574), .B2(new_n575), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n577), .A2(new_n617), .A3(new_n573), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n628), .A2(KEYINPUT10), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n576), .B2(new_n579), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n635), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n642), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n642), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g450(.A(KEYINPUT103), .B(new_n635), .C1(new_n639), .C2(new_n641), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n643), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n649), .B1(new_n653), .B2(new_n648), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n632), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n556), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n447), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g458(.A(G8gat), .B1(new_n656), .B2(new_n482), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT42), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT16), .B(G8gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT104), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n656), .A2(new_n482), .A3(new_n663), .ZN(new_n664));
  MUX2_X1   g463(.A(new_n661), .B(KEYINPUT42), .S(new_n664), .Z(G1325gat));
  NAND2_X1  g464(.A1(new_n493), .A2(new_n495), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(G15gat), .B1(new_n656), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n492), .ZN(new_n669));
  INV_X1    g468(.A(G15gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n668), .B1(new_n656), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT105), .ZN(G1326gat));
  NAND2_X1  g472(.A1(new_n488), .A2(new_n490), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n656), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  INV_X1    g476(.A(new_n631), .ZN(new_n678));
  INV_X1    g477(.A(new_n654), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n607), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n556), .A2(new_n517), .A3(new_n447), .A4(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT45), .Z(new_n683));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684));
  INV_X1    g483(.A(new_n553), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n685), .B2(new_n551), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n552), .A2(KEYINPUT106), .A3(new_n553), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n446), .A2(KEYINPUT107), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n472), .B2(new_n483), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n441), .A2(new_n694), .A3(new_n445), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n691), .A2(new_n693), .A3(new_n698), .A4(new_n695), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n607), .A2(KEYINPUT44), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n501), .B2(new_n607), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n690), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n517), .B1(new_n703), .B2(new_n447), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n683), .A2(new_n704), .ZN(G1328gat));
  AND2_X1   g504(.A1(new_n484), .A2(new_n500), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n554), .B(new_n681), .C1(new_n706), .C2(new_n446), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n482), .A2(G36gat), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT109), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n556), .A2(new_n712), .A3(new_n681), .A4(new_n708), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n482), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n518), .B1(new_n703), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n711), .B1(new_n710), .B2(new_n713), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n716), .A2(new_n720), .ZN(G1329gat));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  INV_X1    g521(.A(G43gat), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n703), .B2(new_n666), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n707), .A2(G43gat), .A3(new_n492), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n701), .A2(new_n702), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n666), .A3(new_n689), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT111), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n703), .A2(new_n730), .A3(new_n666), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n723), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n725), .A2(new_n722), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n726), .B1(new_n732), .B2(new_n733), .ZN(G1330gat));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735));
  INV_X1    g534(.A(G50gat), .ZN(new_n736));
  INV_X1    g535(.A(new_n674), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n703), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n674), .A2(G50gat), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n707), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n735), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743));
  INV_X1    g542(.A(new_n368), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n744), .A3(new_n689), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT48), .B1(new_n707), .B2(new_n740), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n743), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  AOI211_X1 g548(.A(KEYINPUT112), .B(new_n747), .C1(new_n745), .C2(G50gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n742), .B1(new_n749), .B2(new_n750), .ZN(G1331gat));
  AND2_X1   g550(.A1(new_n697), .A2(new_n699), .ZN(new_n752));
  INV_X1    g551(.A(new_n688), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n632), .A2(new_n679), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n447), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  INV_X1    g557(.A(KEYINPUT49), .ZN(new_n759));
  INV_X1    g558(.A(G64gat), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n756), .B(new_n717), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1333gat));
  INV_X1    g562(.A(G71gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n756), .A2(new_n764), .A3(new_n669), .ZN(new_n765));
  OAI21_X1  g564(.A(G71gat), .B1(new_n755), .B2(new_n667), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(KEYINPUT50), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1334gat));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n737), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g572(.A1(new_n678), .A2(new_n654), .A3(new_n688), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n701), .B2(new_n702), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(KEYINPUT113), .A3(new_n447), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT113), .B1(new_n775), .B2(new_n447), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n565), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n607), .A2(new_n631), .A3(new_n753), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n696), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT114), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n696), .A2(new_n783), .A3(KEYINPUT51), .A4(new_n779), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT51), .B1(new_n696), .B2(new_n779), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n654), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n438), .A2(new_n565), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n778), .B1(new_n787), .B2(new_n788), .ZN(G1336gat));
  INV_X1    g588(.A(new_n774), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n727), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G92gat), .B1(new_n791), .B2(new_n482), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n717), .A2(new_n569), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n792), .B(new_n793), .C1(new_n787), .C2(new_n794), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n782), .A2(new_n784), .B1(new_n781), .B2(new_n780), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n796), .A2(new_n679), .A3(new_n794), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n569), .B1(new_n775), .B2(new_n717), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT52), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n791), .B2(new_n667), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n669), .A2(new_n562), .A3(new_n654), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT115), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n796), .B2(new_n803), .ZN(G1338gat));
  OAI21_X1  g603(.A(G106gat), .B1(new_n791), .B2(new_n368), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n744), .A2(new_n563), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n805), .B(new_n806), .C1(new_n787), .C2(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n796), .A2(new_n679), .A3(new_n807), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n563), .B1(new_n775), .B2(new_n737), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT53), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(G1339gat));
  AOI21_X1  g611(.A(new_n508), .B1(new_n548), .B2(new_n538), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n543), .A2(new_n544), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n505), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n654), .A2(new_n553), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n651), .A2(new_n652), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n585), .A2(new_n586), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n634), .B(new_n821), .C1(new_n822), .C2(new_n640), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n642), .A2(new_n823), .A3(KEYINPUT54), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n647), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n817), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n647), .A4(new_n824), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n649), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n816), .B1(new_n688), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(KEYINPUT117), .B(new_n816), .C1(new_n688), .C2(new_n828), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n607), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n607), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n553), .A2(new_n815), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT116), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n828), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n631), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n632), .A2(new_n654), .A3(new_n753), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n737), .A2(new_n492), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n717), .A2(new_n438), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n841), .A2(new_n554), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n844), .A2(new_n845), .A3(G113gat), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n844), .B2(G113gat), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n841), .A2(new_n843), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n370), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n753), .A2(new_n212), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n846), .A2(new_n847), .B1(new_n849), .B2(new_n850), .ZN(G1340gat));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n842), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n852), .A2(new_n210), .A3(new_n679), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n848), .A2(new_n370), .A3(new_n654), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n210), .B2(new_n854), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n852), .B2(new_n678), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n631), .A2(new_n205), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n849), .B2(new_n857), .ZN(G1342gat));
  NOR2_X1   g657(.A1(new_n444), .A2(G134gat), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n841), .A2(new_n834), .A3(new_n843), .A4(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n860), .A2(new_n861), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT56), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n860), .A2(new_n861), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n862), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n841), .A2(new_n834), .A3(new_n842), .A4(new_n843), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G134gat), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT120), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n869), .A2(new_n872), .A3(G134gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n865), .A2(new_n868), .A3(new_n874), .ZN(G1343gat));
  NAND2_X1  g674(.A1(new_n667), .A2(new_n843), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n554), .A2(new_n826), .A3(new_n649), .A4(new_n827), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n816), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n607), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n631), .B1(new_n838), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n737), .B1(new_n880), .B2(new_n840), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n881), .B2(KEYINPUT57), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n883), .B(new_n744), .C1(new_n839), .C2(new_n840), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n884), .A3(new_n554), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT121), .A4(new_n554), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(G141gat), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n666), .A2(new_n368), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n555), .A2(G141gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n848), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n882), .A2(new_n884), .ZN(new_n895));
  OAI21_X1  g694(.A(G141gat), .B1(new_n895), .B2(new_n688), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT58), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n894), .A2(new_n898), .ZN(G1344gat));
  XOR2_X1   g698(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n900));
  NAND2_X1  g699(.A1(new_n655), .A2(new_n555), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n607), .A2(new_n836), .A3(new_n828), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n877), .A2(new_n816), .B1(new_n604), .B2(new_n606), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n678), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n674), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT123), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT57), .B(new_n744), .C1(new_n839), .C2(new_n840), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n632), .A2(new_n554), .A3(new_n654), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n737), .B1(new_n880), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n910), .A3(new_n883), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n906), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n912), .A2(new_n667), .A3(new_n654), .A4(new_n843), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n900), .B1(new_n913), .B2(G148gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n895), .A2(new_n679), .ZN(new_n915));
  INV_X1    g714(.A(G148gat), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n915), .A2(KEYINPUT59), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n848), .A2(new_n891), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n654), .A2(new_n916), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n914), .A2(new_n917), .B1(new_n918), .B2(new_n919), .ZN(G1345gat));
  OAI21_X1  g719(.A(G155gat), .B1(new_n895), .B2(new_n678), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n678), .A2(G155gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n918), .B2(new_n922), .ZN(G1346gat));
  NAND2_X1  g722(.A1(new_n848), .A2(new_n834), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925));
  INV_X1    g724(.A(G162gat), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n891), .A2(new_n926), .ZN(new_n927));
  OR3_X1    g726(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G162gat), .B1(new_n895), .B2(new_n607), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n925), .B1(new_n924), .B2(new_n927), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n482), .A2(new_n447), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n841), .A2(new_n370), .A3(new_n753), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n219), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n841), .A2(new_n932), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n842), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n555), .A2(new_n219), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT125), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n941), .B(new_n934), .C1(new_n936), .C2(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1348gat));
  OAI21_X1  g742(.A(G176gat), .B1(new_n936), .B2(new_n679), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n935), .A2(new_n370), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n654), .A2(new_n220), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1349gat));
  NAND4_X1  g746(.A1(new_n841), .A2(new_n631), .A3(new_n842), .A4(new_n932), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G183gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n631), .A2(new_n251), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT60), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT60), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n953), .B(new_n949), .C1(new_n945), .C2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1350gat));
  NAND4_X1  g754(.A1(new_n841), .A2(new_n834), .A3(new_n842), .A4(new_n932), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n956), .A2(new_n957), .A3(G190gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n956), .B2(G190gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n834), .A2(new_n248), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n958), .A2(new_n959), .B1(new_n945), .B2(new_n960), .ZN(G1351gat));
  NOR3_X1   g760(.A1(new_n666), .A2(new_n447), .A3(new_n482), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n912), .A2(new_n554), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n912), .A2(new_n965), .A3(new_n554), .A4(new_n962), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n964), .A2(G197gat), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n841), .A2(new_n891), .A3(new_n932), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n969), .A2(new_n316), .A3(new_n753), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n967), .A2(new_n971), .ZN(G1352gat));
  NOR2_X1   g771(.A1(new_n679), .A2(G204gat), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n841), .A2(new_n891), .A3(new_n932), .A4(new_n973), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT62), .Z(new_n975));
  AND3_X1   g774(.A1(new_n912), .A2(new_n654), .A3(new_n962), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n314), .B2(new_n976), .ZN(G1353gat));
  NOR2_X1   g776(.A1(new_n678), .A2(G211gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n969), .A2(new_n970), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n912), .A2(new_n631), .A3(new_n962), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  NOR2_X1   g782(.A1(new_n607), .A2(G218gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n970), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n912), .A2(new_n834), .A3(new_n962), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(G218gat), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(new_n987), .ZN(G1355gat));
endmodule


