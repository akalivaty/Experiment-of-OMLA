//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(G1gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n211), .B2(KEYINPUT91), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT16), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n213), .B2(G1gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n212), .B(new_n215), .Z(new_n216));
  XOR2_X1   g015(.A(G43gat), .B(G50gat), .Z(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n218), .B2(KEYINPUT14), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n219), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n217), .B1(new_n223), .B2(KEYINPUT15), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(KEYINPUT15), .B2(new_n223), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(KEYINPUT15), .A3(new_n217), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n216), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n226), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n216), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(KEYINPUT17), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n228), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT92), .Z(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n216), .B(new_n227), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n236), .B(KEYINPUT13), .Z(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT93), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT93), .B1(new_n238), .B2(new_n239), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n237), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT18), .B1(new_n234), .B2(new_n236), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n208), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n240), .B(new_n241), .ZN(new_n247));
  INV_X1    g046(.A(new_n245), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n237), .A4(new_n207), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(G211gat), .B(G218gat), .Z(new_n252));
  XNOR2_X1  g051(.A(G197gat), .B(G204gat), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT74), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT74), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(new_n258), .A3(new_n255), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n252), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n252), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT77), .ZN(new_n265));
  INV_X1    g064(.A(G148gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(G141gat), .ZN(new_n267));
  INV_X1    g066(.A(G141gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n268), .A2(G148gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n265), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(G148gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(G141gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT77), .ZN(new_n273));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT2), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n270), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n274), .ZN(new_n277));
  NOR2_X1   g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT78), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(new_n268), .A3(G148gat), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n281), .B(new_n275), .C1(new_n277), .C2(new_n278), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G141gat), .B(G148gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT78), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n276), .A2(new_n279), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT3), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT29), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n264), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(new_n260), .B2(new_n262), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n286), .B1(new_n291), .B2(new_n287), .ZN(new_n292));
  INV_X1    g091(.A(G228gat), .ZN(new_n293));
  INV_X1    g092(.A(G233gat), .ZN(new_n294));
  OAI22_X1  g093(.A1(new_n289), .A2(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n293), .A2(new_n294), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT84), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n263), .B1(new_n288), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n275), .B1(new_n284), .B2(KEYINPUT77), .ZN(new_n299));
  INV_X1    g098(.A(new_n273), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n279), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n285), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n297), .B(new_n290), .C1(new_n303), .C2(KEYINPUT3), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n296), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT3), .B1(new_n291), .B2(KEYINPUT83), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT83), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n308), .B(new_n290), .C1(new_n260), .C2(new_n262), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n286), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n295), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G22gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT85), .ZN(new_n313));
  INV_X1    g112(.A(new_n252), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n253), .A2(new_n258), .A3(new_n255), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n258), .B1(new_n253), .B2(new_n255), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n317), .B2(new_n261), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n287), .B1(new_n318), .B2(new_n308), .ZN(new_n319));
  INV_X1    g118(.A(new_n309), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n303), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n301), .A2(new_n302), .A3(new_n287), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT84), .B1(new_n322), .B2(KEYINPUT29), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(new_n263), .A3(new_n304), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n324), .A3(new_n296), .ZN(new_n325));
  INV_X1    g124(.A(G22gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n295), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n313), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT86), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT86), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n312), .A2(new_n313), .A3(new_n330), .A4(new_n327), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G78gat), .B(G106gat), .ZN(new_n333));
  INV_X1    g132(.A(G50gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT82), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n336), .B(KEYINPUT31), .Z(new_n337));
  AND3_X1   g136(.A1(new_n325), .A2(new_n326), .A3(new_n295), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n326), .B1(new_n325), .B2(new_n295), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n340), .B2(new_n313), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n337), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n312), .A2(new_n327), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(KEYINPUT85), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(new_n329), .A3(new_n331), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G226gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(new_n294), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT26), .ZN(new_n350));
  INV_X1    g149(.A(G169gat), .ZN(new_n351));
  INV_X1    g150(.A(G176gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  AND3_X1   g153(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n353), .B(new_n354), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT27), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(G183gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT27), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT68), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(G190gat), .B1(new_n364), .B2(KEYINPUT68), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n362), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n364), .A2(new_n366), .ZN(new_n372));
  INV_X1    g171(.A(G190gat), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n372), .A2(KEYINPUT28), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n360), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT65), .B(KEYINPUT25), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n377));
  AND2_X1   g176(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n358), .A2(new_n377), .B1(new_n378), .B2(G190gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT23), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT23), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(G169gat), .B2(G176gat), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n380), .B(new_n382), .C1(new_n355), .C2(new_n356), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT67), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT66), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n390), .A2(KEYINPUT67), .A3(new_n382), .A4(new_n380), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n376), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n383), .A2(new_n379), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n375), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n349), .B1(new_n395), .B2(new_n290), .ZN(new_n396));
  INV_X1    g195(.A(new_n349), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n383), .A2(new_n384), .ZN(new_n398));
  INV_X1    g197(.A(new_n379), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n391), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n376), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n394), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n397), .B1(new_n404), .B2(new_n375), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT75), .B1(new_n396), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n364), .A2(KEYINPUT68), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n373), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT68), .B1(new_n364), .B2(new_n366), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n361), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n372), .A2(KEYINPUT28), .A3(new_n373), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n359), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n412), .B1(new_n402), .B2(new_n403), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n397), .B1(new_n413), .B2(KEYINPUT29), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n406), .A2(new_n264), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n395), .A2(new_n349), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n263), .ZN(new_n420));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT30), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(KEYINPUT76), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n417), .A2(KEYINPUT30), .A3(new_n420), .A4(new_n423), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n417), .A2(new_n420), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n428), .B1(new_n429), .B2(new_n423), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT76), .B1(new_n424), .B2(new_n425), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G127gat), .B(G134gat), .ZN(new_n433));
  INV_X1    g232(.A(G113gat), .ZN(new_n434));
  INV_X1    g233(.A(G120gat), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT1), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(KEYINPUT70), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT70), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G113gat), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n435), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT1), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n442), .B1(G113gat), .B2(G120gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(G113gat), .A2(G120gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI22_X1  g245(.A1(new_n437), .A2(new_n441), .B1(new_n446), .B2(new_n433), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT71), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI221_X1 g248(.A(KEYINPUT71), .B1(new_n446), .B2(new_n433), .C1(new_n437), .C2(new_n441), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n404), .A2(new_n449), .A3(new_n450), .A4(new_n375), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n450), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n395), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n455), .B(KEYINPUT64), .Z(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT72), .B(KEYINPUT33), .Z(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XOR2_X1   g258(.A(G15gat), .B(G43gat), .Z(new_n460));
  XNOR2_X1  g259(.A(G71gat), .B(G99gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n456), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n451), .A2(new_n453), .A3(new_n465), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n466), .A2(KEYINPUT34), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(KEYINPUT34), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n457), .A2(KEYINPUT32), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n467), .A2(new_n468), .B1(KEYINPUT32), .B2(new_n457), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n470), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n467), .A2(KEYINPUT32), .A3(new_n457), .A4(new_n468), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n463), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n347), .A2(new_n432), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480));
  XOR2_X1   g279(.A(G1gat), .B(G29gat), .Z(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G57gat), .B(G85gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n487));
  INV_X1    g286(.A(G134gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G127gat), .ZN(new_n489));
  INV_X1    g288(.A(G127gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G134gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(new_n443), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n438), .A2(new_n440), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G120gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n436), .A2(new_n444), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n493), .A2(new_n495), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT79), .B1(new_n286), .B2(new_n497), .ZN(new_n498));
  AND4_X1   g297(.A1(KEYINPUT79), .A2(new_n301), .A3(new_n497), .A4(new_n302), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n487), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n286), .A2(new_n449), .A3(KEYINPUT4), .A4(new_n450), .ZN(new_n501));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n497), .B1(new_n303), .B2(KEYINPUT3), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(KEYINPUT3), .B2(new_n303), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  OAI22_X1  g305(.A1(new_n498), .A2(new_n499), .B1(new_n286), .B2(new_n497), .ZN(new_n507));
  INV_X1    g306(.A(new_n502), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n506), .A2(new_n509), .A3(KEYINPUT5), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT79), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n303), .B2(new_n447), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n286), .A2(KEYINPUT79), .A3(new_n497), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(KEYINPUT4), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n487), .B1(new_n452), .B2(new_n303), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n505), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  AOI211_X1 g316(.A(new_n480), .B(new_n486), .C1(new_n510), .C2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(KEYINPUT88), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n512), .A2(new_n513), .B1(new_n303), .B2(new_n447), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT5), .B1(new_n520), .B2(new_n502), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n447), .B1(new_n286), .B2(new_n287), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n502), .B(new_n501), .C1(new_n522), .C2(new_n322), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT4), .B1(new_n512), .B2(new_n513), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n517), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n485), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n486), .A3(new_n517), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n480), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(KEYINPUT6), .A3(new_n485), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n519), .B1(new_n531), .B2(KEYINPUT88), .ZN(new_n532));
  OR3_X1    g331(.A1(new_n479), .A2(KEYINPUT35), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n423), .B1(new_n417), .B2(new_n420), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n417), .A2(new_n420), .A3(new_n423), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(KEYINPUT30), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n424), .A2(new_n425), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n531), .A2(new_n536), .A3(new_n539), .A4(new_n426), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT81), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n430), .A2(new_n431), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n543), .A2(KEYINPUT81), .A3(new_n531), .A4(new_n426), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n347), .A2(new_n542), .A3(new_n544), .A4(new_n478), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n545), .A2(KEYINPUT89), .A3(KEYINPUT35), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT89), .B1(new_n545), .B2(KEYINPUT35), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n533), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT36), .B1(new_n477), .B2(KEYINPUT73), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT73), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT36), .ZN(new_n551));
  AOI211_X1 g350(.A(new_n550), .B(new_n551), .C1(new_n473), .C2(new_n476), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n530), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT6), .B1(new_n526), .B2(new_n485), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n518), .B1(new_n528), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n424), .B(new_n555), .C1(new_n557), .C2(new_n554), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT38), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n417), .A2(new_n560), .A3(new_n420), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT87), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT87), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n417), .A2(new_n563), .A3(new_n560), .A4(new_n420), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n423), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n429), .A2(new_n560), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n559), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n406), .A2(new_n263), .A3(new_n416), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n560), .B1(new_n419), .B2(new_n264), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n559), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n423), .B(new_n571), .C1(new_n562), .C2(new_n564), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n558), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n345), .A2(new_n329), .A3(new_n331), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n344), .A2(KEYINPUT85), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n329), .A2(new_n331), .B1(new_n575), .B2(new_n337), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT40), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n505), .A2(new_n515), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n502), .B1(new_n578), .B2(new_n514), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT39), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n486), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT39), .B1(new_n507), .B2(new_n508), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n577), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n485), .B1(new_n579), .B2(new_n580), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n586), .B(KEYINPUT40), .C1(new_n579), .C2(new_n583), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n587), .A3(new_n527), .ZN(new_n588));
  OAI22_X1  g387(.A1(new_n574), .A2(new_n576), .B1(new_n432), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n553), .B1(new_n573), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n347), .B1(new_n542), .B2(new_n544), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n251), .B1(new_n548), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(KEYINPUT9), .ZN(new_n595));
  XNOR2_X1  g394(.A(G57gat), .B(G64gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n594), .A2(KEYINPUT94), .ZN(new_n600));
  OR3_X1    g399(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n599), .B1(new_n597), .B2(new_n600), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n603), .B(KEYINPUT96), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT21), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n216), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(KEYINPUT21), .ZN(new_n607));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT95), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n610), .B(new_n616), .Z(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT7), .ZN(new_n619));
  NAND2_X1  g418(.A1(G99gat), .A2(G106gat), .ZN(new_n620));
  INV_X1    g419(.A(G85gat), .ZN(new_n621));
  INV_X1    g420(.A(G92gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(KEYINPUT8), .A2(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G99gat), .B(G106gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  NAND3_X1  g425(.A1(new_n233), .A2(new_n231), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  AND2_X1   g427(.A1(G232gat), .A2(G233gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n628), .A2(new_n229), .B1(KEYINPUT41), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G190gat), .B(G218gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n634));
  XOR2_X1   g433(.A(G134gat), .B(G162gat), .Z(new_n635));
  NOR2_X1   g434(.A1(new_n629), .A2(KEYINPUT41), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  OR3_X1    g436(.A1(new_n633), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(KEYINPUT97), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n617), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n628), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n626), .B(new_n603), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n644), .A2(KEYINPUT98), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT98), .B1(new_n644), .B2(new_n645), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(G230gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n294), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n651), .B2(new_n644), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n642), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n593), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT99), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n593), .A2(KEYINPUT99), .A3(new_n660), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n557), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  INV_X1    g465(.A(new_n432), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT16), .B(G8gat), .Z(new_n668));
  AND3_X1   g467(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n209), .B1(new_n664), .B2(new_n667), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT42), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(KEYINPUT42), .B2(new_n669), .ZN(G1325gat));
  INV_X1    g471(.A(G15gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n664), .A2(new_n673), .A3(new_n478), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n553), .B1(new_n662), .B2(new_n663), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n675), .B2(new_n673), .ZN(G1326gat));
  INV_X1    g475(.A(new_n347), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n664), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NAND2_X1  g479(.A1(new_n548), .A2(new_n592), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n641), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n659), .A2(new_n617), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n250), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n246), .A2(new_n249), .A3(KEYINPUT101), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n542), .A2(new_n544), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n692), .A2(new_n677), .A3(KEYINPUT102), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT102), .B1(new_n692), .B2(new_n677), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n693), .A2(new_n590), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n548), .B2(KEYINPUT103), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n479), .A2(KEYINPUT35), .A3(new_n532), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n478), .B1(new_n574), .B2(new_n576), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT35), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT89), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n545), .A2(KEYINPUT89), .A3(KEYINPUT35), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n641), .B1(new_n696), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n684), .B(new_n691), .C1(new_n706), .C2(KEYINPUT44), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT104), .B1(new_n707), .B2(new_n531), .ZN(new_n708));
  INV_X1    g507(.A(new_n684), .ZN(new_n709));
  INV_X1    g508(.A(new_n641), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n590), .A2(new_n694), .ZN(new_n711));
  INV_X1    g510(.A(new_n693), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n703), .B2(new_n704), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n548), .A2(KEYINPUT103), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n710), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n709), .B1(new_n716), .B2(new_n682), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n717), .A2(new_n718), .A3(new_n557), .A4(new_n691), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n708), .A2(G29gat), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n686), .A2(new_n641), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n681), .A2(new_n250), .A3(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n722), .A2(G29gat), .A3(new_n531), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT100), .B(KEYINPUT45), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT105), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n720), .A2(new_n728), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1328gat));
  OAI21_X1  g529(.A(G36gat), .B1(new_n707), .B2(new_n432), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n667), .A2(new_n221), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n722), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT106), .Z(G1329gat));
  INV_X1    g535(.A(new_n553), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G43gat), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n477), .ZN(new_n739));
  OAI22_X1  g538(.A1(new_n707), .A2(new_n738), .B1(G43gat), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1330gat));
  OAI21_X1  g541(.A(G50gat), .B1(new_n707), .B2(new_n347), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n677), .A2(new_n334), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n743), .B(KEYINPUT48), .C1(new_n722), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n722), .A2(new_n744), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT108), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT48), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(KEYINPUT109), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n750), .B(KEYINPUT48), .C1(new_n743), .C2(new_n747), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n745), .B1(new_n749), .B2(new_n751), .ZN(G1331gat));
  NAND4_X1  g551(.A1(new_n690), .A2(new_n617), .A3(new_n641), .A4(new_n659), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n696), .B2(new_n705), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n557), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT110), .B(G57gat), .Z(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1332gat));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n758));
  INV_X1    g557(.A(G64gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n667), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT111), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n759), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1333gat));
  INV_X1    g563(.A(G71gat), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n754), .A2(new_n765), .A3(new_n478), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n754), .A2(new_n737), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n765), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n677), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  INV_X1    g570(.A(new_n617), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n690), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT112), .Z(new_n774));
  NOR3_X1   g573(.A1(new_n716), .A2(KEYINPUT51), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  INV_X1    g575(.A(new_n774), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n706), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n659), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n775), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n621), .A3(new_n557), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n774), .A2(new_n779), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n684), .B(new_n782), .C1(new_n706), .C2(KEYINPUT44), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n716), .A2(new_n682), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n786), .A2(KEYINPUT113), .A3(new_n684), .A4(new_n782), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n785), .A2(new_n557), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n781), .B1(new_n788), .B2(new_n621), .ZN(G1336gat));
  NAND3_X1  g588(.A1(new_n785), .A2(new_n667), .A3(new_n787), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n432), .A2(G92gat), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n790), .A2(G92gat), .B1(new_n780), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n780), .A2(new_n791), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n793), .ZN(new_n795));
  INV_X1    g594(.A(new_n783), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n622), .B1(new_n796), .B2(new_n667), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n792), .A2(new_n793), .B1(new_n795), .B2(new_n797), .ZN(G1337gat));
  INV_X1    g597(.A(G99gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n799), .A3(new_n478), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n737), .A3(new_n787), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G99gat), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n800), .B1(new_n804), .B2(new_n805), .ZN(G1338gat));
  NAND3_X1  g605(.A1(new_n785), .A2(new_n677), .A3(new_n787), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n347), .A2(G106gat), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n807), .A2(G106gat), .B1(new_n780), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n780), .A2(new_n808), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n810), .ZN(new_n812));
  INV_X1    g611(.A(G106gat), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n796), .B2(new_n677), .ZN(new_n814));
  OAI22_X1  g613(.A1(new_n809), .A2(new_n810), .B1(new_n812), .B2(new_n814), .ZN(G1339gat));
  NAND2_X1  g614(.A1(new_n660), .A2(new_n690), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n234), .A2(new_n236), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n238), .A2(new_n239), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n206), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n659), .A2(new_n249), .A3(new_n820), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n652), .A2(KEYINPUT54), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n650), .B(new_n643), .C1(new_n646), .C2(new_n647), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n652), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n656), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n656), .A4(new_n824), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n657), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n821), .B1(new_n829), .B2(new_n690), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n641), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n249), .A2(new_n820), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT115), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n827), .A2(new_n710), .A3(new_n657), .A4(new_n828), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n817), .B1(new_n837), .B2(new_n772), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n531), .A3(new_n479), .ZN(new_n839));
  INV_X1    g638(.A(new_n690), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n839), .A2(new_n438), .A3(new_n440), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n667), .A2(new_n531), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n838), .A2(KEYINPUT116), .A3(new_n677), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n835), .B1(new_n641), .B2(new_n830), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n816), .B1(new_n845), .B2(new_n617), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n846), .B2(new_n347), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n478), .B(new_n842), .C1(new_n843), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT117), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT116), .B1(new_n838), .B2(new_n677), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n846), .A2(new_n844), .A3(new_n347), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n478), .A4(new_n842), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n849), .A2(new_n250), .A3(new_n854), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n855), .A2(KEYINPUT118), .A3(G113gat), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT118), .B1(new_n855), .B2(G113gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n841), .B1(new_n856), .B2(new_n857), .ZN(G1340gat));
  AND4_X1   g657(.A1(G120gat), .A2(new_n849), .A3(new_n659), .A4(new_n854), .ZN(new_n859));
  AOI21_X1  g658(.A(G120gat), .B1(new_n839), .B2(new_n659), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(G1341gat));
  NAND3_X1  g660(.A1(new_n839), .A2(new_n490), .A3(new_n617), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n849), .A2(new_n617), .A3(new_n854), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n490), .ZN(G1342gat));
  NAND3_X1  g663(.A1(new_n839), .A2(new_n488), .A3(new_n710), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT56), .Z(new_n866));
  AND3_X1   g665(.A1(new_n849), .A2(new_n710), .A3(new_n854), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n488), .ZN(G1343gat));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n553), .A2(new_n842), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n827), .A2(new_n250), .A3(new_n657), .A4(new_n828), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n710), .B1(new_n872), .B2(new_n821), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n772), .B1(new_n873), .B2(new_n835), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n816), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(KEYINPUT57), .A3(new_n677), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n846), .B2(new_n677), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(KEYINPUT119), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n879), .B(KEYINPUT57), .C1(new_n846), .C2(new_n677), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n871), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n869), .B1(new_n881), .B2(new_n251), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n838), .B2(new_n347), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n879), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n877), .A2(KEYINPUT119), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(new_n876), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n887), .A2(KEYINPUT120), .A3(new_n250), .A4(new_n871), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(G141gat), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n846), .A2(new_n557), .ZN(new_n890));
  NOR4_X1   g689(.A1(new_n890), .A2(new_n667), .A3(new_n347), .A4(new_n737), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n268), .A3(new_n250), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G141gat), .B1(new_n881), .B2(new_n690), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n892), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT58), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(G1344gat));
  NAND3_X1  g698(.A1(new_n891), .A2(new_n266), .A3(new_n659), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n660), .A2(new_n251), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n874), .A2(KEYINPUT121), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n677), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT121), .B1(new_n874), .B2(new_n902), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n883), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n846), .A2(KEYINPUT57), .A3(new_n677), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n779), .B(new_n870), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n266), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n779), .B1(new_n906), .B2(new_n907), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT122), .B1(new_n912), .B2(new_n870), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n901), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n881), .A2(new_n779), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(KEYINPUT59), .A3(new_n266), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n900), .B1(new_n914), .B2(new_n916), .ZN(G1345gat));
  OAI21_X1  g716(.A(G155gat), .B1(new_n881), .B2(new_n772), .ZN(new_n918));
  INV_X1    g717(.A(G155gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n891), .A2(new_n919), .A3(new_n617), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n881), .B2(new_n641), .ZN(new_n922));
  INV_X1    g721(.A(G162gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n891), .A2(new_n923), .A3(new_n710), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n432), .A2(new_n557), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n478), .B(new_n926), .C1(new_n843), .C2(new_n847), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(new_n351), .A3(new_n251), .ZN(new_n928));
  NOR4_X1   g727(.A1(new_n838), .A2(new_n557), .A3(new_n432), .A4(new_n698), .ZN(new_n929));
  AOI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n840), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n928), .A2(new_n930), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n927), .B2(new_n779), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n929), .A2(new_n352), .A3(new_n659), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1349gat));
  OAI21_X1  g733(.A(G183gat), .B1(new_n927), .B2(new_n772), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n929), .A2(new_n372), .A3(new_n617), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  OAI221_X1 g738(.A(G190gat), .B1(KEYINPUT123), .B2(new_n939), .C1(new_n927), .C2(new_n641), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n939), .A2(KEYINPUT123), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n929), .A2(new_n373), .A3(new_n710), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(G1351gat));
  NOR2_X1   g744(.A1(new_n838), .A2(new_n557), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n737), .A2(new_n432), .A3(new_n347), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n840), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n553), .A2(new_n926), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n951), .B1(new_n906), .B2(new_n907), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n250), .A2(G197gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(G1352gat));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  XOR2_X1   g754(.A(KEYINPUT124), .B(G204gat), .Z(new_n956));
  NAND4_X1  g755(.A1(new_n946), .A2(new_n659), .A3(new_n947), .A4(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n957), .B2(new_n959), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n951), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n956), .B1(new_n911), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n955), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n961), .A2(new_n962), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n912), .A2(new_n951), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n967), .B(KEYINPUT126), .C1(new_n968), .C2(new_n956), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n966), .A2(new_n969), .ZN(G1353gat));
  OR3_X1    g769(.A1(new_n948), .A2(G211gat), .A3(new_n772), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n952), .A2(new_n617), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  INV_X1    g774(.A(G218gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n949), .A2(new_n976), .A3(new_n710), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n952), .A2(new_n710), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(new_n976), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n981), .B(new_n977), .C1(new_n978), .C2(new_n976), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1355gat));
endmodule


