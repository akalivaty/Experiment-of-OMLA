//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n537,
    new_n538, new_n539, new_n540, new_n542, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n587, new_n588,
    new_n591, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1109, new_n1110, new_n1111;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n462), .A2(new_n466), .ZN(G160));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n463), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n472), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  NAND3_X1  g055(.A1(new_n469), .A2(new_n471), .A3(G126), .ZN(new_n481));
  NAND2_X1  g056(.A1(G114), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n469), .A2(new_n471), .A3(G138), .A4(new_n463), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n483), .A2(G2105), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT68), .A2(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(G138), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n492), .B2(new_n472), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(new_n463), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  NAND2_X1  g071(.A1(G75), .A2(G543), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G62), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(new_n498), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n504), .A2(G651), .B1(new_n508), .B2(G50), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n511), .B1(new_n502), .B2(new_n507), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n513), .B(KEYINPUT69), .C1(new_n506), .C2(new_n505), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n509), .B1(new_n510), .B2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  AND3_X1   g092(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XOR2_X1   g094(.A(new_n519), .B(KEYINPUT7), .Z(new_n520));
  AOI211_X1 g095(.A(new_n518), .B(new_n520), .C1(G51), .C2(new_n508), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n512), .A2(new_n514), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(G286));
  INV_X1    g099(.A(G286), .ZN(G168));
  AOI22_X1  g100(.A1(new_n522), .A2(G90), .B1(G52), .B2(new_n508), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT70), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n527), .A2(KEYINPUT71), .A3(new_n530), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  NAND2_X1  g111(.A1(new_n508), .A2(G43), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n529), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n522), .B2(G81), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  AND3_X1   g116(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G36), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G188));
  NAND3_X1  g121(.A1(new_n508), .A2(KEYINPUT72), .A3(G53), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT9), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n529), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n522), .A2(G91), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(G299));
  NAND2_X1  g128(.A1(new_n508), .A2(G49), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G87), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT73), .B1(new_n515), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n512), .A2(new_n514), .A3(new_n558), .A4(G87), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n555), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(G288));
  NAND2_X1  g137(.A1(new_n522), .A2(G86), .ZN(new_n563));
  NAND2_X1  g138(.A1(G73), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G61), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n502), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(new_n508), .B2(G48), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G305));
  AOI22_X1  g143(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n529), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT74), .Z(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(G47), .B2(new_n508), .ZN(new_n572));
  XNOR2_X1  g147(.A(KEYINPUT75), .B(G85), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n522), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(new_n522), .A2(G92), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT10), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n508), .A2(G54), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n529), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G868), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n584), .B1(G171), .B2(new_n583), .ZN(G284));
  OAI21_X1  g160(.A(new_n584), .B1(G171), .B2(new_n583), .ZN(G321));
  NAND2_X1  g161(.A1(G286), .A2(G868), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n552), .B(KEYINPUT76), .Z(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n588), .B2(G868), .ZN(G280));
  XNOR2_X1  g164(.A(G280), .B(KEYINPUT77), .ZN(G297));
  AND3_X1   g165(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n591));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G860), .ZN(G148));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g172(.A1(new_n475), .A2(G2104), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT12), .Z(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT13), .Z(new_n600));
  NOR2_X1   g175(.A1(KEYINPUT78), .A2(G2100), .ZN(new_n601));
  AND2_X1   g176(.A1(KEYINPUT78), .A2(G2100), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n473), .A2(G123), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n475), .A2(G135), .ZN(new_n605));
  NOR2_X1   g180(.A1(G99), .A2(G2105), .ZN(new_n606));
  OAI21_X1  g181(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n604), .B(new_n605), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(G2096), .Z(new_n609));
  OAI211_X1 g184(.A(new_n603), .B(new_n609), .C1(new_n600), .C2(new_n601), .ZN(G156));
  XNOR2_X1  g185(.A(G2451), .B(G2454), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT16), .ZN(new_n612));
  XOR2_X1   g187(.A(G2443), .B(G2446), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(G1341), .B(G1348), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT80), .B(G2438), .ZN(new_n617));
  XNOR2_X1  g192(.A(G2427), .B(G2430), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT15), .B(G2435), .Z(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(KEYINPUT79), .A2(KEYINPUT14), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n620), .A2(new_n621), .ZN(new_n624));
  OR2_X1    g199(.A1(KEYINPUT79), .A2(KEYINPUT14), .ZN(new_n625));
  NAND4_X1  g200(.A1(new_n622), .A2(new_n623), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n616), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G14), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(G401));
  INV_X1    g204(.A(KEYINPUT18), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2067), .B(G2678), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT81), .Z(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  AND2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(KEYINPUT17), .B1(new_n633), .B2(new_n634), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n630), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2072), .B(G2078), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n630), .B2(new_n635), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT82), .B(G2096), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(G227));
  XNOR2_X1  g218(.A(G1971), .B(G1976), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1956), .B(G2474), .Z(new_n648));
  XOR2_X1   g223(.A(G1961), .B(G1966), .Z(new_n649));
  AND2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n648), .A2(new_n649), .ZN(new_n653));
  AOI22_X1  g228(.A1(new_n651), .A2(new_n652), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  OR3_X1    g229(.A1(new_n647), .A2(new_n650), .A3(new_n653), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n654), .B(new_n655), .C1(new_n651), .C2(new_n652), .ZN(new_n656));
  XOR2_X1   g231(.A(G1991), .B(G1996), .Z(new_n657));
  XNOR2_X1  g232(.A(G1981), .B(G1986), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(G229));
  INV_X1    g238(.A(G16), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G22), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(G166), .B2(new_n664), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT89), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G1971), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(G23), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n560), .A2(KEYINPUT88), .A3(new_n561), .ZN(new_n670));
  AOI21_X1  g245(.A(KEYINPUT88), .B1(new_n560), .B2(new_n561), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n669), .B1(new_n672), .B2(new_n664), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT33), .B(G1976), .Z(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n664), .A2(G6), .ZN(new_n676));
  INV_X1    g251(.A(G305), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n677), .B2(new_n664), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT32), .B(G1981), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  NAND4_X1  g256(.A1(new_n668), .A2(new_n675), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(KEYINPUT34), .ZN(new_n683));
  AOI22_X1  g258(.A1(G119), .A2(new_n473), .B1(new_n475), .B2(G131), .ZN(new_n684));
  OR3_X1    g259(.A1(KEYINPUT86), .A2(G95), .A3(G2105), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n463), .A2(G107), .ZN(new_n686));
  OAI21_X1  g261(.A(KEYINPUT86), .B1(G95), .B2(G2105), .ZN(new_n687));
  NAND4_X1  g262(.A1(new_n685), .A2(new_n686), .A3(G2104), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  MUX2_X1   g264(.A(G25), .B(new_n689), .S(G29), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT35), .B(G1991), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n664), .A2(G24), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G290), .B2(G16), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT87), .B(G1986), .Z(new_n695));
  AOI22_X1  g270(.A1(new_n694), .A2(new_n695), .B1(new_n691), .B2(new_n690), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n694), .B2(new_n695), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n682), .B2(KEYINPUT34), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n683), .A2(new_n692), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT36), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT36), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n683), .A2(new_n698), .A3(new_n701), .A4(new_n692), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G26), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n473), .A2(G128), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n475), .A2(G140), .ZN(new_n707));
  OR2_X1    g282(.A1(G104), .A2(G2105), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n708), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(new_n704), .ZN(new_n712));
  MUX2_X1   g287(.A(new_n705), .B(new_n712), .S(KEYINPUT28), .Z(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(G2067), .ZN(new_n714));
  NOR2_X1   g289(.A1(G5), .A2(G16), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G171), .B2(G16), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1961), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT92), .B(KEYINPUT23), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n664), .A2(G20), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n552), .B2(new_n664), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1956), .ZN(new_n722));
  INV_X1    g297(.A(G1966), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G21), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G168), .B2(G16), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n722), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n704), .A2(G27), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G164), .B2(new_n704), .ZN(new_n729));
  INV_X1    g304(.A(G2078), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n664), .A2(G4), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n591), .B2(new_n664), .ZN(new_n733));
  INV_X1    g308(.A(G1348), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n727), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G29), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n475), .A2(G139), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n739), .B(new_n740), .C1(new_n463), .C2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(G29), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G2072), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(G2072), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n664), .A2(G19), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n540), .B2(new_n664), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n747), .A2(new_n748), .B1(G1341), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n704), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n704), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT29), .Z(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  INV_X1    g330(.A(new_n748), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(new_n745), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n751), .B(new_n757), .C1(G1341), .C2(new_n750), .ZN(new_n758));
  INV_X1    g333(.A(new_n754), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n759), .A2(G2090), .B1(G2067), .B2(new_n713), .ZN(new_n760));
  INV_X1    g335(.A(G28), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n761), .B2(KEYINPUT30), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(KEYINPUT30), .B2(new_n761), .ZN(new_n763));
  OR2_X1    g338(.A1(G29), .A2(G32), .ZN(new_n764));
  AOI22_X1  g339(.A1(G129), .A2(new_n473), .B1(new_n475), .B2(G141), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT26), .Z(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n764), .B1(new_n769), .B2(new_n704), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT27), .B(G1996), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n763), .B1(new_n704), .B2(new_n608), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G1966), .B2(new_n725), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT31), .B(G11), .ZN(new_n774));
  OR2_X1    g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n775), .A2(new_n704), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G160), .B2(new_n704), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2084), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n770), .B2(new_n771), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n760), .A2(new_n773), .A3(new_n774), .A4(new_n780), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n717), .A2(new_n736), .A3(new_n758), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n703), .A2(new_n714), .A3(new_n782), .ZN(G150));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n784));
  NAND2_X1  g359(.A1(G150), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n703), .A2(KEYINPUT93), .A3(new_n714), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(G311));
  NAND2_X1  g362(.A1(new_n508), .A2(G55), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT95), .B(G93), .ZN(new_n790));
  OAI221_X1 g365(.A(new_n788), .B1(new_n529), .B2(new_n789), .C1(new_n515), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G860), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT37), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n591), .A2(G559), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT39), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n540), .B(new_n791), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n795), .B(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n793), .B1(new_n799), .B2(G860), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT96), .ZN(G145));
  XOR2_X1   g376(.A(KEYINPUT99), .B(G37), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n473), .A2(G130), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n475), .A2(G142), .ZN(new_n804));
  NOR2_X1   g379(.A1(G106), .A2(G2105), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n803), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n689), .B(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT97), .ZN(new_n809));
  INV_X1    g384(.A(new_n599), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n744), .A2(new_n769), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n744), .A2(new_n769), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n711), .B(new_n495), .ZN(new_n814));
  OR3_X1    g389(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n812), .B2(new_n813), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT98), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n809), .B(new_n599), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n815), .A2(new_n816), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n817), .A2(KEYINPUT100), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n817), .A2(KEYINPUT100), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(new_n811), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(G160), .B(new_n608), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G162), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n823), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n811), .A2(new_n817), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n823), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n802), .B(new_n830), .C1(new_n832), .C2(new_n829), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT101), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g410(.A1(new_n670), .A2(new_n671), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G303), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n836), .A2(G303), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n677), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n839), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(new_n837), .A3(G305), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G290), .ZN(new_n844));
  INV_X1    g419(.A(G290), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n840), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT42), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n847), .A2(KEYINPUT103), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n848), .B1(new_n847), .B2(KEYINPUT103), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n591), .A2(new_n552), .ZN(new_n852));
  NAND2_X1  g427(.A1(G299), .A2(new_n582), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT41), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n856), .A3(new_n853), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT102), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n859));
  INV_X1    g434(.A(new_n854), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n859), .B1(new_n860), .B2(new_n856), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n594), .B(new_n796), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n854), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n851), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n868), .A2(new_n850), .A3(new_n849), .ZN(new_n869));
  OAI21_X1  g444(.A(G868), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n791), .A2(new_n583), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(G295));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n871), .ZN(G331));
  XNOR2_X1  g448(.A(new_n796), .B(G286), .ZN(new_n874));
  AND2_X1   g449(.A1(G301), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(G301), .A2(new_n874), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n860), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G301), .B(new_n874), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n862), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  INV_X1    g455(.A(new_n846), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n845), .B1(new_n840), .B2(new_n842), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n844), .A2(new_n846), .A3(KEYINPUT104), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n881), .A2(new_n882), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n886), .B(new_n877), .C1(new_n862), .C2(new_n878), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n877), .A2(KEYINPUT105), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n878), .A2(new_n892), .A3(new_n860), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n878), .B1(new_n857), .B2(new_n855), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n884), .B(new_n883), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n802), .A4(new_n887), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n890), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n889), .A2(new_n897), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n896), .A2(KEYINPUT43), .A3(new_n802), .A4(new_n887), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  MUX2_X1   g477(.A(new_n899), .B(new_n902), .S(KEYINPUT44), .Z(G397));
  AOI21_X1  g478(.A(G1384), .B1(new_n489), .B2(new_n494), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(KEYINPUT45), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n466), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n907), .B(G40), .C1(G2105), .C2(new_n461), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  INV_X1    g485(.A(G1986), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n845), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n910), .ZN(new_n913));
  NAND2_X1  g488(.A1(G290), .A2(G1986), .ZN(new_n914));
  MUX2_X1   g489(.A(new_n910), .B(new_n913), .S(new_n914), .Z(new_n915));
  XNOR2_X1  g490(.A(new_n769), .B(G1996), .ZN(new_n916));
  INV_X1    g491(.A(G2067), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n710), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n689), .B(new_n691), .Z(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n909), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n924));
  OAI21_X1  g499(.A(G1976), .B1(new_n670), .B2(new_n671), .ZN(new_n925));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n488), .A2(new_n487), .ZN(new_n927));
  INV_X1    g502(.A(new_n482), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n460), .B2(G126), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n929), .B2(new_n463), .ZN(new_n930));
  INV_X1    g505(.A(G138), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(KEYINPUT68), .B2(KEYINPUT4), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n460), .A2(new_n486), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(G2105), .B1(new_n933), .B2(new_n490), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n926), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT107), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n495), .A2(new_n937), .A3(new_n926), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n908), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G8), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(KEYINPUT109), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  INV_X1    g517(.A(new_n908), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n937), .B1(new_n495), .B2(new_n926), .ZN(new_n944));
  AOI211_X1 g519(.A(KEYINPUT107), .B(G1384), .C1(new_n489), .C2(new_n494), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n942), .B1(new_n946), .B2(G8), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n925), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT52), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT109), .B1(new_n939), .B2(new_n940), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n942), .A3(G8), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n953));
  INV_X1    g528(.A(G1976), .ZN(new_n954));
  NAND2_X1  g529(.A1(G288), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n952), .A2(new_n953), .A3(new_n955), .A4(new_n925), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n924), .B1(new_n949), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n924), .ZN(new_n958));
  XNOR2_X1  g533(.A(G305), .B(G1981), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT49), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n960), .A2(new_n952), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n908), .B1(new_n904), .B2(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n906), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(G1971), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n944), .B2(new_n945), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n935), .A2(KEYINPUT50), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(new_n943), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(G2090), .ZN(new_n971));
  OAI21_X1  g546(.A(G8), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(G303), .A2(G8), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT55), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT108), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n962), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n936), .A2(KEYINPUT50), .A3(new_n938), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n904), .A2(new_n967), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n943), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT112), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n980), .A2(new_n984), .A3(new_n943), .A4(new_n981), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(new_n755), .A3(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n965), .A2(G1971), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n940), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n974), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n979), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(G2090), .B1(new_n982), .B2(KEYINPUT112), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n966), .B1(new_n991), .B2(new_n985), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT113), .B(new_n974), .C1(new_n992), .C2(new_n940), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n978), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n936), .A2(new_n996), .A3(new_n938), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n963), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n723), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT114), .ZN(new_n1000));
  INV_X1    g575(.A(G2084), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n968), .A2(new_n1001), .A3(new_n969), .A4(new_n943), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(new_n1003), .A3(new_n723), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(G8), .A3(G286), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1000), .A2(new_n1002), .A3(G168), .A4(new_n1004), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT121), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(G8), .A3(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1014), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1009), .A2(G8), .A3(new_n1012), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1008), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT62), .ZN(new_n1020));
  AOI21_X1  g595(.A(G301), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT62), .B1(new_n1008), .B2(new_n1018), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT124), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n965), .B2(new_n730), .ZN(new_n1024));
  INV_X1    g599(.A(G1961), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(new_n970), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n730), .A2(KEYINPUT53), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n998), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT124), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(KEYINPUT62), .C1(new_n1008), .C2(new_n1018), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1021), .A2(new_n1023), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT57), .B1(new_n548), .B2(KEYINPUT117), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n552), .B(new_n1032), .Z(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT56), .B(G2072), .ZN(new_n1034));
  INV_X1    g609(.A(G1956), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n965), .A2(new_n1034), .B1(new_n982), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n970), .A2(new_n734), .B1(new_n917), .B2(new_n939), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n591), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT61), .B1(new_n1037), .B2(KEYINPUT119), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n964), .A2(G1996), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT58), .B(G1341), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n939), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n540), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1046));
  XNOR2_X1  g621(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT61), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1033), .A2(new_n1048), .A3(new_n1049), .A4(new_n1036), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1038), .A2(new_n1051), .A3(new_n591), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1041), .A2(new_n1047), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1039), .A2(new_n591), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1038), .A2(new_n582), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI221_X1 g631(.A(new_n1040), .B1(new_n1033), .B2(new_n1036), .C1(new_n1053), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1019), .ZN(new_n1058));
  XOR2_X1   g633(.A(G301), .B(KEYINPUT54), .Z(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1028), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n935), .A2(new_n996), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT122), .B1(new_n462), .B2(new_n466), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(G40), .C1(KEYINPUT122), .C2(new_n462), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(KEYINPUT123), .ZN(new_n1065));
  OR4_X1    g640(.A1(new_n1062), .A2(new_n1065), .A3(new_n905), .A4(new_n1027), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1059), .A2(new_n1026), .A3(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1057), .A2(new_n1058), .A3(new_n1061), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n995), .B1(new_n1031), .B2(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1005), .A2(G8), .A3(G168), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n962), .A2(new_n977), .A3(new_n994), .A4(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT115), .B(KEYINPUT63), .Z(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT116), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n972), .A2(new_n974), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n978), .A2(KEYINPUT63), .A3(new_n1070), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1071), .A2(new_n1077), .A3(new_n1072), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n962), .A2(new_n976), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n961), .A2(G1976), .A3(G288), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G305), .A2(G1981), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n952), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1079), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n923), .B1(new_n1069), .B2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT126), .B(KEYINPUT46), .ZN(new_n1089));
  INV_X1    g664(.A(new_n909), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(G1996), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n909), .B1(new_n769), .B2(new_n919), .ZN(new_n1092));
  INV_X1    g667(.A(G1996), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n909), .B(new_n1093), .C1(KEYINPUT126), .C2(KEYINPUT46), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n1095), .B(KEYINPUT47), .Z(new_n1096));
  NOR2_X1   g671(.A1(new_n689), .A2(new_n691), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n920), .B2(new_n1090), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(G2067), .B2(new_n710), .ZN(new_n1099));
  XOR2_X1   g674(.A(new_n1099), .B(KEYINPUT125), .Z(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n1090), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n912), .A2(new_n1090), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT127), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT48), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n922), .A2(new_n909), .ZN(new_n1105));
  AOI211_X1 g680(.A(new_n1096), .B(new_n1101), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1088), .A2(new_n1106), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g682(.A(G229), .ZN(new_n1109));
  NAND2_X1  g683(.A1(new_n1109), .A2(G319), .ZN(new_n1110));
  NOR2_X1   g684(.A1(G227), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g685(.A1(new_n899), .A2(new_n834), .A3(new_n628), .A4(new_n1111), .ZN(G225));
  INV_X1    g686(.A(G225), .ZN(G308));
endmodule


