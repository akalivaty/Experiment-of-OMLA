//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NAND2_X1  g002(.A1(G234), .A2(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AND3_X1   g004(.A1(new_n189), .A2(G952), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT67), .B(G953), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n194), .A2(G902), .A3(new_n189), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT21), .B(G898), .Z(new_n197));
  OAI21_X1  g011(.A(new_n192), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT79), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT77), .A2(G104), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT77), .A2(G104), .ZN(new_n202));
  OAI21_X1  g016(.A(G107), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n201), .A2(new_n202), .A3(G107), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT78), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR4_X1   g025(.A1(new_n208), .A2(KEYINPUT78), .A3(KEYINPUT3), .A4(G107), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n200), .B1(new_n206), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n207), .A3(new_n210), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n205), .A2(new_n210), .A3(G104), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT78), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OR2_X1    g032(.A1(KEYINPUT77), .A2(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT77), .A2(G104), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n210), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n218), .A2(new_n222), .A3(KEYINPUT79), .A4(new_n203), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n214), .A2(G101), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G101), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n218), .A2(new_n222), .A3(new_n225), .A4(new_n203), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n226), .A2(KEYINPUT4), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n214), .A2(new_n229), .A3(G101), .A4(new_n223), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G119), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G116), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT66), .B(G119), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n232), .B(new_n235), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n233), .A2(KEYINPUT66), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n236), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n231), .B1(new_n242), .B2(new_n234), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n228), .A2(new_n230), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n210), .A2(G104), .ZN(new_n246));
  OAI21_X1  g060(.A(G101), .B1(new_n204), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n226), .A2(KEYINPUT81), .A3(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n247), .A2(KEYINPUT81), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT5), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n240), .A2(G119), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n233), .A2(KEYINPUT66), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n251), .B(G116), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT84), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n242), .A2(KEYINPUT84), .A3(new_n251), .ZN(new_n257));
  OAI211_X1 g071(.A(KEYINPUT5), .B(new_n235), .C1(new_n237), .C2(new_n236), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n256), .A2(new_n257), .A3(G113), .A4(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n250), .A2(new_n238), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n245), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g075(.A(G110), .B(G122), .Z(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n262), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n245), .A2(new_n264), .A3(new_n260), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n263), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n245), .A2(new_n264), .A3(new_n260), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n245), .B2(new_n260), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n261), .A2(new_n269), .A3(new_n262), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT85), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n266), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G125), .ZN(new_n275));
  XNOR2_X1  g089(.A(G143), .B(G146), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT0), .ZN(new_n277));
  INV_X1    g091(.A(G128), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G146), .ZN(new_n281));
  INV_X1    g095(.A(G146), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(G143), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n277), .A2(new_n278), .ZN(new_n284));
  NOR2_X1   g098(.A1(KEYINPUT0), .A2(G128), .ZN(new_n285));
  OAI22_X1  g099(.A1(new_n281), .A2(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n275), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n276), .A2(new_n288), .A3(G128), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n280), .B(G146), .C1(new_n278), .C2(KEYINPUT1), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n278), .A2(new_n282), .A3(G143), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n290), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n289), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n287), .B1(new_n275), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n190), .A2(G224), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n274), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT88), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n302), .A2(KEYINPUT86), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n297), .B1(KEYINPUT86), .B2(new_n302), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n296), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT87), .ZN(new_n306));
  INV_X1    g120(.A(new_n297), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n295), .A2(new_n275), .ZN(new_n308));
  INV_X1    g122(.A(new_n287), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n306), .B1(new_n310), .B2(KEYINPUT7), .ZN(new_n311));
  NOR4_X1   g125(.A1(new_n296), .A2(KEYINPUT87), .A3(new_n302), .A4(new_n307), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n305), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n262), .B(KEYINPUT8), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n259), .A2(new_n238), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n248), .A3(new_n249), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n260), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n301), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n308), .A2(new_n309), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT7), .A3(new_n297), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT87), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n310), .A2(new_n306), .A3(KEYINPUT7), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n314), .ZN(new_n324));
  INV_X1    g138(.A(new_n316), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n315), .B1(new_n248), .B2(new_n249), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n323), .A2(new_n327), .A3(KEYINPUT88), .A4(new_n305), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n318), .A2(new_n265), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G902), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(G210), .B1(G237), .B2(G902), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT89), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n300), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n263), .A2(KEYINPUT6), .A3(new_n265), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT85), .B1(new_n268), .B2(new_n269), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n298), .B1(new_n339), .B2(new_n266), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n334), .B1(new_n340), .B2(new_n331), .ZN(new_n341));
  AOI211_X1 g155(.A(new_n188), .B(new_n199), .C1(new_n336), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G478), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(KEYINPUT15), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT9), .B(G234), .Z(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(G217), .A3(new_n190), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n236), .A2(G122), .ZN(new_n348));
  INV_X1    g162(.A(G122), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G116), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT14), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n236), .A2(KEYINPUT14), .A3(G122), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n352), .A2(G107), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n278), .A2(G143), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n280), .A2(G128), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n355), .B2(new_n356), .ZN(new_n359));
  OAI21_X1  g173(.A(G134), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n356), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT92), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n363));
  INV_X1    g177(.A(G134), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n354), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n348), .A2(new_n350), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT93), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n367), .A2(new_n368), .A3(new_n210), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n367), .B2(new_n210), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT94), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT94), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n366), .A2(new_n374), .A3(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n367), .B(new_n210), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT13), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n378), .B(G134), .C1(KEYINPUT13), .C2(new_n356), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n365), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n347), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n380), .ZN(new_n382));
  AOI211_X1 g196(.A(new_n382), .B(new_n346), .C1(new_n373), .C2(new_n375), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n330), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n344), .B1(new_n384), .B2(KEYINPUT95), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(KEYINPUT95), .ZN(new_n386));
  INV_X1    g200(.A(new_n375), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n374), .B1(new_n366), .B2(new_n371), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n380), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n346), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n376), .A2(new_n380), .A3(new_n347), .ZN(new_n391));
  AOI21_X1  g205(.A(G902), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT95), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n385), .B1(new_n395), .B2(new_n344), .ZN(new_n396));
  XNOR2_X1  g210(.A(G113), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n208), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n275), .A2(KEYINPUT16), .A3(G140), .ZN(new_n399));
  XNOR2_X1  g213(.A(G125), .B(G140), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n399), .B1(new_n400), .B2(KEYINPUT16), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n401), .A2(G146), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(G146), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT17), .ZN(new_n405));
  INV_X1    g219(.A(G131), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT64), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT64), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G131), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G237), .ZN(new_n411));
  AND2_X1   g225(.A1(KEYINPUT67), .A2(G953), .ZN(new_n412));
  NOR2_X1   g226(.A1(KEYINPUT67), .A2(G953), .ZN(new_n413));
  OAI211_X1 g227(.A(G214), .B(new_n411), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n280), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n193), .A2(G143), .A3(G214), .A4(new_n411), .ZN(new_n416));
  AOI211_X1 g230(.A(new_n405), .B(new_n410), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT90), .B1(new_n404), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n416), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n407), .A2(new_n409), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n415), .A2(new_n416), .A3(new_n410), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n405), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(KEYINPUT17), .A3(new_n420), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n402), .A4(new_n403), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n418), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(KEYINPUT18), .A2(G131), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n419), .B(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n400), .A2(new_n282), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT75), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n282), .B2(new_n400), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n398), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n427), .A2(new_n398), .A3(new_n433), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT91), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT91), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n427), .A2(new_n437), .A3(new_n398), .A4(new_n433), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n434), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G475), .B1(new_n439), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  INV_X1    g255(.A(new_n398), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n421), .A2(new_n422), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n400), .B(KEYINPUT19), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n282), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n403), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n433), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n436), .A2(new_n438), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(G475), .A2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n441), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n436), .A2(new_n438), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(new_n442), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT20), .A3(new_n449), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n396), .A2(new_n440), .A3(new_n451), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n364), .A2(G137), .ZN(new_n457));
  INV_X1    g271(.A(G137), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G134), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G131), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT11), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n364), .B2(G137), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n458), .A2(KEYINPUT11), .A3(G134), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n457), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n461), .B1(new_n465), .B2(new_n420), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n290), .A2(new_n292), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT65), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n466), .B1(new_n470), .B2(new_n289), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n465), .A2(G131), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n410), .A2(new_n457), .A3(new_n464), .A4(new_n463), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n472), .A2(new_n473), .B1(new_n279), .B2(new_n286), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n471), .A2(KEYINPUT30), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n463), .A2(new_n457), .A3(new_n464), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n477), .A2(new_n410), .B1(G131), .B2(new_n460), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n295), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n472), .A2(new_n473), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n279), .A2(new_n286), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n476), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n244), .B1(new_n475), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n193), .A2(G210), .A3(new_n411), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n485), .B(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT26), .B(G101), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n238), .A2(new_n243), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n479), .A2(new_n490), .A3(new_n482), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n484), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT31), .ZN(new_n493));
  INV_X1    g307(.A(new_n489), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n244), .B1(new_n471), .B2(new_n474), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(new_n491), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT28), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n494), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT31), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n484), .A2(new_n502), .A3(new_n489), .A4(new_n491), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n493), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(G472), .A2(G902), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT32), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT70), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n510), .A3(new_n505), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n508), .B1(new_n512), .B2(new_n507), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n494), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT72), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n491), .A2(new_n517), .A3(new_n498), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT71), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n496), .A2(new_n491), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n520), .B1(new_n521), .B2(KEYINPUT28), .ZN(new_n522));
  AOI211_X1 g336(.A(KEYINPUT71), .B(new_n498), .C1(new_n496), .C2(new_n491), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n515), .B(new_n519), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n330), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT73), .ZN(new_n526));
  OR3_X1    g340(.A1(new_n500), .A2(new_n497), .A3(new_n494), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n484), .A2(new_n491), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n494), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n514), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT73), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n531), .A3(new_n330), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G472), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n456), .B1(new_n513), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n345), .ZN(new_n536));
  OAI21_X1  g350(.A(G221), .B1(new_n536), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n228), .A2(new_n481), .A3(new_n230), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT80), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT80), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n228), .A2(new_n541), .A3(new_n481), .A4(new_n230), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n480), .ZN(new_n544));
  INV_X1    g358(.A(new_n467), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n289), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n250), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT82), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT10), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n248), .A2(new_n249), .B1(new_n289), .B2(new_n545), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT82), .B1(new_n551), .B2(KEYINPUT10), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n250), .A2(KEYINPUT10), .A3(new_n295), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n543), .A2(new_n544), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n193), .A2(G227), .ZN(new_n556));
  XNOR2_X1  g370(.A(G110), .B(G140), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n543), .A2(new_n553), .A3(new_n554), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n480), .ZN(new_n561));
  INV_X1    g375(.A(new_n295), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n248), .A2(new_n249), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n480), .B1(new_n563), .B2(new_n551), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT12), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(KEYINPUT12), .B(new_n480), .C1(new_n563), .C2(new_n551), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n555), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n558), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n559), .A2(new_n561), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G469), .B1(new_n571), .B2(G902), .ZN(new_n572));
  INV_X1    g386(.A(G469), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n558), .B1(new_n561), .B2(new_n555), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT83), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n248), .A2(new_n249), .A3(new_n562), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n547), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT12), .B1(new_n577), .B2(new_n480), .ZN(new_n578));
  INV_X1    g392(.A(new_n567), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n566), .A2(KEYINPUT83), .A3(new_n567), .ZN(new_n581));
  AND4_X1   g395(.A1(new_n555), .A2(new_n580), .A3(new_n558), .A4(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n573), .B(new_n330), .C1(new_n574), .C2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n538), .B1(new_n572), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT23), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n237), .A2(new_n585), .A3(new_n278), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n233), .A2(G128), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n237), .B2(new_n278), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n586), .B1(new_n589), .B2(new_n585), .ZN(new_n590));
  INV_X1    g404(.A(G110), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n589), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT24), .B(G110), .Z(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n403), .B(new_n431), .C1(new_n592), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n594), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n404), .B(new_n597), .C1(new_n591), .C2(new_n590), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(KEYINPUT22), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G137), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n601), .B(new_n458), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n596), .A3(new_n598), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n605), .A3(new_n330), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n607));
  INV_X1    g421(.A(G217), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(G234), .B2(new_n330), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT74), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n609), .A2(KEYINPUT74), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT76), .B(KEYINPUT25), .Z(new_n612));
  NAND4_X1  g426(.A1(new_n603), .A2(new_n605), .A3(new_n330), .A4(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n607), .A2(new_n610), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n603), .A2(new_n605), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n609), .A2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n342), .A2(new_n535), .A3(new_n584), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G101), .ZN(G3));
  NAND2_X1  g435(.A1(G469), .A2(G902), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n561), .A2(new_n555), .A3(new_n558), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n569), .A2(new_n570), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(G469), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n583), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G472), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n504), .B2(new_n330), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n509), .B2(new_n511), .ZN(new_n629));
  AND4_X1   g443(.A1(new_n537), .A2(new_n626), .A3(new_n619), .A4(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n188), .B1(new_n336), .B2(new_n341), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n390), .A2(new_n391), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT33), .B1(new_n632), .B2(KEYINPUT96), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT96), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n634), .B(new_n635), .C1(new_n390), .C2(new_n391), .ZN(new_n636));
  OAI211_X1 g450(.A(G478), .B(new_n330), .C1(new_n633), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n384), .A2(new_n343), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n455), .A2(new_n451), .A3(new_n440), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n631), .A2(new_n198), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n630), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND2_X1  g461(.A1(new_n336), .A2(new_n341), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n640), .A2(new_n396), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n648), .A2(new_n187), .A3(new_n198), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n630), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  OR2_X1    g468(.A1(new_n599), .A2(KEYINPUT97), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n599), .A2(KEYINPUT97), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n602), .A2(KEYINPUT36), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n655), .A2(new_n658), .A3(new_n656), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n616), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n614), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n629), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n456), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n342), .A2(new_n584), .A3(new_n664), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT37), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n591), .ZN(G12));
  AND3_X1   g483(.A1(new_n504), .A2(new_n510), .A3(new_n505), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n510), .B1(new_n504), .B2(new_n505), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n507), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n508), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n534), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n674), .A2(new_n648), .A3(new_n187), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n192), .B1(new_n196), .B2(G900), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n640), .A2(new_n396), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n675), .A2(new_n584), .A3(new_n664), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT98), .B(G128), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G30));
  XOR2_X1   g495(.A(new_n648), .B(KEYINPUT99), .Z(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT38), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n648), .B(KEYINPUT99), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT38), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n528), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n494), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n330), .B1(new_n521), .B2(new_n489), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n513), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n392), .A2(new_n393), .ZN(new_n693));
  AOI211_X1 g507(.A(KEYINPUT95), .B(G902), .C1(new_n390), .C2(new_n391), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n344), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n385), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n640), .A2(new_n697), .A3(new_n187), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n687), .A2(new_n663), .A3(new_n692), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n676), .B(KEYINPUT39), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n584), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT40), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT100), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n280), .ZN(G45));
  NOR2_X1   g520(.A1(new_n641), .A2(new_n677), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n675), .A2(new_n584), .A3(new_n664), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  OAI21_X1  g523(.A(new_n330), .B1(new_n574), .B2(new_n582), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n537), .A3(new_n583), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n674), .A2(new_n619), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n644), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n651), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  AND3_X1   g533(.A1(new_n711), .A2(new_n537), .A3(new_n583), .ZN(new_n720));
  AOI211_X1 g534(.A(new_n188), .B(new_n663), .C1(new_n336), .C2(new_n341), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n342), .A3(new_n721), .A4(new_n535), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT101), .B(G119), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G21));
  NOR2_X1   g538(.A1(new_n522), .A2(new_n523), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n516), .B2(new_n518), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n493), .B(new_n503), .C1(new_n726), .C2(new_n489), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n628), .B1(new_n727), .B2(new_n505), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n619), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n199), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n698), .B1(new_n341), .B2(new_n336), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n720), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  INV_X1    g547(.A(new_n728), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n734), .A2(new_n641), .A3(new_n677), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n720), .A2(new_n721), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  NOR2_X1   g551(.A1(new_n648), .A2(new_n188), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n584), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n506), .B(KEYINPUT32), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n618), .B1(new_n740), .B2(new_n534), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n707), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n713), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n584), .A3(new_n707), .A4(new_n738), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  AND4_X1   g562(.A1(new_n584), .A2(new_n743), .A3(new_n738), .A4(new_n678), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n364), .ZN(G36));
  NAND2_X1  g564(.A1(new_n571), .A2(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n623), .A2(new_n624), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(new_n754), .A3(G469), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT46), .B1(new_n755), .B2(new_n622), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(KEYINPUT102), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(KEYINPUT102), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n622), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n583), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n538), .ZN(new_n762));
  INV_X1    g576(.A(new_n640), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n639), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT103), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT43), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n665), .A3(new_n664), .A4(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n762), .A2(new_n701), .A3(new_n772), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n738), .B(KEYINPUT104), .Z(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n770), .B2(new_n771), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  NAND2_X1  g592(.A1(new_n762), .A2(KEYINPUT47), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n761), .B2(new_n538), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n674), .A2(new_n619), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n707), .A3(new_n738), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  NAND3_X1  g599(.A1(new_n768), .A2(new_n191), .A3(new_n769), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n729), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(new_n774), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n711), .A2(new_n538), .A3(new_n583), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT115), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n791), .B1(new_n782), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n788), .A2(new_n789), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n720), .A2(new_n738), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT116), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n734), .A2(new_n663), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n729), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n187), .B1(new_n683), .B2(new_n686), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n795), .A2(new_n720), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n790), .A2(KEYINPUT50), .A3(new_n720), .A4(new_n801), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n692), .A2(new_n618), .A3(new_n192), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n797), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n639), .A2(new_n640), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n794), .A2(new_n806), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n810), .B(new_n799), .C1(new_n804), .C2(new_n805), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n779), .A2(new_n781), .A3(new_n792), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n813), .B1(new_n815), .B2(new_n791), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n812), .A2(new_n813), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n795), .A2(new_n741), .A3(new_n797), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT48), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n795), .A2(new_n631), .A3(new_n720), .A4(new_n800), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n797), .A2(new_n642), .A3(new_n807), .ZN(new_n821));
  AND4_X1   g635(.A1(G952), .A2(new_n820), .A3(new_n190), .A4(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n819), .A2(new_n822), .A3(KEYINPUT117), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT117), .B1(new_n819), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n676), .B(KEYINPUT111), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n614), .A2(new_n662), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT112), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n731), .A2(new_n584), .A3(new_n692), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n679), .A2(new_n708), .A3(new_n736), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT113), .ZN(new_n831));
  INV_X1    g645(.A(new_n555), .ZN(new_n832));
  INV_X1    g646(.A(new_n554), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n540), .B2(new_n542), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n544), .B1(new_n834), .B2(new_n553), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n570), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n555), .A2(new_n580), .A3(new_n558), .A4(new_n581), .ZN(new_n837));
  AOI211_X1 g651(.A(G469), .B(G902), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n625), .A2(new_n622), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n537), .B(new_n664), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n674), .A2(new_n648), .A3(new_n187), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n335), .B1(new_n300), .B2(new_n332), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n340), .A2(new_n334), .A3(new_n331), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n187), .B(new_n664), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n712), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n842), .A2(new_n678), .B1(new_n846), .B2(new_n735), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n708), .A4(new_n829), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n831), .A2(new_n849), .A3(KEYINPUT52), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(new_n831), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT106), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT106), .B1(new_n639), .B2(new_n640), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n648), .A2(new_n187), .A3(new_n198), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT107), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT106), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n641), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT106), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT107), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n342), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n857), .A2(new_n863), .A3(new_n630), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n620), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT108), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(KEYINPUT108), .A3(new_n620), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n535), .A2(new_n676), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n870), .A2(new_n735), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n584), .A3(new_n664), .A4(new_n738), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n749), .B1(new_n742), .B2(new_n746), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n722), .A2(new_n667), .A3(new_n732), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n713), .B(new_n712), .C1(new_n643), .C2(new_n650), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n649), .A2(KEYINPUT109), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n649), .A2(KEYINPUT109), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n342), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n584), .A2(new_n619), .A3(new_n629), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n874), .A2(new_n875), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n869), .A2(new_n872), .A3(new_n873), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n852), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n679), .A2(new_n736), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(KEYINPUT110), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(KEYINPUT110), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n829), .A2(KEYINPUT52), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n886), .A2(new_n708), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n831), .A2(new_n849), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(KEYINPUT52), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n864), .A2(KEYINPUT108), .A3(new_n620), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT108), .B1(new_n864), .B2(new_n620), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n881), .B(new_n873), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n872), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT53), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT54), .B1(new_n884), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n883), .B1(new_n852), .B2(new_n882), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n891), .A2(new_n896), .A3(KEYINPUT53), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n817), .A2(new_n825), .A3(new_n898), .A4(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(G952), .A2(G953), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT118), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n711), .A2(new_n583), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n618), .B1(new_n907), .B2(KEYINPUT49), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n764), .A2(new_n188), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n537), .A3(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT105), .Z(new_n911));
  NOR2_X1   g725(.A1(new_n907), .A2(KEYINPUT49), .ZN(new_n912));
  OR4_X1    g726(.A1(new_n692), .A2(new_n911), .A3(new_n687), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n906), .A2(new_n913), .ZN(G75));
  NAND2_X1  g728(.A1(new_n899), .A2(new_n900), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(G902), .A3(new_n334), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n274), .B(KEYINPUT119), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n298), .B(KEYINPUT55), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n920), .B1(new_n916), .B2(new_n917), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n193), .A2(G952), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G51));
  XOR2_X1   g738(.A(new_n622), .B(KEYINPUT57), .Z(new_n925));
  AND3_X1   g739(.A1(new_n899), .A2(new_n901), .A3(new_n900), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n901), .B1(new_n899), .B2(new_n900), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n574), .A2(new_n582), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n330), .B1(new_n899), .B2(new_n900), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n755), .B(KEYINPUT120), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n923), .B1(new_n931), .B2(new_n934), .ZN(G54));
  NAND3_X1  g749(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n448), .ZN(new_n937));
  INV_X1    g751(.A(new_n923), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .A4(new_n454), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(G60));
  OR2_X1    g754(.A1(new_n633), .A2(new_n636), .ZN(new_n941));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT59), .Z(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n941), .B(new_n944), .C1(new_n926), .C2(new_n927), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n898), .B2(new_n902), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n945), .B(new_n938), .C1(new_n946), .C2(new_n941), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(G63));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  XNOR2_X1  g763(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT122), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n608), .A2(new_n330), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n915), .A2(new_n661), .A3(new_n660), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n938), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n615), .B1(new_n915), .B2(new_n953), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n956), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n958), .A2(KEYINPUT61), .A3(new_n938), .A4(new_n954), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(G66));
  AOI21_X1  g774(.A(new_n190), .B1(new_n197), .B2(G224), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n869), .A2(new_n881), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n962), .B2(new_n193), .ZN(new_n963));
  INV_X1    g777(.A(G898), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n918), .B1(new_n964), .B2(new_n194), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n963), .B(new_n965), .ZN(G69));
  NAND3_X1  g780(.A1(new_n886), .A2(new_n708), .A3(new_n887), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n762), .A2(new_n701), .A3(new_n731), .A4(new_n741), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n969), .A2(new_n873), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n784), .A2(new_n777), .A3(new_n968), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n193), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n475), .A2(new_n483), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT123), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(new_n444), .Z(new_n975));
  NAND2_X1  g789(.A1(new_n194), .A2(G900), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n972), .B(new_n975), .C1(G227), .C2(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n704), .B2(new_n967), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n876), .A2(new_n877), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n855), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n701), .A2(new_n981), .A3(new_n743), .A4(new_n739), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n773), .B2(new_n776), .ZN(new_n983));
  NAND2_X1  g797(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n968), .B(new_n984), .C1(new_n700), .C2(new_n703), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n784), .A2(new_n979), .A3(new_n983), .A4(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(G227), .ZN(new_n987));
  OAI22_X1  g801(.A1(new_n986), .A2(new_n194), .B1(new_n987), .B2(new_n976), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n977), .B1(new_n975), .B2(new_n988), .ZN(G72));
  XNOR2_X1  g803(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n971), .B2(new_n962), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n494), .A3(new_n688), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n993), .B1(new_n986), .B2(new_n962), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n689), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n529), .A2(new_n492), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n993), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT127), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n884), .B2(new_n897), .ZN(new_n1001));
  AND4_X1   g815(.A1(new_n938), .A2(new_n995), .A3(new_n997), .A4(new_n1001), .ZN(G57));
endmodule


