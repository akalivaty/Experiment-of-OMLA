//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G211gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G231gat), .A2(G233gat), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT16), .ZN(new_n206));
  INV_X1    g005(.A(G15gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G15gat), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(G1gat), .B1(new_n208), .B2(new_n210), .ZN(new_n212));
  OAI21_X1  g011(.A(G8gat), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n210), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(new_n205), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n216));
  INV_X1    g015(.A(G8gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G64gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT86), .B1(new_n220), .B2(G57gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT86), .ZN(new_n222));
  INV_X1    g021(.A(G57gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(G64gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n221), .B(new_n224), .C1(new_n223), .C2(G64gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(G71gat), .B(G78gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227));
  INV_X1    g026(.A(G71gat), .ZN(new_n228));
  INV_X1    g027(.A(G78gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n225), .A2(new_n226), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n226), .ZN(new_n232));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n219), .B1(new_n236), .B2(KEYINPUT21), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(G183gat), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n236), .A2(KEYINPUT21), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(new_n239), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n204), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n240), .A2(new_n241), .A3(new_n204), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n203), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n244), .ZN(new_n246));
  INV_X1    g045(.A(new_n203), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n242), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n245), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n245), .B2(new_n248), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(KEYINPUT90), .A2(G99gat), .A3(G106gat), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT90), .B1(G99gat), .B2(G106gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G85gat), .ZN(new_n257));
  INV_X1    g056(.A(G92gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n256), .A2(KEYINPUT8), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G99gat), .B(G106gat), .Z(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G85gat), .A2(G92gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT89), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT7), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n263), .ZN(new_n266));
  NAND3_X1  g065(.A1(KEYINPUT89), .A2(G85gat), .A3(G92gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n259), .A2(new_n261), .A3(new_n265), .A4(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n255), .ZN(new_n270));
  NAND3_X1  g069(.A1(KEYINPUT90), .A2(G99gat), .A3(G106gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(KEYINPUT8), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n258), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n265), .A4(new_n268), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n260), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G29gat), .A2(G36gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT14), .ZN(new_n278));
  INV_X1    g077(.A(G29gat), .ZN(new_n279));
  INV_X1    g078(.A(G36gat), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .A4(KEYINPUT80), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(G29gat), .A2(G36gat), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT80), .B1(new_n284), .B2(new_n278), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n277), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G43gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G50gat), .ZN(new_n288));
  INV_X1    g087(.A(G50gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G43gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n290), .A3(KEYINPUT15), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n289), .B2(G43gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n287), .A2(KEYINPUT82), .A3(G50gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT15), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n278), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n300), .A2(new_n282), .B1(G29gat), .B2(G36gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT81), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n288), .A2(new_n290), .A3(KEYINPUT81), .A4(KEYINPUT15), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n299), .A2(new_n301), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT17), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n293), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n306), .B1(new_n293), .B2(new_n305), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n276), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT91), .ZN(new_n310));
  INV_X1    g109(.A(new_n276), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n305), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT91), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n314), .B(new_n276), .C1(new_n307), .C2(new_n308), .ZN(new_n315));
  AND2_X1   g114(.A1(G232gat), .A2(G233gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT41), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n310), .A2(new_n313), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT92), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n309), .A2(KEYINPUT91), .B1(KEYINPUT41), .B2(new_n316), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n321), .A2(KEYINPUT92), .A3(new_n313), .A4(new_n315), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G190gat), .B(G218gat), .Z(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n320), .A2(new_n324), .A3(new_n322), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(KEYINPUT88), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n316), .A2(KEYINPUT41), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT87), .ZN(new_n330));
  XNOR2_X1  g129(.A(G134gat), .B(G162gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n326), .A2(KEYINPUT88), .A3(new_n327), .A4(new_n332), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n253), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT93), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n235), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n231), .A2(KEYINPUT93), .A3(new_n234), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n276), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n269), .A2(new_n275), .A3(new_n235), .A4(new_n339), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT10), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT94), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n276), .A2(new_n345), .A3(new_n235), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G230gat), .A2(G233gat), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT10), .B1(new_n342), .B2(new_n343), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT94), .B1(new_n352), .B2(new_n348), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n351), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n342), .A2(new_n355), .A3(new_n343), .ZN(new_n356));
  XNOR2_X1  g155(.A(G120gat), .B(G148gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(G176gat), .B(G204gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT95), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT95), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n354), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n352), .A2(new_n348), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n356), .B1(new_n366), .B2(new_n355), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n363), .A2(new_n365), .B1(new_n359), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n338), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n213), .A2(new_n218), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n307), .B2(new_n308), .ZN(new_n371));
  NAND2_X1  g170(.A1(G229gat), .A2(G233gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n312), .A2(new_n219), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n371), .A2(KEYINPUT18), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n312), .B2(new_n219), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n370), .A2(KEYINPUT83), .A3(new_n293), .A4(new_n305), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n372), .B(KEYINPUT13), .Z(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT84), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n382), .A3(new_n379), .ZN(new_n383));
  XNOR2_X1  g182(.A(G113gat), .B(G141gat), .ZN(new_n384));
  INV_X1    g183(.A(G197gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT11), .B(G169gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(KEYINPUT12), .ZN(new_n389));
  AND4_X1   g188(.A1(new_n374), .A2(new_n381), .A3(new_n383), .A4(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT18), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT85), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n395), .A3(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n381), .A2(new_n393), .A3(new_n374), .A4(new_n383), .ZN(new_n399));
  INV_X1    g198(.A(new_n389), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT27), .B(G183gat), .ZN(new_n404));
  INV_X1    g203(.A(G190gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409));
  INV_X1    g208(.A(G169gat), .ZN(new_n410));
  INV_X1    g209(.A(G176gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT26), .ZN(new_n413));
  NOR2_X1   g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n413), .B2(new_n414), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n408), .A2(new_n409), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n412), .B1(KEYINPUT23), .B2(new_n414), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT24), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n409), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n420), .B(new_n421), .C1(G183gat), .C2(G190gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT25), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n414), .A2(KEYINPUT23), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n418), .A2(new_n422), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT64), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n418), .B(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n409), .A2(KEYINPUT65), .A3(new_n419), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(G183gat), .B2(G190gat), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n409), .B1(KEYINPUT65), .B2(new_n419), .ZN(new_n430));
  OR2_X1    g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n427), .A2(new_n424), .A3(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n417), .B(new_n425), .C1(new_n432), .C2(new_n423), .ZN(new_n433));
  INV_X1    g232(.A(G120gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(G113gat), .ZN(new_n435));
  INV_X1    g234(.A(G113gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G120gat), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT1), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT67), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G127gat), .B(G134gat), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n438), .A2(new_n439), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n433), .B(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G15gat), .B(G43gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT34), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n448), .B2(KEYINPUT32), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n448), .A2(KEYINPUT32), .A3(new_n455), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n446), .A2(new_n447), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n457), .B2(new_n458), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n454), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n463), .ZN(new_n465));
  INV_X1    g264(.A(new_n454), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n461), .ZN(new_n467));
  XNOR2_X1  g266(.A(G197gat), .B(G204gat), .ZN(new_n468));
  AND2_X1   g267(.A1(G211gat), .A2(G218gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(KEYINPUT22), .B2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(G211gat), .B(G218gat), .Z(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT29), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT3), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G141gat), .B(G148gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(G155gat), .B(G162gat), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT72), .B(G155gat), .Z(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT73), .B(G162gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI211_X1 g279(.A(new_n475), .B(new_n477), .C1(new_n480), .C2(KEYINPUT2), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n475), .A2(KEYINPUT2), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n476), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT3), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n473), .ZN(new_n488));
  INV_X1    g287(.A(new_n472), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G228gat), .A2(G233gat), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n490), .B(new_n491), .Z(new_n492));
  XNOR2_X1  g291(.A(G78gat), .B(G106gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT31), .B(G50gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT76), .A3(G22gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(G22gat), .B2(new_n495), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n492), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n464), .A2(new_n467), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G1gat), .B(G29gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(G85gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT0), .B(G57gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n502), .B(new_n503), .Z(new_n504));
  INV_X1    g303(.A(new_n484), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT3), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(new_n445), .A3(new_n487), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n484), .A2(new_n444), .A3(new_n442), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT4), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n509), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G225gat), .A2(G233gat), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT74), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n505), .A2(new_n445), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n508), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(new_n518), .B2(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n515), .A2(new_n519), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n504), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n515), .A2(new_n519), .ZN(new_n524));
  INV_X1    g323(.A(new_n504), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n526), .A2(new_n527), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n523), .A2(new_n526), .A3(KEYINPUT75), .A4(new_n527), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT71), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n433), .A2(G226gat), .A3(G233gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n433), .A2(new_n473), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT69), .ZN(new_n537));
  NAND2_X1  g336(.A1(G226gat), .A2(G233gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n489), .B(new_n535), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(new_n538), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n535), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n472), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G8gat), .B(G36gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(new_n258), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT70), .B(G64gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n548), .B(new_n549), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT30), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n534), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n546), .A2(KEYINPUT71), .A3(KEYINPUT30), .A4(new_n550), .ZN(new_n555));
  INV_X1    g354(.A(new_n550), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n542), .A2(new_n545), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n500), .A2(new_n533), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n464), .A2(new_n467), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(new_n558), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT35), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT77), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n528), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n523), .A2(new_n526), .A3(KEYINPUT77), .A4(new_n527), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n531), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n563), .A2(new_n564), .A3(new_n499), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT39), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n571), .B(new_n514), .C1(new_n517), .C2(new_n508), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n512), .B(new_n571), .ZN(new_n573));
  AOI211_X1 g372(.A(new_n525), .B(new_n572), .C1(new_n573), .C2(new_n514), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT40), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n576), .A3(new_n526), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT37), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n546), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n542), .A2(KEYINPUT37), .A3(new_n545), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n556), .A3(new_n580), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n581), .A2(KEYINPUT38), .B1(new_n546), .B2(new_n550), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n582), .A2(new_n566), .A3(new_n531), .A4(new_n567), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT38), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n544), .A2(new_n489), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n585), .A2(KEYINPUT79), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n472), .B(new_n535), .C1(new_n540), .C2(new_n541), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT78), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n541), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(new_n539), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n591), .A2(KEYINPUT78), .A3(new_n472), .A4(new_n535), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n585), .A2(KEYINPUT79), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n586), .A2(new_n589), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT37), .ZN(new_n595));
  AND4_X1   g394(.A1(new_n584), .A2(new_n595), .A3(new_n556), .A4(new_n579), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n577), .B(new_n499), .C1(new_n583), .C2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n533), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n498), .B1(new_n598), .B2(new_n558), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n562), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n464), .A2(new_n467), .A3(KEYINPUT36), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n369), .B(new_n403), .C1(new_n570), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n598), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n558), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT96), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n610), .A3(new_n558), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(G8gat), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n611), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT16), .B(G8gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT97), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT42), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n605), .A2(KEYINPUT42), .A3(new_n558), .A4(new_n617), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n614), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n614), .A2(new_n620), .A3(KEYINPUT99), .A4(new_n621), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(G1325gat));
  INV_X1    g425(.A(new_n605), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n207), .B1(new_n627), .B2(new_n562), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT100), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n627), .A2(new_n207), .A3(new_n603), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(G1326gat));
  NAND2_X1  g430(.A1(new_n605), .A2(new_n498), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G22gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(G1327gat));
  AOI21_X1  g434(.A(new_n336), .B1(new_n570), .B2(new_n604), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n367), .A2(new_n359), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n354), .A2(new_n364), .A3(new_n361), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n364), .B1(new_n354), .B2(new_n361), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n252), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n636), .A2(new_n402), .A3(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n642), .A2(G29gat), .A3(new_n533), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT45), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n604), .A2(KEYINPUT103), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n597), .A2(new_n599), .A3(new_n646), .A4(new_n603), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n570), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n337), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI211_X1 g450(.A(new_n650), .B(new_n336), .C1(new_n570), .C2(new_n604), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654));
  AOI221_X4 g453(.A(new_n654), .B1(new_n399), .B2(new_n400), .C1(new_n390), .C2(new_n397), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT102), .B1(new_n398), .B2(new_n401), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n651), .A2(new_n653), .A3(new_n658), .A4(new_n641), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT104), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT44), .B1(new_n648), .B2(new_n337), .ZN(new_n661));
  INV_X1    g460(.A(new_n641), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n661), .A2(new_n662), .A3(new_n652), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n658), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n533), .B1(new_n660), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n644), .B1(new_n666), .B2(new_n279), .ZN(G1328gat));
  INV_X1    g466(.A(new_n642), .ZN(new_n668));
  NAND2_X1  g467(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n668), .A2(new_n280), .A3(new_n558), .A4(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n559), .B1(new_n660), .B2(new_n665), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n672), .B1(new_n673), .B2(new_n280), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n672), .B(KEYINPUT106), .C1(new_n673), .C2(new_n280), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(G1329gat));
  OAI21_X1  g477(.A(G43gat), .B1(new_n659), .B2(new_n603), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n642), .A2(G43gat), .A3(new_n562), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(KEYINPUT47), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n603), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n659), .A2(KEYINPUT104), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n664), .B1(new_n663), .B2(new_n658), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n680), .B1(new_n686), .B2(G43gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n687), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g487(.A(G50gat), .B1(new_n659), .B2(new_n499), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n642), .A2(G50gat), .A3(new_n499), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(KEYINPUT48), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n498), .B1(new_n684), .B2(new_n685), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n690), .B1(new_n693), .B2(G50gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n694), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g494(.A1(new_n658), .A2(new_n368), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n648), .A2(new_n338), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n533), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(new_n223), .ZN(G1332gat));
  INV_X1    g498(.A(KEYINPUT49), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n697), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n558), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT108), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n702), .A2(new_n706), .A3(new_n558), .A4(new_n703), .ZN(new_n707));
  AND4_X1   g506(.A1(new_n700), .A2(new_n705), .A3(new_n220), .A4(new_n707), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n705), .A2(new_n707), .B1(new_n700), .B2(new_n220), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(G1333gat));
  OR3_X1    g509(.A1(new_n697), .A2(G71gat), .A3(new_n562), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n702), .A2(new_n683), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(new_n228), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT50), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1334gat));
  NAND2_X1  g514(.A1(new_n702), .A2(new_n498), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT109), .B(G78gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1335gat));
  NOR3_X1   g517(.A1(new_n661), .A2(new_n252), .A3(new_n652), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n696), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(new_n257), .A3(new_n533), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n252), .A2(new_n658), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n648), .A2(new_n337), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(new_n640), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n598), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n721), .B1(new_n727), .B2(new_n257), .ZN(G1336gat));
  AND4_X1   g527(.A1(new_n258), .A2(new_n725), .A3(new_n640), .A4(new_n558), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT52), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n720), .A2(new_n559), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n730), .B(new_n731), .C1(new_n258), .C2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n258), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT52), .B1(new_n734), .B2(new_n729), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1337gat));
  NOR2_X1   g535(.A1(new_n661), .A2(new_n652), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n737), .A2(new_n253), .A3(new_n683), .A4(new_n696), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n719), .A2(KEYINPUT110), .A3(new_n683), .A4(new_n696), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(G99gat), .A3(new_n741), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n562), .A2(G99gat), .A3(new_n368), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT111), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n725), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n742), .A2(KEYINPUT112), .A3(new_n745), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1338gat));
  OAI211_X1 g549(.A(KEYINPUT53), .B(G106gat), .C1(new_n720), .C2(new_n499), .ZN(new_n751));
  INV_X1    g550(.A(G106gat), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n725), .A2(new_n752), .A3(new_n640), .A4(new_n498), .ZN(new_n753));
  OR2_X1    g552(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n751), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n753), .A2(KEYINPUT113), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT114), .B1(new_n720), .B2(new_n499), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n719), .A2(new_n758), .A3(new_n498), .A4(new_n696), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(G106gat), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n755), .B1(new_n761), .B2(new_n762), .ZN(G1339gat));
  NOR2_X1   g562(.A1(new_n378), .A2(new_n379), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n388), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT115), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n398), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n640), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n771), .B(new_n351), .C1(new_n352), .C2(new_n348), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n359), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(new_n366), .B2(new_n355), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n354), .B2(new_n774), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n363), .A2(new_n365), .B1(new_n775), .B2(KEYINPUT55), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n354), .A2(new_n774), .ZN(new_n777));
  INV_X1    g576(.A(new_n773), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT55), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n770), .B1(new_n657), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n336), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n638), .A2(new_n639), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785));
  AOI211_X1 g584(.A(new_n785), .B(new_n773), .C1(new_n354), .C2(new_n774), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n784), .A2(new_n786), .A3(new_n779), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n337), .A2(new_n787), .A3(new_n769), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n252), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n252), .A2(new_n336), .A3(new_n368), .A4(new_n657), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT116), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n334), .A2(new_n335), .A3(new_n780), .A4(new_n776), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n336), .A2(new_n782), .B1(new_n795), .B2(new_n769), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n793), .B(new_n790), .C1(new_n796), .C2(new_n252), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n798), .A2(new_n598), .A3(new_n499), .A4(new_n563), .ZN(new_n799));
  OAI21_X1  g598(.A(G113gat), .B1(new_n799), .B2(new_n403), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n658), .A2(new_n436), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(G1340gat));
  NOR2_X1   g601(.A1(new_n799), .A2(new_n368), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(new_n434), .ZN(G1341gat));
  NOR2_X1   g603(.A1(new_n799), .A2(new_n253), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g605(.A1(new_n799), .A2(new_n336), .ZN(new_n807));
  NOR2_X1   g606(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n808));
  AND2_X1   g607(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n807), .B2(new_n808), .ZN(G1343gat));
  NOR3_X1   g610(.A1(new_n683), .A2(new_n533), .A3(new_n558), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n368), .B2(new_n768), .ZN(new_n815));
  XOR2_X1   g614(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n816));
  OAI21_X1  g615(.A(KEYINPUT119), .B1(new_n775), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n777), .A2(new_n778), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819));
  INV_X1    g618(.A(new_n816), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n776), .A2(new_n402), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n769), .A2(KEYINPUT117), .A3(new_n640), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n815), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n336), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n252), .B1(new_n825), .B2(new_n788), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n498), .B1(new_n826), .B2(new_n791), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n813), .B1(KEYINPUT57), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n792), .A2(new_n498), .A3(new_n797), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G141gat), .B1(new_n832), .B2(new_n403), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n829), .A2(new_n812), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(G141gat), .A3(new_n403), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n832), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n658), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n836), .B1(new_n840), .B2(G141gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n841), .B2(new_n834), .ZN(G1344gat));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n792), .A2(new_n498), .A3(new_n797), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(KEYINPUT120), .A3(new_n830), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n794), .A2(KEYINPUT121), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n787), .A2(new_n847), .A3(new_n335), .A4(new_n334), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n769), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n825), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n253), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n338), .A2(new_n368), .A3(new_n403), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT57), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n498), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n829), .B2(new_n830), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n845), .B1(new_n855), .B2(KEYINPUT120), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n640), .A3(new_n812), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(G148gat), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n857), .B2(new_n858), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n843), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g661(.A(KEYINPUT59), .B(new_n860), .C1(new_n839), .C2(new_n640), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n640), .A2(new_n860), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n862), .A2(new_n863), .B1(new_n835), .B2(new_n864), .ZN(G1345gat));
  INV_X1    g664(.A(new_n478), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n832), .A2(new_n866), .A3(new_n253), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n829), .A2(new_n252), .A3(new_n812), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n866), .B2(new_n868), .ZN(G1346gat));
  INV_X1    g668(.A(new_n479), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n832), .A2(new_n870), .A3(new_n336), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n829), .A2(new_n337), .A3(new_n812), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n870), .B2(new_n872), .ZN(G1347gat));
  AND2_X1   g672(.A1(new_n798), .A2(new_n500), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n598), .A2(new_n559), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G169gat), .B1(new_n876), .B2(new_n403), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n658), .A2(new_n410), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(G1348gat));
  NOR2_X1   g678(.A1(new_n876), .A2(new_n368), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(new_n411), .ZN(G1349gat));
  NOR2_X1   g680(.A1(new_n876), .A2(new_n253), .ZN(new_n882));
  MUX2_X1   g681(.A(G183gat), .B(new_n404), .S(new_n882), .Z(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g683(.A1(new_n874), .A2(new_n337), .A3(new_n875), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G190gat), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(KEYINPUT61), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(KEYINPUT123), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n886), .A2(KEYINPUT124), .A3(KEYINPUT61), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(KEYINPUT123), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT124), .B1(new_n886), .B2(KEYINPUT61), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(G190gat), .B2(new_n885), .ZN(G1351gat));
  NOR2_X1   g692(.A1(new_n830), .A2(KEYINPUT120), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n829), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n875), .A2(new_n603), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n844), .A2(KEYINPUT57), .B1(new_n853), .B2(new_n498), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G197gat), .B1(new_n899), .B2(new_n403), .ZN(new_n900));
  INV_X1    g699(.A(new_n896), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n844), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n385), .A3(new_n658), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(G1352gat));
  INV_X1    g703(.A(new_n902), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(G204gat), .A3(new_n368), .ZN(new_n906));
  XNOR2_X1  g705(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n856), .A2(new_n640), .A3(new_n896), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G204gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1353gat));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n856), .A2(new_n912), .A3(new_n252), .A4(new_n896), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT126), .B1(new_n899), .B2(new_n253), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(G211gat), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n905), .A2(G211gat), .A3(new_n253), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT127), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n919), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1354gat));
  OAI21_X1  g724(.A(G218gat), .B1(new_n899), .B2(new_n336), .ZN(new_n926));
  OR3_X1    g725(.A1(new_n905), .A2(G218gat), .A3(new_n336), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1355gat));
endmodule


