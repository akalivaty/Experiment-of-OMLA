//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1251,
    new_n1252;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n207));
  INV_X1    g0007(.A(G226), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n207), .B1(new_n202), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g0009(.A(new_n209), .B1(G116), .B2(G270), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT65), .Z(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT66), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n211), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n221), .A2(G50), .A3(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n206), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR3_X1   g0029(.A1(new_n220), .A2(new_n226), .A3(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  OAI211_X1 g0049(.A(G1), .B(G13), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT81), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT81), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n253), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n216), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n257), .B(new_n259), .C1(G264), .C2(new_n258), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n252), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G303), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n250), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT5), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n265), .B(G45), .C1(new_n266), .C2(G41), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G274), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT85), .ZN(new_n271));
  INV_X1    g0071(.A(new_n250), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G270), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n264), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G190), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n265), .A2(G20), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G116), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n225), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n285), .B(G116), .C1(G1), .C2(new_n248), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G283), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(new_n224), .C1(G33), .C2(new_n215), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n288), .B(new_n284), .C1(new_n224), .C2(G116), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT20), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n289), .A2(new_n290), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n282), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G200), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n277), .B(new_n294), .C1(new_n295), .C2(new_n276), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G238), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n250), .A2(new_n297), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n252), .A2(new_n261), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G226), .A2(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(G232), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(G1698), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n303), .A2(new_n306), .B1(G33), .B2(G97), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n300), .B1(new_n301), .B2(new_n302), .C1(new_n307), .C2(new_n250), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n308), .A2(KEYINPUT13), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n308), .A2(KEYINPUT13), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT78), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n308), .A2(KEYINPUT78), .A3(KEYINPUT13), .ZN(new_n314));
  OAI211_X1 g0114(.A(G179), .B(new_n310), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(G169), .B1(new_n309), .B2(new_n311), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT14), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n308), .B(KEYINPUT13), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT14), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(G169), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n315), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n202), .A2(G20), .A3(G33), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT79), .ZN(new_n323));
  INV_X1    g0123(.A(G77), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n224), .A2(G33), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n323), .B1(new_n224), .B2(G68), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n284), .B(KEYINPUT70), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n326), .A2(new_n330), .A3(new_n327), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G68), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n280), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g0134(.A(new_n334), .B(KEYINPUT12), .Z(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n285), .A2(G68), .A3(new_n278), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n321), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n338), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n318), .A2(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT77), .ZN(new_n342));
  OAI211_X1 g0142(.A(G190), .B(new_n310), .C1(new_n313), .C2(new_n314), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT77), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n318), .A2(new_n344), .A3(G200), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n340), .A2(new_n342), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT80), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT7), .B1(new_n257), .B2(G20), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT81), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n248), .ZN(new_n351));
  NAND2_X1  g0151(.A1(KEYINPUT81), .A2(G33), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(KEYINPUT3), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n252), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT7), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(new_n224), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n349), .A2(G68), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G58), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n333), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n201), .ZN(new_n360));
  NOR2_X1   g0160(.A1(G20), .A2(G33), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G159), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT82), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n360), .A2(KEYINPUT82), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n357), .A2(new_n367), .A3(KEYINPUT16), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT3), .B1(new_n351), .B2(new_n352), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT83), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n251), .B2(G33), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n248), .A2(KEYINPUT83), .A3(KEYINPUT3), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(KEYINPUT7), .B(new_n224), .C1(new_n370), .C2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n355), .B1(new_n303), .B2(G20), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n333), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n369), .B1(new_n377), .B2(new_n363), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n368), .A2(new_n378), .A3(new_n284), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n358), .A2(KEYINPUT8), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n380), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n358), .A2(KEYINPUT8), .ZN(new_n383));
  MUX2_X1   g0183(.A(new_n380), .B(new_n382), .S(new_n383), .Z(new_n384));
  INV_X1    g0184(.A(new_n278), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n327), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n384), .A2(new_n280), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G223), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n258), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n208), .A2(G1698), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n353), .A2(new_n252), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n272), .ZN(new_n398));
  INV_X1    g0198(.A(G190), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n302), .A2(new_n305), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n398), .A2(new_n399), .A3(new_n300), .A4(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n250), .B1(new_n395), .B2(new_n396), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n403), .A2(new_n299), .A3(new_n400), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n402), .B1(new_n404), .B2(G200), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n379), .A2(new_n391), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT17), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n379), .A2(new_n391), .A3(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n379), .A2(new_n391), .ZN(new_n411));
  INV_X1    g0211(.A(G169), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n299), .B1(new_n397), .B2(new_n272), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(new_n401), .ZN(new_n414));
  INV_X1    g0214(.A(G179), .ZN(new_n415));
  NOR4_X1   g0215(.A1(new_n403), .A2(new_n415), .A3(new_n299), .A4(new_n400), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n411), .A2(KEYINPUT18), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT18), .B1(new_n411), .B2(new_n418), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n408), .B(new_n410), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n303), .A2(G232), .A3(new_n258), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n303), .A2(G238), .A3(G1698), .ZN(new_n424));
  INV_X1    g0224(.A(G107), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n423), .B(new_n424), .C1(new_n425), .C2(new_n303), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n299), .B1(new_n426), .B2(new_n272), .ZN(new_n427));
  INV_X1    g0227(.A(G244), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(new_n302), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT73), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n430), .A2(G169), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n285), .A2(G77), .A3(new_n278), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n280), .A2(new_n324), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT75), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT15), .B(G87), .Z(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n436), .A2(new_n325), .B1(new_n224), .B2(new_n324), .ZN(new_n437));
  INV_X1    g0237(.A(new_n383), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(new_n381), .ZN(new_n439));
  XOR2_X1   g0239(.A(new_n439), .B(KEYINPUT74), .Z(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n440), .B2(new_n361), .ZN(new_n441));
  INV_X1    g0241(.A(new_n284), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n432), .B(new_n434), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n430), .A2(new_n415), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n431), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n348), .A2(new_n422), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n392), .A2(G1698), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(G222), .B2(G1698), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n250), .B1(new_n303), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(G77), .B2(new_n303), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n450), .B(new_n300), .C1(new_n208), .C2(new_n302), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n451), .A2(KEYINPUT69), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(KEYINPUT69), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n452), .A2(KEYINPUT76), .A3(G200), .A4(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n361), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n384), .B2(new_n325), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n327), .ZN(new_n457));
  INV_X1    g0257(.A(new_n280), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n278), .A2(G50), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT72), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n387), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n457), .B(new_n461), .C1(G50), .C2(new_n458), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT9), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n454), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n452), .A2(new_n453), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT76), .B1(new_n466), .B2(new_n399), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(G200), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n462), .A2(new_n463), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT10), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT10), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n473), .A3(new_n470), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n466), .A2(G179), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n466), .A2(new_n412), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n462), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n443), .B1(new_n430), .B2(G190), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n295), .B2(new_n430), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n446), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n276), .A2(G179), .A3(new_n293), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT21), .ZN(new_n484));
  INV_X1    g0284(.A(new_n264), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT85), .ZN(new_n486));
  XNOR2_X1  g0286(.A(new_n270), .B(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n274), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n293), .A2(G169), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n484), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n276), .A2(new_n489), .A3(KEYINPUT21), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n483), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n214), .A2(new_n258), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n216), .A2(G1698), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n353), .A2(new_n252), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G294), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(new_n256), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n272), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n487), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n250), .B(G264), .C1(new_n267), .C2(new_n268), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n501), .B(KEYINPUT88), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n487), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n502), .A2(new_n412), .B1(new_n415), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n425), .A2(G20), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n507), .B(KEYINPUT23), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n353), .A2(KEYINPUT22), .A3(G87), .A4(new_n252), .ZN(new_n509));
  OAI21_X1  g0309(.A(G116), .B1(new_n254), .B2(new_n255), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n511), .B2(new_n224), .ZN(new_n512));
  NOR2_X1   g0312(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n262), .A2(G20), .A3(new_n213), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n515), .A2(KEYINPUT22), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n512), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n512), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n506), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n284), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n387), .B(new_n458), .C1(G1), .C2(new_n248), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G107), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n280), .A2(new_n425), .ZN(new_n524));
  XOR2_X1   g0324(.A(new_n524), .B(KEYINPUT25), .Z(new_n525));
  NAND3_X1  g0325(.A1(new_n520), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n493), .B1(new_n505), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n487), .A2(new_n399), .A3(new_n499), .A4(new_n501), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n504), .A2(new_n295), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(new_n520), .A3(new_n523), .A4(new_n525), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n273), .A2(G257), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n353), .A2(G244), .A3(new_n258), .A4(new_n252), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT4), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n428), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(new_n258), .A3(new_n252), .A4(new_n261), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n252), .A2(new_n261), .A3(G250), .A4(G1698), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n539), .A2(new_n287), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n487), .B(new_n534), .C1(new_n542), .C2(new_n250), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n399), .B2(new_n543), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n280), .A2(new_n215), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n546), .B(KEYINPUT84), .ZN(new_n547));
  XOR2_X1   g0347(.A(G97), .B(G107), .Z(new_n548));
  NAND2_X1  g0348(.A1(new_n425), .A2(G97), .ZN(new_n549));
  MUX2_X1   g0349(.A(new_n548), .B(new_n549), .S(KEYINPUT6), .Z(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n224), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n425), .B1(new_n375), .B2(new_n376), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n324), .A2(G20), .A3(G33), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OAI221_X1 g0354(.A(new_n547), .B1(new_n215), .B2(new_n521), .C1(new_n554), .C2(new_n442), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n545), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G238), .A2(G1698), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n428), .B2(G1698), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n257), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n250), .B1(new_n559), .B2(new_n510), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n265), .A2(G45), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(new_n298), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n250), .A2(G250), .A3(new_n562), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(new_n399), .ZN(new_n567));
  INV_X1    g0367(.A(new_n565), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n560), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(new_n295), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G97), .A2(G107), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n224), .A2(new_n572), .B1(new_n573), .B2(new_n213), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n574), .B(KEYINPUT86), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n224), .A2(G68), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n325), .A2(new_n215), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n354), .A2(new_n576), .B1(KEYINPUT19), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n284), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n436), .A2(new_n280), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(G87), .B2(new_n522), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n569), .A2(G179), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n569), .B2(new_n412), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n579), .B(new_n580), .C1(new_n521), .C2(new_n436), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n571), .A2(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n543), .A2(new_n412), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n250), .B1(new_n537), .B2(new_n541), .ZN(new_n588));
  INV_X1    g0388(.A(new_n534), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n271), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n415), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n555), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  AND4_X1   g0392(.A1(new_n533), .A2(new_n556), .A3(new_n586), .A4(new_n592), .ZN(new_n593));
  AND4_X1   g0393(.A1(new_n296), .A2(new_n482), .A3(new_n527), .A4(new_n593), .ZN(G372));
  AND2_X1   g0394(.A1(new_n526), .A2(new_n505), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT90), .B1(new_n595), .B2(new_n493), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT90), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n527), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT26), .ZN(new_n600));
  INV_X1    g0400(.A(new_n586), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(new_n592), .ZN(new_n602));
  INV_X1    g0402(.A(new_n592), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n586), .A3(KEYINPUT26), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n602), .A2(new_n604), .B1(new_n585), .B2(new_n584), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n482), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n607), .B(KEYINPUT91), .ZN(new_n608));
  INV_X1    g0408(.A(new_n478), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n419), .A2(new_n420), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n445), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(new_n346), .B1(new_n338), .B2(new_n321), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n410), .A2(new_n408), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n609), .B1(new_n615), .B2(new_n475), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n608), .A2(new_n616), .ZN(G369));
  NOR2_X1   g0417(.A1(new_n279), .A2(G20), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n265), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(G213), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(G343), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n595), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n625), .B(KEYINPUT92), .ZN(new_n626));
  INV_X1    g0426(.A(new_n595), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n526), .A2(new_n624), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(new_n533), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n624), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n294), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n493), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n296), .ZN(new_n634));
  INV_X1    g0434(.A(G330), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n627), .A2(new_n624), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n626), .A2(new_n629), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n493), .A2(new_n631), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n644), .ZN(G399));
  INV_X1    g0445(.A(new_n227), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(G41), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR4_X1   g0448(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G1), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n223), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT93), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT28), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n624), .B1(new_n599), .B2(new_n605), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT29), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n593), .B1(new_n595), .B2(new_n493), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n624), .B1(new_n605), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT29), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT30), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n590), .A2(G179), .A3(new_n499), .A4(new_n569), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n276), .A2(new_n503), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n583), .A2(new_n543), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n274), .A2(new_n485), .A3(new_n487), .A4(new_n503), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT30), .A4(new_n499), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n543), .A2(new_n504), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT94), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT94), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n543), .A2(new_n669), .A3(new_n504), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n668), .A2(new_n415), .A3(new_n566), .A4(new_n670), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n663), .B(new_n666), .C1(new_n671), .C2(new_n276), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n624), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT95), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n624), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT31), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n593), .A2(new_n296), .A3(new_n527), .A4(new_n631), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT95), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(new_n677), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n659), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n653), .B1(new_n683), .B2(G1), .ZN(G364));
  NAND2_X1  g0484(.A1(new_n415), .A2(new_n295), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT100), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(G20), .A3(new_n399), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G159), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT32), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n224), .A2(G179), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n399), .A3(G200), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n224), .A2(new_n415), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT99), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n697), .A2(G190), .A3(new_n295), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI221_X1 g0499(.A(new_n303), .B1(new_n425), .B2(new_n695), .C1(new_n699), .C2(new_n358), .ZN(new_n700));
  NOR4_X1   g0500(.A1(new_n224), .A2(new_n399), .A3(new_n295), .A4(G179), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n213), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n696), .A2(G200), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G190), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n704), .A2(new_n399), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n706), .A2(new_n333), .B1(new_n708), .B2(new_n202), .ZN(new_n709));
  NOR4_X1   g0509(.A1(new_n693), .A2(new_n700), .A3(new_n703), .A4(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n697), .A2(new_n399), .A3(new_n295), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n686), .A2(G190), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI221_X1 g0515(.A(new_n710), .B1(new_n324), .B2(new_n712), .C1(new_n215), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT102), .ZN(new_n717));
  INV_X1    g0517(.A(G322), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n699), .A2(new_n718), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n691), .A2(G329), .B1(G326), .B2(new_n707), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT103), .ZN(new_n721));
  INV_X1    g0521(.A(G303), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n262), .B1(new_n702), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g0523(.A(KEYINPUT33), .B(G317), .Z(new_n724));
  OAI221_X1 g0524(.A(new_n720), .B1(new_n721), .B2(new_n723), .C1(new_n706), .C2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(G294), .B2(new_n714), .ZN(new_n726));
  INV_X1    g0526(.A(new_n695), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n711), .A2(G311), .B1(G283), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n723), .A2(new_n721), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n717), .B1(new_n719), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n225), .B1(G20), .B2(new_n412), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n224), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n732), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT98), .Z(new_n737));
  NAND3_X1  g0537(.A1(new_n303), .A2(G355), .A3(new_n227), .ZN(new_n738));
  INV_X1    g0538(.A(G45), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n243), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n257), .A2(new_n646), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G45), .B2(new_n223), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT97), .Z(new_n743));
  OAI221_X1 g0543(.A(new_n738), .B1(G116), .B2(new_n227), .C1(new_n740), .C2(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n731), .A2(new_n732), .B1(new_n737), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n618), .A2(G45), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT96), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(KEYINPUT96), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n747), .A2(G1), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n647), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n634), .A2(new_n735), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n634), .A2(new_n635), .ZN(new_n753));
  INV_X1    g0553(.A(new_n750), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n637), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n752), .A2(new_n755), .ZN(G396));
  NOR2_X1   g0556(.A1(new_n445), .A2(new_n624), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n443), .A2(new_n624), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n480), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n757), .B1(new_n759), .B2(new_n445), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n654), .B(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(new_n682), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n754), .ZN(new_n763));
  INV_X1    g0563(.A(new_n760), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n733), .ZN(new_n765));
  AOI22_X1  g0565(.A1(G143), .A2(new_n698), .B1(new_n711), .B2(G159), .ZN(new_n766));
  INV_X1    g0566(.A(G137), .ZN(new_n767));
  INV_X1    g0567(.A(G150), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n766), .B1(new_n767), .B2(new_n708), .C1(new_n768), .C2(new_n706), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT34), .Z(new_n770));
  NOR2_X1   g0570(.A1(new_n702), .A2(new_n202), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n715), .A2(new_n358), .ZN(new_n772));
  INV_X1    g0572(.A(G132), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n257), .B1(new_n333), .B2(new_n695), .C1(new_n690), .C2(new_n773), .ZN(new_n774));
  NOR4_X1   g0574(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n699), .A2(new_n497), .B1(new_n425), .B2(new_n702), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n695), .A2(new_n213), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n776), .A2(new_n303), .A3(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n715), .A2(new_n215), .B1(new_n722), .B2(new_n708), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G283), .B2(new_n705), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n691), .A2(G311), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G116), .B2(new_n711), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n732), .B1(new_n775), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n732), .A2(new_n733), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n324), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n765), .A2(new_n750), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n763), .A2(new_n787), .ZN(G384));
  INV_X1    g0588(.A(KEYINPUT110), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n673), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n672), .A2(KEYINPUT110), .A3(KEYINPUT31), .A4(new_n624), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n679), .A2(new_n790), .A3(new_n677), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n338), .A2(new_n624), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n339), .A2(new_n346), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n321), .A2(new_n338), .A3(new_n624), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT104), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n794), .A2(KEYINPUT104), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n792), .A2(new_n800), .A3(new_n760), .ZN(new_n801));
  INV_X1    g0601(.A(new_n622), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n357), .A2(new_n367), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n387), .B1(new_n803), .B2(new_n369), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n390), .B1(new_n804), .B2(new_n368), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n421), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT107), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n622), .B1(new_n379), .B2(new_n391), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n409), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n411), .A2(new_n418), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT106), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n417), .B1(new_n391), .B2(new_n379), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(KEYINPUT106), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n810), .A2(new_n813), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n414), .A2(new_n416), .A3(new_n802), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n406), .B1(new_n805), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT105), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT37), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n820), .B1(new_n819), .B2(KEYINPUT37), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n808), .B(new_n817), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n355), .B1(new_n354), .B2(new_n224), .ZN(new_n826));
  AOI211_X1 g0626(.A(KEYINPUT7), .B(G20), .C1(new_n353), .C2(new_n252), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n826), .A2(new_n827), .A3(new_n333), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n365), .A2(new_n366), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n369), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n830), .A2(new_n327), .A3(new_n368), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n831), .A2(new_n391), .B1(new_n417), .B2(new_n622), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT37), .B1(new_n832), .B2(new_n409), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT105), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n821), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n808), .B1(new_n835), .B2(new_n817), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n807), .B1(new_n825), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(KEYINPUT38), .B(new_n807), .C1(new_n825), .C2(new_n836), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n801), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(KEYINPUT40), .ZN(new_n842));
  AND3_X1   g0642(.A1(new_n792), .A2(new_n800), .A3(new_n760), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n814), .A2(new_n409), .A3(new_n809), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n817), .B1(new_n816), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n421), .A2(new_n809), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n838), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n843), .A2(new_n849), .A3(KEYINPUT40), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n842), .A2(new_n482), .A3(new_n792), .A4(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n850), .B(G330), .C1(new_n841), .C2(KEYINPUT40), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n446), .A2(new_n481), .A3(new_n635), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n792), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n851), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n655), .A2(new_n482), .A3(new_n658), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n616), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n857), .B(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT39), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n839), .B2(new_n840), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n840), .A2(new_n861), .A3(new_n848), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT108), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n817), .B1(new_n822), .B2(new_n823), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT107), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n824), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n867), .B2(new_n807), .ZN(new_n868));
  INV_X1    g0668(.A(new_n807), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n838), .B(new_n869), .C1(new_n866), .C2(new_n824), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT39), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT108), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n840), .A2(new_n861), .A3(new_n848), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n864), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n339), .A2(new_n624), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n757), .B1(new_n654), .B2(new_n760), .ZN(new_n878));
  INV_X1    g0678(.A(new_n800), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n839), .A2(new_n840), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n880), .A2(new_n881), .B1(new_n610), .B2(new_n622), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n877), .A2(KEYINPUT109), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT109), .ZN(new_n884));
  INV_X1    g0684(.A(new_n876), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n864), .B2(new_n874), .ZN(new_n886));
  INV_X1    g0686(.A(new_n882), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n860), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n265), .B2(new_n618), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT35), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n224), .B(new_n225), .C1(new_n550), .C2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n893), .B(G116), .C1(new_n892), .C2(new_n550), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n223), .A2(new_n324), .A3(new_n359), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n333), .A2(G50), .ZN(new_n897));
  OAI211_X1 g0697(.A(G1), .B(new_n279), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n891), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT111), .Z(G367));
  NAND2_X1  g0700(.A1(new_n641), .A2(new_n643), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n555), .A2(new_n624), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n556), .A2(new_n592), .A3(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT113), .Z(new_n904));
  NAND2_X1  g0704(.A1(new_n603), .A2(new_n624), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  OR3_X1    g0707(.A1(new_n901), .A2(KEYINPUT42), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n592), .B1(new_n904), .B2(new_n627), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n631), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT42), .B1(new_n901), .B2(new_n907), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n586), .B1(new_n582), .B2(new_n631), .ZN(new_n913));
  INV_X1    g0713(.A(new_n582), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n914), .A2(new_n584), .A3(new_n585), .A4(new_n624), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT112), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n912), .A2(new_n917), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n922), .B2(new_n912), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n639), .A2(new_n907), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n647), .B(KEYINPUT41), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT44), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n644), .B2(new_n906), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n642), .B1(new_n626), .B2(new_n629), .ZN(new_n931));
  OAI211_X1 g0731(.A(KEYINPUT44), .B(new_n907), .C1(new_n931), .C2(new_n640), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n644), .A2(KEYINPUT45), .A3(new_n906), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT45), .B1(new_n644), .B2(new_n906), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n638), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n641), .B(new_n642), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(new_n636), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n636), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n933), .B(new_n639), .C1(new_n934), .C2(new_n935), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n937), .A2(new_n942), .A3(new_n683), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n928), .B1(new_n944), .B2(new_n683), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n926), .B1(new_n945), .B2(new_n749), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n303), .B1(new_n699), .B2(new_n768), .C1(new_n202), .C2(new_n712), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n691), .A2(G137), .B1(G77), .B2(new_n727), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n714), .A2(G68), .B1(G143), .B2(new_n707), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(new_n358), .C2(new_n702), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n947), .B(new_n950), .C1(G159), .C2(new_n705), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n702), .A2(new_n281), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(KEYINPUT46), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G311), .B2(new_n707), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n257), .B1(new_n711), .B2(G283), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(new_n497), .C2(new_n706), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n698), .A2(G303), .B1(KEYINPUT46), .B2(new_n952), .ZN(new_n957));
  INV_X1    g0757(.A(G317), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n957), .B1(new_n215), .B2(new_n695), .C1(new_n690), .C2(new_n958), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n956), .B(new_n959), .C1(G107), .C2(new_n714), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n951), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT47), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n732), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n913), .A2(new_n735), .A3(new_n915), .ZN(new_n964));
  INV_X1    g0764(.A(new_n741), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n736), .B1(new_n227), .B2(new_n436), .C1(new_n965), .C2(new_n238), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n963), .A2(new_n750), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n946), .A2(new_n967), .ZN(G387));
  NOR2_X1   g0768(.A1(new_n384), .A2(new_n706), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n727), .A2(G97), .B1(new_n701), .B2(G77), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n257), .B(new_n970), .C1(new_n690), .C2(new_n768), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT116), .Z(new_n972));
  AOI22_X1  g0772(.A1(new_n714), .A2(new_n435), .B1(G159), .B2(new_n707), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(new_n202), .C2(new_n699), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n969), .B(new_n974), .C1(G68), .C2(new_n711), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT117), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G303), .A2(new_n711), .B1(new_n698), .B2(G317), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n718), .B2(new_n708), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G311), .B2(new_n705), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT48), .Z(new_n980));
  INV_X1    g0780(.A(G283), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n980), .B1(new_n981), .B2(new_n715), .C1(new_n497), .C2(new_n702), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT49), .Z(new_n983));
  INV_X1    g0783(.A(G326), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n354), .B1(new_n281), .B2(new_n695), .C1(new_n690), .C2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n976), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n986), .A2(new_n732), .B1(new_n630), .B2(new_n735), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n235), .A2(new_n739), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT114), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n440), .A2(new_n202), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(G45), .B1(G68), .B2(G77), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n992), .A2(new_n649), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n741), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n303), .A2(new_n227), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(G107), .B2(new_n227), .C1(new_n649), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n737), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n987), .A2(new_n750), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT118), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n942), .A2(new_n683), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n941), .B1(new_n682), .B2(new_n659), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1001), .A2(new_n647), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n942), .A2(new_n749), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1000), .A2(new_n1003), .A3(new_n1004), .ZN(G393));
  AOI21_X1  g0805(.A(new_n754), .B1(new_n907), .B2(new_n735), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n702), .A2(new_n981), .B1(new_n425), .B2(new_n695), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n303), .B(new_n1007), .C1(new_n691), .C2(G322), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT119), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n711), .A2(G294), .B1(G303), .B2(new_n705), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n698), .A2(G311), .B1(G317), .B2(new_n707), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT52), .Z(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G116), .B2(new_n714), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n698), .A2(G159), .B1(G150), .B2(new_n707), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT51), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n714), .A2(G77), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n440), .A2(new_n711), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n701), .A2(G68), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n257), .B1(new_n706), .B2(new_n202), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n691), .A2(G143), .ZN(new_n1022));
  NOR4_X1   g0822(.A1(new_n1020), .A2(new_n777), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n732), .B1(new_n1014), .B2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n736), .B1(new_n215), .B2(new_n227), .C1(new_n965), .C2(new_n246), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1006), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n937), .A2(new_n943), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n749), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n648), .B1(new_n1027), .B2(new_n1001), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1029), .B1(new_n944), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(G390));
  OAI21_X1  g0832(.A(new_n885), .B1(new_n878), .B2(new_n879), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n864), .A2(new_n874), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n682), .A2(new_n760), .A3(new_n800), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n759), .A2(new_n445), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n757), .B1(new_n657), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n849), .B(new_n885), .C1(new_n1037), .C2(new_n879), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1034), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n843), .A2(G330), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n858), .A2(new_n855), .A3(new_n616), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n792), .A2(G330), .A3(new_n760), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n879), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT120), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(KEYINPUT120), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1046), .A2(new_n1035), .A3(new_n1037), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n878), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n681), .A2(G330), .A3(new_n760), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1050), .A2(new_n879), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1040), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1043), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n648), .B1(new_n1042), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1054), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1042), .A2(new_n749), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n864), .A2(new_n874), .A3(new_n733), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT53), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n702), .A2(new_n768), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n691), .A2(G125), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT54), .B(G143), .Z(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1063), .B1(new_n1061), .B2(new_n1062), .C1(new_n712), .C2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n706), .A2(new_n767), .ZN(new_n1067));
  INV_X1    g0867(.A(G159), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n715), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n707), .A2(G128), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n262), .B1(new_n727), .B2(G50), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n699), .C2(new_n773), .ZN(new_n1072));
  NOR4_X1   g0872(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .A4(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n262), .B1(new_n708), .B2(new_n981), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n691), .A2(G294), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n711), .A2(G97), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n714), .A2(G77), .B1(G107), .B2(new_n705), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n703), .B1(G68), .B2(new_n727), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1074), .B(new_n1079), .C1(G116), .C2(new_n698), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n732), .B1(new_n1073), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n384), .A2(new_n785), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1060), .A2(new_n750), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1058), .A2(new_n1059), .A3(new_n1083), .ZN(G378));
  INV_X1    g0884(.A(KEYINPUT57), .ZN(new_n1085));
  XOR2_X1   g0885(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n469), .A2(new_n473), .A3(new_n470), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n473), .B1(new_n469), .B2(new_n470), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n478), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT55), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n475), .A2(KEYINPUT55), .A3(new_n478), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n462), .A2(new_n802), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1094), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1087), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1094), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n1086), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n852), .B(new_n1103), .Z(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT109), .B1(new_n877), .B2(new_n882), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n886), .A2(new_n887), .A3(new_n884), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n852), .B(new_n1103), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n883), .A2(new_n1108), .A3(new_n888), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1043), .B1(new_n1042), .B2(new_n1054), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1085), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1052), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1034), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n1115), .A3(new_n1054), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1043), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1118), .A2(KEYINPUT57), .A3(new_n1109), .A4(new_n1107), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1112), .A2(new_n647), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1107), .A2(new_n749), .A3(new_n1109), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1097), .A2(new_n1102), .A3(new_n733), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G107), .A2(new_n698), .B1(new_n714), .B2(G68), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n215), .B2(new_n706), .C1(new_n690), .C2(new_n981), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G58), .B2(new_n727), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n354), .B1(new_n702), .B2(new_n324), .C1(new_n708), .C2(new_n281), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n711), .B2(new_n435), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n249), .A3(new_n1127), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT58), .Z(new_n1129));
  OAI22_X1  g0929(.A1(new_n712), .A2(new_n767), .B1(new_n702), .B2(new_n1065), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G128), .B2(new_n698), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G125), .A2(new_n707), .B1(new_n705), .B2(G132), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n768), .C2(new_n715), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT59), .ZN(new_n1134));
  AOI21_X1  g0934(.A(G33), .B1(new_n727), .B2(G159), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n249), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n691), .B2(G124), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT121), .ZN(new_n1138));
  AOI21_X1  g0938(.A(G41), .B1(new_n254), .B2(KEYINPUT3), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1134), .A2(new_n1138), .B1(G50), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n732), .B1(new_n1129), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n785), .A2(new_n202), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1122), .A2(new_n750), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1121), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1120), .A2(new_n1145), .ZN(G375));
  NAND3_X1  g0946(.A1(new_n1048), .A2(new_n1053), .A3(new_n1043), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1056), .A2(new_n927), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1028), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n879), .A2(new_n733), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n691), .A2(G128), .B1(new_n705), .B2(new_n1064), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n358), .B2(new_n695), .C1(new_n768), .C2(new_n712), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n708), .A2(new_n773), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n715), .A2(new_n202), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n257), .B1(new_n1068), .B2(new_n702), .C1(new_n699), .C2(new_n767), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n691), .A2(G303), .B1(G77), .B2(new_n727), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n981), .B2(new_n699), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n706), .A2(new_n281), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n714), .A2(new_n435), .B1(G294), .B2(new_n707), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n712), .B2(new_n425), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n262), .B1(new_n702), .B2(new_n215), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n732), .B1(new_n1156), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n785), .A2(new_n333), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1150), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1149), .B1(new_n750), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1148), .A2(new_n1167), .ZN(G381));
  NOR2_X1   g0968(.A1(G375), .A2(G378), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1170), .A2(G384), .A3(G381), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n946), .A2(new_n1031), .A3(new_n967), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1172), .A2(G396), .A3(G393), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1173), .ZN(G407));
  OAI211_X1 g0974(.A(G407), .B(G213), .C1(G343), .C2(new_n1170), .ZN(G409));
  XNOR2_X1  g0975(.A(G393), .B(G396), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1172), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1031), .B1(new_n946), .B2(new_n967), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1179), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(G375), .A2(G378), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT62), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT60), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1147), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1147), .A2(new_n1186), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1187), .A2(new_n647), .A3(new_n1056), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1167), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT123), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(G384), .B(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n763), .A2(new_n1191), .A3(new_n787), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1190), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(G213), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(G343), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1118), .A2(new_n927), .A3(new_n1109), .A4(new_n1107), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1201), .A2(new_n1121), .A3(new_n1143), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1059), .A2(new_n1083), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1057), .B2(new_n1055), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1200), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1184), .A2(new_n1185), .A3(new_n1198), .A4(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT125), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1184), .B2(new_n1205), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1204), .B1(new_n1120), .B2(new_n1145), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1201), .A2(new_n1121), .A3(new_n1143), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n1211), .A2(G378), .B1(new_n1199), .B2(G343), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1210), .A2(new_n1212), .A3(KEYINPUT125), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1198), .B1(new_n1209), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1207), .B1(new_n1214), .B2(KEYINPUT62), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1118), .A2(new_n1109), .A3(new_n1107), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n648), .B1(new_n1216), .B2(new_n1085), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1144), .B1(new_n1217), .B2(new_n1119), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1205), .B(new_n1208), .C1(new_n1204), .C2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(KEYINPUT125), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1200), .A2(G2897), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1221), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1193), .B(new_n1223), .C1(new_n1195), .C2(new_n1190), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1219), .A2(new_n1220), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n1228));
  OR2_X1    g1028(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1183), .B1(new_n1215), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT61), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1180), .A2(new_n1182), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT124), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1233), .B(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1197), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT63), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1184), .A2(new_n1198), .A3(new_n1205), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1225), .B1(new_n1184), .B2(new_n1205), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT63), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1235), .A2(new_n1237), .A3(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(KEYINPUT127), .B1(new_n1231), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT127), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1235), .A2(new_n1237), .A3(new_n1241), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1206), .B1(new_n1236), .B2(new_n1185), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1244), .B(new_n1245), .C1(new_n1248), .C2(new_n1183), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1243), .A2(new_n1249), .ZN(G405));
  XNOR2_X1  g1050(.A(new_n1183), .B(new_n1198), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1170), .A2(new_n1184), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1251), .B(new_n1252), .ZN(G402));
endmodule


