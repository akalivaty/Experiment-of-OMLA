//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n457), .A2(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(G137), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(G2104), .ZN(new_n473));
  OAI22_X1  g048(.A1(new_n466), .A2(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI221_X1 g051(.A(KEYINPUT71), .B1(new_n472), .B2(new_n473), .C1(new_n466), .C2(new_n471), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n469), .A2(new_n470), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n482), .A2(new_n463), .A3(KEYINPUT68), .ZN(new_n483));
  AOI21_X1  g058(.A(KEYINPUT68), .B1(new_n482), .B2(new_n463), .ZN(new_n484));
  OAI21_X1  g059(.A(G125), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(G113), .A2(G2104), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n481), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n479), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G160));
  NOR2_X1   g066(.A1(new_n466), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  INV_X1    g068(.A(G124), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n481), .A2(new_n466), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G112), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n480), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n501));
  OAI221_X1 g076(.A(new_n493), .B1(new_n494), .B2(new_n495), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G162));
  NAND4_X1  g078(.A1(new_n462), .A2(new_n465), .A3(G126), .A4(new_n463), .ZN(new_n504));
  NAND2_X1  g079(.A1(G114), .A2(G2104), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n468), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n473), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G102), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n461), .A2(G2104), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n482), .A2(new_n463), .A3(KEYINPUT68), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n469), .A2(KEYINPUT73), .A3(G138), .A4(new_n470), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n469), .A2(G138), .A3(new_n470), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT4), .B1(new_n466), .B2(new_n521), .ZN(new_n522));
  AOI211_X1 g097(.A(new_n506), .B(new_n509), .C1(new_n520), .C2(new_n522), .ZN(G164));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n526), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n528), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G168));
  INV_X1    g117(.A(new_n526), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G90), .ZN(new_n544));
  INV_X1    g119(.A(new_n528), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G52), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n544), .B(new_n546), .C1(new_n532), .C2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n526), .A2(new_n550), .B1(new_n528), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n532), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND3_X1  g135(.A1(new_n524), .A2(G53), .A3(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n543), .A2(G91), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n532), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(G299));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n543), .A2(G87), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n545), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n525), .A2(G61), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT74), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT75), .ZN(new_n578));
  INV_X1    g153(.A(new_n576), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n532), .B1(new_n579), .B2(new_n573), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n526), .A2(new_n583), .B1(new_n528), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n578), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n578), .A2(new_n582), .A3(new_n590), .A4(new_n586), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n526), .A2(new_n595), .B1(new_n528), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n532), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n543), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n526), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(new_n525), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT77), .B(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(new_n545), .B2(G54), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n602), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n602), .B1(new_n614), .B2(G868), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  XOR2_X1   g194(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  NOR2_X1   g197(.A1(new_n555), .A2(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n614), .A2(new_n621), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n515), .A2(new_n507), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n628), .B(new_n629), .Z(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT82), .Z(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n495), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  INV_X1    g215(.A(G111), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n640), .B1(new_n480), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n492), .B2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  INV_X1    g220(.A(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(new_n646), .A3(new_n643), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n632), .A2(new_n633), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n635), .A2(new_n645), .A3(new_n647), .A4(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT14), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n655), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(new_n664), .A3(G14), .ZN(G401));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT17), .Z(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  INV_X1    g246(.A(new_n668), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(new_n666), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n670), .B(new_n671), .C1(new_n669), .C2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n666), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT18), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(new_n646), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2100), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT84), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT85), .B(G1981), .Z(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(G229));
  NAND2_X1  g273(.A1(new_n593), .A2(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G6), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1971), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(G288), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n704), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT33), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(G1976), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(G1976), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n707), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n702), .A2(new_n703), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n702), .A2(new_n714), .A3(new_n717), .A4(new_n703), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n492), .A2(G131), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  INV_X1    g297(.A(G107), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n480), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n481), .A2(new_n466), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(G119), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G29), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G25), .B2(G29), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT35), .B(G1991), .Z(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n704), .A2(G24), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n600), .B2(new_n704), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1986), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n732), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n716), .A2(new_n718), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(KEYINPUT36), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n716), .A2(new_n740), .A3(new_n718), .A4(new_n737), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n704), .A2(G21), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G168), .B2(new_n704), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G1966), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n704), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n555), .B2(new_n704), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n745), .B1(G1341), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G33), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT25), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n515), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(new_n481), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n752), .B(new_n754), .C1(G139), .C2(new_n492), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n750), .B1(new_n755), .B2(new_n749), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n748), .B1(G1341), .B2(new_n747), .C1(new_n756), .C2(G2072), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(G2072), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n704), .A2(G4), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n614), .B2(new_n704), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT87), .B(G1348), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n760), .B(new_n762), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n757), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n749), .A2(G35), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G162), .B2(new_n749), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT29), .B(G2090), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n704), .A2(G20), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n618), .B2(new_n704), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n768), .A2(new_n769), .A3(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n764), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n749), .A2(G27), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G164), .B2(new_n749), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT93), .B(G2078), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n749), .A2(G32), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n492), .A2(G141), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT89), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n725), .A2(G129), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G105), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n473), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n783), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n781), .B1(new_n790), .B2(new_n749), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT27), .B(G1996), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT91), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT92), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n704), .A2(G5), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G171), .B2(new_n704), .ZN(new_n797));
  INV_X1    g372(.A(G1961), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT30), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n800), .A2(G28), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n749), .B1(new_n800), .B2(G28), .ZN(new_n802));
  AND2_X1   g377(.A1(KEYINPUT31), .A2(G11), .ZN(new_n803));
  NOR2_X1   g378(.A1(KEYINPUT31), .A2(G11), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n801), .A2(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n744), .B2(G1966), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n799), .B(new_n806), .C1(new_n749), .C2(new_n644), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n749), .A2(G26), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT28), .ZN(new_n809));
  OAI221_X1 g384(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n481), .C2(G116), .ZN(new_n810));
  INV_X1    g385(.A(G128), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n495), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G140), .B2(new_n492), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n809), .B1(new_n813), .B2(new_n749), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G2067), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n807), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n749), .B1(KEYINPUT24), .B2(G34), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(KEYINPUT24), .B2(G34), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n490), .B2(G29), .ZN(new_n819));
  INV_X1    g394(.A(G2084), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT88), .Z(new_n822));
  AOI22_X1  g397(.A1(new_n791), .A2(new_n793), .B1(new_n820), .B2(new_n819), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n816), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NOR4_X1   g399(.A1(new_n776), .A2(new_n780), .A3(new_n795), .A4(new_n824), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n742), .A2(KEYINPUT94), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(KEYINPUT94), .B1(new_n742), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(G311));
  NAND2_X1  g403(.A1(new_n742), .A2(new_n825), .ZN(G150));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  INV_X1    g405(.A(G55), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n526), .A2(new_n830), .B1(new_n528), .B2(new_n831), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n532), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n555), .B(new_n835), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n614), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n836), .B1(new_n844), .B2(KEYINPUT39), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n838), .B1(new_n845), .B2(new_n846), .ZN(G145));
  OAI21_X1  g422(.A(new_n519), .B1(new_n483), .B2(new_n484), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n516), .A2(new_n517), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n522), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n506), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n851), .A3(new_n508), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n790), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n790), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n813), .B(KEYINPUT96), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n813), .B(KEYINPUT96), .Z(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(new_n853), .A3(new_n854), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n755), .B2(KEYINPUT97), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n861), .B2(new_n755), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n864), .A2(new_n857), .A3(new_n859), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n725), .A2(G130), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT99), .Z(new_n869));
  INV_X1    g444(.A(G118), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT100), .B1(new_n480), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n480), .A2(KEYINPUT100), .A3(new_n870), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n873), .A2(new_n874), .B1(G142), .B2(new_n492), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n728), .ZN(new_n877));
  INV_X1    g452(.A(new_n630), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n876), .B(new_n727), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n630), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n881), .A3(KEYINPUT101), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n881), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n866), .A2(new_n867), .A3(new_n882), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n863), .A2(new_n865), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT102), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n882), .A2(new_n885), .B1(new_n863), .B2(new_n865), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n502), .B(new_n490), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n644), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n863), .A2(new_n865), .A3(new_n883), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n897), .A2(new_n894), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n898), .B2(new_n891), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n896), .A2(KEYINPUT40), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT40), .B1(new_n896), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(G395));
  NOR2_X1   g477(.A1(new_n835), .A2(G868), .ZN(new_n903));
  AOI21_X1  g478(.A(G290), .B1(new_n588), .B2(new_n591), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(G166), .B(G288), .Z(new_n906));
  NAND3_X1  g481(.A1(new_n588), .A2(new_n591), .A3(G290), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n906), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n588), .A2(new_n591), .A3(G290), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(new_n904), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n618), .A2(new_n613), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT103), .B1(new_n618), .B2(new_n613), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n618), .A2(new_n613), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n918), .B2(new_n921), .ZN(new_n924));
  NOR4_X1   g499(.A1(new_n917), .A2(new_n919), .A3(KEYINPUT41), .A4(new_n920), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n839), .B(new_n624), .ZN(new_n927));
  MUX2_X1   g502(.A(new_n922), .B(new_n926), .S(new_n927), .Z(new_n928));
  OR2_X1    g503(.A1(new_n914), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n914), .A2(new_n928), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n930), .A3(G868), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n903), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n932), .B2(new_n931), .ZN(G295));
  OAI21_X1  g509(.A(new_n933), .B1(new_n932), .B2(new_n931), .ZN(G331));
  XNOR2_X1  g510(.A(G301), .B(G168), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n839), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(new_n924), .B2(new_n925), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n839), .A2(new_n936), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n839), .A2(new_n936), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n939), .A2(new_n918), .A3(new_n921), .A4(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n912), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n912), .A3(new_n941), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n945));
  INV_X1    g520(.A(G37), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n944), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(new_n946), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n950), .B2(new_n942), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(KEYINPUT44), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n953));
  INV_X1    g528(.A(new_n942), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n947), .B2(new_n948), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n943), .A2(new_n946), .A3(new_n944), .ZN(new_n957));
  AOI211_X1 g532(.A(new_n953), .B(KEYINPUT44), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n950), .A2(KEYINPUT106), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n942), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n957), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT107), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n952), .B1(new_n958), .B2(new_n965), .ZN(G397));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n852), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n479), .A2(G40), .A3(new_n489), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n790), .B(G1996), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n813), .B(G2067), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n728), .A2(new_n731), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n728), .A2(new_n731), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n600), .B(G1986), .Z(new_n978));
  OAI21_X1  g553(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(KEYINPUT108), .Z(new_n980));
  INV_X1    g555(.A(G40), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n478), .A2(new_n488), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n509), .B1(new_n520), .B2(new_n522), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n983), .B2(new_n851), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n984), .B2(KEYINPUT45), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n852), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT109), .B(G1971), .Z(new_n989));
  OAI21_X1  g564(.A(KEYINPUT110), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT45), .B1(new_n852), .B2(new_n967), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(new_n971), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n992), .B2(new_n986), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n968), .A2(KEYINPUT50), .ZN(new_n996));
  INV_X1    g571(.A(G2090), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n852), .A2(new_n967), .A3(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n982), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n990), .B(new_n995), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G303), .A2(G8), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1006));
  XNOR2_X1  g581(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(G8), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n984), .A2(new_n982), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G8), .ZN(new_n1010));
  OAI21_X1  g585(.A(G1981), .B1(new_n580), .B2(new_n585), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n587), .B2(G1981), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1010), .B1(KEYINPUT49), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(KEYINPUT49), .B2(new_n1014), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1010), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(G288), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1017), .B(new_n1019), .C1(new_n1018), .C2(G288), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G288), .A2(new_n1018), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n1010), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1016), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n587), .A2(G1981), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G288), .A2(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1016), .B2(new_n1025), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n1008), .A2(new_n1023), .B1(new_n1010), .B2(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1016), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1028));
  NOR2_X1   g603(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT115), .B1(G164), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n852), .A2(new_n1032), .A3(new_n1029), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n982), .B1(new_n984), .B2(new_n998), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1034), .A2(new_n1035), .A3(G2090), .ZN(new_n1036));
  OAI21_X1  g611(.A(G8), .B1(new_n1036), .B2(new_n993), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1007), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n991), .B2(new_n971), .ZN(new_n1041));
  OAI211_X1 g616(.A(KEYINPUT116), .B(new_n982), .C1(new_n984), .C2(KEYINPUT45), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1042), .A3(new_n986), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n999), .A2(new_n982), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n984), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1043), .A2(new_n1044), .B1(new_n1048), .B2(new_n820), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1049), .A2(new_n1050), .A3(G286), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1008), .A2(new_n1028), .A3(new_n1039), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT63), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1004), .A2(G8), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1038), .ZN(new_n1056));
  NOR4_X1   g631(.A1(new_n1049), .A2(new_n1053), .A3(new_n1050), .A4(G286), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(new_n1008), .A3(new_n1028), .A4(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1027), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n773), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G299), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT57), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT56), .B(G2072), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n992), .A2(new_n986), .A3(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1060), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1048), .A2(new_n762), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1009), .A2(G2067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n614), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1063), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1033), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1032), .B1(new_n852), .B2(new_n1029), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n998), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n971), .B1(new_n968), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1956), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1064), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n985), .A2(new_n987), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1070), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1066), .B1(new_n1069), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n996), .A2(new_n982), .A3(new_n999), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1068), .B1(new_n1081), .B2(new_n761), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT60), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n614), .A2(KEYINPUT120), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n613), .B(KEYINPUT120), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(KEYINPUT60), .A3(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1082), .A2(KEYINPUT60), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1063), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1090), .B1(new_n1066), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1060), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1079), .A2(KEYINPUT61), .A3(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n971), .B2(new_n968), .ZN(new_n1096));
  INV_X1    g671(.A(G1996), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n986), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n985), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n555), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT118), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1102), .A3(new_n555), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(KEYINPUT59), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  INV_X1    g680(.A(new_n555), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n970), .A2(new_n1097), .A3(new_n982), .A4(new_n986), .ZN(new_n1107));
  AOI211_X1 g682(.A(KEYINPUT118), .B(new_n1106), .C1(new_n1107), .C2(new_n1096), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1102), .B1(new_n1099), .B2(new_n555), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1105), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1092), .A2(new_n1094), .A3(new_n1104), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1089), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(KEYINPUT119), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1080), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT121), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT51), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1050), .B1(new_n1049), .B2(G168), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1049), .A2(G168), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT51), .B(new_n1117), .C1(new_n1121), .C2(new_n1050), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1049), .A2(new_n1050), .A3(G168), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G2078), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n970), .A2(new_n1126), .A3(new_n982), .A4(new_n986), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1081), .A2(new_n798), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1128), .A2(G2078), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1041), .A2(new_n1042), .A3(new_n986), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(G171), .ZN(new_n1135));
  OR2_X1    g710(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1136));
  NAND2_X1  g711(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1137));
  AOI211_X1 g712(.A(new_n1128), .B(new_n981), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n479), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n485), .A2(new_n487), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1141), .A2(KEYINPUT122), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n481), .B1(new_n1141), .B2(KEYINPUT122), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(new_n970), .A3(new_n986), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1129), .A2(new_n1130), .A3(new_n1145), .ZN(new_n1146));
  OR3_X1    g721(.A1(new_n1146), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT124), .B1(new_n1146), .B2(G171), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1135), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT54), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1146), .A2(G171), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1129), .A2(new_n1133), .A3(G301), .A4(new_n1130), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(KEYINPUT54), .A3(new_n1153), .ZN(new_n1154));
  AND4_X1   g729(.A1(new_n1039), .A2(new_n1008), .A3(new_n1154), .A4(new_n1028), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1125), .A2(new_n1151), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1059), .B1(new_n1116), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1123), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n1122), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1158), .B2(new_n1122), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1135), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1162), .A2(new_n1039), .A3(new_n1008), .A4(new_n1028), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n980), .B1(new_n1157), .B2(new_n1164), .ZN(new_n1165));
  NOR4_X1   g740(.A1(new_n970), .A2(new_n971), .A3(G1986), .A4(G290), .ZN(new_n1166));
  XNOR2_X1  g741(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n977), .A2(new_n972), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1168), .B1(new_n1169), .B2(KEYINPUT126), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(KEYINPUT126), .B2(new_n1169), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n974), .A2(new_n790), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n972), .A2(new_n1097), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT46), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1172), .A2(new_n972), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n1174), .B2(new_n1173), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT47), .Z(new_n1177));
  INV_X1    g752(.A(G2067), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n813), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n975), .B(KEYINPUT125), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n973), .A2(new_n974), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g757(.A(new_n1171), .B(new_n1177), .C1(new_n972), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1165), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g759(.A1(new_n896), .A2(new_n899), .ZN(new_n1186));
  INV_X1    g760(.A(G319), .ZN(new_n1187));
  NOR4_X1   g761(.A1(G229), .A2(new_n1187), .A3(G401), .A4(G227), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n1186), .A2(new_n963), .A3(new_n1188), .ZN(G225));
  INV_X1    g763(.A(G225), .ZN(G308));
endmodule


