

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750;

  BUF_X1 U372 ( .A(n447), .Z(n350) );
  NOR2_X1 U373 ( .A1(n579), .A2(n667), .ZN(n620) );
  XNOR2_X1 U374 ( .A(n509), .B(n349), .ZN(n507) );
  XNOR2_X1 U375 ( .A(n467), .B(n504), .ZN(n349) );
  XNOR2_X1 U376 ( .A(n473), .B(n472), .ZN(n513) );
  XNOR2_X1 U377 ( .A(G107), .B(G104), .ZN(n501) );
  INV_X2 U378 ( .A(G953), .ZN(n741) );
  NOR2_X1 U379 ( .A1(n750), .A2(n749), .ZN(n575) );
  XNOR2_X1 U380 ( .A(n573), .B(KEYINPUT40), .ZN(n750) );
  XNOR2_X1 U381 ( .A(KEYINPUT93), .B(G110), .ZN(n426) );
  NOR2_X1 U382 ( .A1(n674), .A2(n617), .ZN(n679) );
  NOR2_X1 U383 ( .A1(n569), .A2(n598), .ZN(n656) );
  NOR2_X2 U384 ( .A1(n598), .A2(n597), .ZN(n425) );
  XNOR2_X2 U385 ( .A(n401), .B(KEYINPUT4), .ZN(n510) );
  NAND2_X1 U386 ( .A1(n661), .A2(n647), .ZN(n624) );
  NOR2_X1 U387 ( .A1(n599), .A2(n667), .ZN(n374) );
  INV_X1 U388 ( .A(KEYINPUT34), .ZN(n410) );
  XOR2_X1 U389 ( .A(KEYINPUT3), .B(G119), .Z(n473) );
  NOR2_X1 U390 ( .A1(G953), .A2(n703), .ZN(n704) );
  NOR2_X1 U391 ( .A1(n643), .A2(n721), .ZN(n644) );
  AND2_X1 U392 ( .A1(n367), .A2(n366), .ZN(n365) );
  XNOR2_X1 U393 ( .A(n422), .B(KEYINPUT42), .ZN(n749) );
  XOR2_X1 U394 ( .A(KEYINPUT31), .B(n619), .Z(n661) );
  AND2_X1 U395 ( .A1(n405), .A2(n408), .ZN(n403) );
  XNOR2_X1 U396 ( .A(n674), .B(KEYINPUT6), .ZN(n616) );
  XNOR2_X1 U397 ( .A(n516), .B(n395), .ZN(n735) );
  XNOR2_X2 U398 ( .A(n351), .B(G469), .ZN(n579) );
  NOR2_X1 U399 ( .A1(n705), .A2(G902), .ZN(n351) );
  XNOR2_X1 U400 ( .A(n411), .B(n410), .ZN(n602) );
  NAND2_X1 U401 ( .A1(n403), .A2(n402), .ZN(n411) );
  XOR2_X2 U402 ( .A(G110), .B(KEYINPUT75), .Z(n354) );
  XOR2_X1 U403 ( .A(G146), .B(G125), .Z(n516) );
  NAND2_X1 U404 ( .A1(n404), .A2(n375), .ZN(n405) );
  NOR2_X1 U405 ( .A1(n600), .A2(n409), .ZN(n375) );
  OR2_X1 U406 ( .A1(n476), .A2(n461), .ZN(n460) );
  NAND2_X1 U407 ( .A1(n477), .A2(n462), .ZN(n461) );
  INV_X1 U408 ( .A(G902), .ZN(n462) );
  OR2_X1 U409 ( .A1(n353), .A2(n577), .ZN(n391) );
  XNOR2_X1 U410 ( .A(n453), .B(G101), .ZN(n502) );
  INV_X1 U411 ( .A(KEYINPUT68), .ZN(n453) );
  NAND2_X1 U412 ( .A1(n741), .A2(G234), .ZN(n481) );
  XNOR2_X1 U413 ( .A(n588), .B(KEYINPUT38), .ZN(n682) );
  INV_X1 U414 ( .A(KEYINPUT72), .ZN(n373) );
  NAND2_X1 U415 ( .A1(n457), .A2(n464), .ZN(n459) );
  NAND2_X1 U416 ( .A1(n465), .A2(G902), .ZN(n464) );
  NAND2_X1 U417 ( .A1(n476), .A2(n465), .ZN(n457) );
  XNOR2_X1 U418 ( .A(n606), .B(n607), .ZN(n611) );
  AND2_X1 U419 ( .A1(n618), .A2(n466), .ZN(n606) );
  INV_X1 U420 ( .A(KEYINPUT10), .ZN(n395) );
  NOR2_X1 U421 ( .A1(n686), .A2(n685), .ZN(n568) );
  OR2_X1 U422 ( .A1(n508), .A2(n579), .ZN(n569) );
  INV_X1 U423 ( .A(KEYINPUT86), .ZN(n444) );
  NAND2_X1 U424 ( .A1(n627), .A2(n372), .ZN(n371) );
  INV_X1 U425 ( .A(n616), .ZN(n600) );
  INV_X1 U426 ( .A(KEYINPUT33), .ZN(n409) );
  NOR2_X1 U427 ( .A1(G953), .A2(G237), .ZN(n529) );
  INV_X1 U428 ( .A(KEYINPUT48), .ZN(n412) );
  XNOR2_X1 U429 ( .A(n393), .B(KEYINPUT81), .ZN(n392) );
  NAND2_X1 U430 ( .A1(n600), .A2(n409), .ZN(n407) );
  INV_X1 U431 ( .A(KEYINPUT88), .ZN(n523) );
  XNOR2_X1 U432 ( .A(n488), .B(n487), .ZN(n604) );
  XNOR2_X1 U433 ( .A(n486), .B(n485), .ZN(n487) );
  NOR2_X1 U434 ( .A1(n717), .A2(G902), .ZN(n488) );
  XOR2_X1 U435 ( .A(G131), .B(G134), .Z(n468) );
  NAND2_X1 U436 ( .A1(n529), .A2(G210), .ZN(n451) );
  XNOR2_X1 U437 ( .A(KEYINPUT5), .B(KEYINPUT74), .ZN(n450) );
  XNOR2_X1 U438 ( .A(n502), .B(n471), .ZN(n452) );
  XNOR2_X1 U439 ( .A(n513), .B(n512), .ZN(n722) );
  XNOR2_X1 U440 ( .A(n511), .B(G122), .ZN(n512) );
  XOR2_X1 U441 ( .A(KEYINPUT16), .B(KEYINPUT71), .Z(n511) );
  XOR2_X1 U442 ( .A(G137), .B(G140), .Z(n506) );
  XNOR2_X1 U443 ( .A(n480), .B(n479), .ZN(n397) );
  XNOR2_X1 U444 ( .A(KEYINPUT92), .B(KEYINPUT23), .ZN(n479) );
  XNOR2_X1 U445 ( .A(n478), .B(n426), .ZN(n480) );
  XNOR2_X1 U446 ( .A(n433), .B(n432), .ZN(n716) );
  XNOR2_X1 U447 ( .A(n549), .B(n547), .ZN(n432) );
  XNOR2_X1 U448 ( .A(n551), .B(n434), .ZN(n433) );
  XNOR2_X1 U449 ( .A(n538), .B(n379), .ZN(n714) );
  XNOR2_X1 U450 ( .A(n539), .B(n735), .ZN(n379) );
  XNOR2_X1 U451 ( .A(n425), .B(KEYINPUT0), .ZN(n618) );
  NAND2_X1 U452 ( .A1(n463), .A2(n460), .ZN(n674) );
  NOR2_X1 U453 ( .A1(n611), .A2(n608), .ZN(n614) );
  NOR2_X1 U454 ( .A1(n702), .A2(n355), .ZN(n455) );
  XNOR2_X1 U455 ( .A(KEYINPUT85), .B(KEYINPUT46), .ZN(n574) );
  NOR2_X1 U456 ( .A1(G902), .A2(G237), .ZN(n522) );
  NAND2_X1 U457 ( .A1(n370), .A2(n369), .ZN(n368) );
  NOR2_X1 U458 ( .A1(n371), .A2(n444), .ZN(n370) );
  INV_X1 U459 ( .A(KEYINPUT44), .ZN(n442) );
  XNOR2_X1 U460 ( .A(n431), .B(KEYINPUT9), .ZN(n546) );
  INV_X1 U461 ( .A(KEYINPUT7), .ZN(n431) );
  XNOR2_X1 U462 ( .A(G134), .B(G116), .ZN(n543) );
  XOR2_X1 U463 ( .A(G122), .B(G107), .Z(n544) );
  XNOR2_X1 U464 ( .A(G140), .B(KEYINPUT98), .ZN(n534) );
  XOR2_X1 U465 ( .A(G104), .B(G113), .Z(n531) );
  XNOR2_X1 U466 ( .A(G131), .B(G143), .ZN(n532) );
  XOR2_X1 U467 ( .A(G902), .B(KEYINPUT15), .Z(n521) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n489) );
  NOR2_X1 U469 ( .A1(n458), .A2(n459), .ZN(n559) );
  NAND2_X1 U470 ( .A1(n460), .A2(n683), .ZN(n458) );
  NAND2_X1 U471 ( .A1(n604), .A2(n670), .ZN(n667) );
  XNOR2_X1 U472 ( .A(n376), .B(KEYINPUT84), .ZN(n388) );
  INV_X1 U473 ( .A(G146), .ZN(n504) );
  XNOR2_X1 U474 ( .A(n722), .B(n518), .ZN(n519) );
  XNOR2_X1 U475 ( .A(n572), .B(n571), .ZN(n590) );
  INV_X1 U476 ( .A(KEYINPUT39), .ZN(n571) );
  INV_X1 U477 ( .A(n407), .ZN(n406) );
  NOR2_X1 U478 ( .A1(n611), .A2(n671), .ZN(n385) );
  XNOR2_X1 U479 ( .A(n616), .B(n386), .ZN(n609) );
  INV_X1 U480 ( .A(KEYINPUT79), .ZN(n386) );
  INV_X1 U481 ( .A(KEYINPUT32), .ZN(n383) );
  OR2_X2 U482 ( .A1(n588), .A2(n558), .ZN(n445) );
  XNOR2_X1 U483 ( .A(n449), .B(n452), .ZN(n474) );
  XNOR2_X1 U484 ( .A(n451), .B(n450), .ZN(n449) );
  XNOR2_X1 U485 ( .A(n396), .B(n394), .ZN(n717) );
  XNOR2_X1 U486 ( .A(n482), .B(n735), .ZN(n394) );
  XNOR2_X1 U487 ( .A(n398), .B(n397), .ZN(n396) );
  NOR2_X1 U488 ( .A1(n700), .A2(n569), .ZN(n422) );
  INV_X1 U489 ( .A(n610), .ZN(n377) );
  XNOR2_X1 U490 ( .A(n583), .B(KEYINPUT36), .ZN(n378) );
  XNOR2_X1 U491 ( .A(n384), .B(n382), .ZN(n748) );
  XNOR2_X1 U492 ( .A(n423), .B(n383), .ZN(n382) );
  NAND2_X1 U493 ( .A1(n385), .A2(n612), .ZN(n384) );
  INV_X1 U494 ( .A(KEYINPUT78), .ZN(n423) );
  AND2_X1 U495 ( .A1(n424), .A2(n421), .ZN(n651) );
  AND2_X1 U496 ( .A1(n448), .A2(n674), .ZN(n421) );
  XNOR2_X1 U497 ( .A(n381), .B(n380), .ZN(n659) );
  INV_X1 U498 ( .A(KEYINPUT104), .ZN(n380) );
  INV_X1 U499 ( .A(KEYINPUT122), .ZN(n427) );
  INV_X1 U500 ( .A(KEYINPUT60), .ZN(n413) );
  XNOR2_X1 U501 ( .A(n454), .B(KEYINPUT118), .ZN(n703) );
  XNOR2_X1 U502 ( .A(KEYINPUT83), .B(n655), .ZN(n352) );
  AND2_X1 U503 ( .A1(n378), .A2(n377), .ZN(n353) );
  XNOR2_X1 U504 ( .A(n568), .B(KEYINPUT41), .ZN(n700) );
  XOR2_X1 U505 ( .A(n701), .B(KEYINPUT117), .Z(n355) );
  XOR2_X1 U506 ( .A(n524), .B(n523), .Z(n356) );
  AND2_X1 U507 ( .A1(n555), .A2(n554), .ZN(n357) );
  XOR2_X1 U508 ( .A(n526), .B(KEYINPUT89), .Z(n683) );
  BUF_X1 U509 ( .A(n604), .Z(n671) );
  INV_X1 U510 ( .A(n671), .ZN(n448) );
  AND2_X1 U511 ( .A1(n408), .A2(n407), .ZN(n358) );
  XOR2_X1 U512 ( .A(n476), .B(KEYINPUT62), .Z(n359) );
  XOR2_X1 U513 ( .A(n714), .B(n713), .Z(n360) );
  XNOR2_X1 U514 ( .A(n716), .B(KEYINPUT121), .ZN(n361) );
  XOR2_X1 U515 ( .A(n642), .B(n641), .Z(n362) );
  AND2_X1 U516 ( .A1(n444), .A2(KEYINPUT44), .ZN(n363) );
  NOR2_X1 U517 ( .A1(G952), .A2(n741), .ZN(n721) );
  INV_X1 U518 ( .A(n721), .ZN(n417) );
  XNOR2_X2 U519 ( .A(n364), .B(n506), .ZN(n736) );
  XNOR2_X1 U520 ( .A(n475), .B(n364), .ZN(n476) );
  XNOR2_X2 U521 ( .A(n510), .B(n468), .ZN(n364) );
  NAND2_X1 U522 ( .A1(n368), .A2(n365), .ZN(n400) );
  NAND2_X1 U523 ( .A1(n628), .A2(n363), .ZN(n366) );
  NAND2_X1 U524 ( .A1(n371), .A2(n444), .ZN(n367) );
  NAND2_X1 U525 ( .A1(n628), .A2(KEYINPUT44), .ZN(n369) );
  INV_X1 U526 ( .A(n645), .ZN(n372) );
  NAND2_X1 U527 ( .A1(n613), .A2(n748), .ZN(n628) );
  XNOR2_X2 U528 ( .A(n374), .B(n373), .ZN(n617) );
  XNOR2_X2 U529 ( .A(n579), .B(KEYINPUT1), .ZN(n599) );
  NOR2_X1 U530 ( .A1(n621), .A2(n406), .ZN(n402) );
  AND2_X2 U531 ( .A1(n711), .A2(n387), .ZN(n447) );
  NAND2_X1 U532 ( .A1(n443), .A2(n442), .ZN(n441) );
  NAND2_X1 U533 ( .A1(n589), .A2(n435), .ZN(n376) );
  NOR2_X1 U534 ( .A1(n566), .A2(n563), .ZN(n381) );
  NAND2_X1 U535 ( .A1(n447), .A2(G472), .ZN(n419) );
  NAND2_X1 U536 ( .A1(n387), .A2(n698), .ZN(n456) );
  NAND2_X1 U537 ( .A1(n438), .A2(n387), .ZN(n437) );
  NAND2_X1 U538 ( .A1(n712), .A2(n387), .ZN(n715) );
  NAND2_X2 U539 ( .A1(n631), .A2(n630), .ZN(n387) );
  NOR2_X1 U540 ( .A1(n388), .A2(n592), .ZN(n629) );
  XNOR2_X1 U541 ( .A(n388), .B(n740), .ZN(n742) );
  XNOR2_X2 U542 ( .A(n389), .B(n412), .ZN(n589) );
  NAND2_X1 U543 ( .A1(n392), .A2(n390), .ZN(n389) );
  NOR2_X1 U544 ( .A1(n578), .A2(n391), .ZN(n390) );
  NAND2_X1 U545 ( .A1(n357), .A2(n352), .ZN(n393) );
  NAND2_X1 U546 ( .A1(n550), .A2(G221), .ZN(n398) );
  XNOR2_X2 U547 ( .A(n399), .B(KEYINPUT45), .ZN(n729) );
  NAND2_X1 U548 ( .A1(n400), .A2(n441), .ZN(n399) );
  XNOR2_X1 U549 ( .A(n401), .B(n548), .ZN(n434) );
  XNOR2_X2 U550 ( .A(n470), .B(n469), .ZN(n401) );
  NAND2_X1 U551 ( .A1(n617), .A2(n409), .ZN(n408) );
  INV_X1 U552 ( .A(n617), .ZN(n404) );
  NAND2_X1 U553 ( .A1(n358), .A2(n405), .ZN(n699) );
  NAND2_X1 U554 ( .A1(n729), .A2(n638), .ZN(n698) );
  NAND2_X1 U555 ( .A1(n447), .A2(G478), .ZN(n430) );
  AND2_X2 U556 ( .A1(n698), .A2(n521), .ZN(n711) );
  XNOR2_X1 U557 ( .A(n430), .B(n361), .ZN(n429) );
  XNOR2_X1 U558 ( .A(n419), .B(n359), .ZN(n418) );
  NAND2_X1 U559 ( .A1(n429), .A2(n417), .ZN(n428) );
  NAND2_X1 U560 ( .A1(n418), .A2(n417), .ZN(n416) );
  XNOR2_X1 U561 ( .A(n414), .B(n413), .ZN(G60) );
  NAND2_X1 U562 ( .A1(n415), .A2(n417), .ZN(n414) );
  XNOR2_X1 U563 ( .A(n437), .B(n362), .ZN(n643) );
  XNOR2_X1 U564 ( .A(n416), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U565 ( .A(n428), .B(n427), .ZN(G63) );
  XNOR2_X1 U566 ( .A(n715), .B(n360), .ZN(n415) );
  AND2_X2 U567 ( .A1(n711), .A2(G210), .ZN(n438) );
  BUF_X1 U568 ( .A(n588), .Z(n420) );
  XNOR2_X1 U569 ( .A(n439), .B(KEYINPUT76), .ZN(n562) );
  NOR2_X1 U570 ( .A1(n590), .A2(n659), .ZN(n573) );
  OR2_X2 U571 ( .A1(n640), .A2(n521), .ZN(n446) );
  INV_X1 U572 ( .A(n459), .ZN(n463) );
  XNOR2_X1 U573 ( .A(n614), .B(KEYINPUT106), .ZN(n424) );
  NAND2_X1 U574 ( .A1(n589), .A2(n666), .ZN(n637) );
  NOR2_X1 U575 ( .A1(n745), .A2(n436), .ZN(n435) );
  INV_X1 U576 ( .A(n666), .ZN(n436) );
  NAND2_X1 U577 ( .A1(n620), .A2(n557), .ZN(n439) );
  XNOR2_X2 U578 ( .A(n440), .B(n503), .ZN(n509) );
  XNOR2_X1 U579 ( .A(n440), .B(G101), .ZN(n723) );
  XNOR2_X2 U580 ( .A(n354), .B(n501), .ZN(n440) );
  INV_X1 U581 ( .A(n628), .ZN(n443) );
  XNOR2_X2 U582 ( .A(n445), .B(n527), .ZN(n598) );
  XNOR2_X2 U583 ( .A(n446), .B(n356), .ZN(n588) );
  NAND2_X1 U584 ( .A1(n350), .A2(G217), .ZN(n718) );
  NAND2_X1 U585 ( .A1(n350), .A2(G469), .ZN(n708) );
  NOR2_X2 U586 ( .A1(n562), .A2(n561), .ZN(n570) );
  NAND2_X1 U587 ( .A1(n456), .A2(n455), .ZN(n454) );
  INV_X1 U588 ( .A(n477), .ZN(n465) );
  INV_X1 U589 ( .A(n502), .ZN(n503) );
  AND2_X1 U590 ( .A1(n605), .A2(n670), .ZN(n466) );
  AND2_X1 U591 ( .A1(G227), .A2(n741), .ZN(n467) );
  INV_X1 U592 ( .A(G143), .ZN(n469) );
  INV_X1 U593 ( .A(KEYINPUT69), .ZN(n497) );
  XNOR2_X1 U594 ( .A(n474), .B(n513), .ZN(n475) );
  INV_X1 U595 ( .A(n599), .ZN(n608) );
  XNOR2_X2 U596 ( .A(G128), .B(KEYINPUT64), .ZN(n470) );
  XNOR2_X1 U597 ( .A(G146), .B(G137), .ZN(n471) );
  XNOR2_X1 U598 ( .A(G116), .B(G113), .ZN(n472) );
  XNOR2_X1 U599 ( .A(G472), .B(KEYINPUT70), .ZN(n477) );
  XNOR2_X1 U600 ( .A(G128), .B(G119), .ZN(n478) );
  XOR2_X1 U601 ( .A(KEYINPUT8), .B(n481), .Z(n550) );
  XNOR2_X1 U602 ( .A(n506), .B(KEYINPUT24), .ZN(n482) );
  INV_X1 U603 ( .A(n521), .ZN(n639) );
  NAND2_X1 U604 ( .A1(G234), .A2(n639), .ZN(n483) );
  XNOR2_X1 U605 ( .A(KEYINPUT20), .B(n483), .ZN(n494) );
  NAND2_X1 U606 ( .A1(n494), .A2(G217), .ZN(n486) );
  XNOR2_X1 U607 ( .A(KEYINPUT25), .B(KEYINPUT77), .ZN(n484) );
  XOR2_X1 U608 ( .A(n484), .B(KEYINPUT94), .Z(n485) );
  XNOR2_X1 U609 ( .A(n489), .B(KEYINPUT90), .ZN(n490) );
  XNOR2_X1 U610 ( .A(KEYINPUT14), .B(n490), .ZN(n491) );
  NAND2_X1 U611 ( .A1(G952), .A2(n491), .ZN(n697) );
  NOR2_X1 U612 ( .A1(G953), .A2(n697), .ZN(n596) );
  NAND2_X1 U613 ( .A1(n491), .A2(G902), .ZN(n594) );
  OR2_X1 U614 ( .A1(n741), .A2(n594), .ZN(n492) );
  NOR2_X1 U615 ( .A1(G900), .A2(n492), .ZN(n493) );
  NOR2_X1 U616 ( .A1(n596), .A2(n493), .ZN(n556) );
  NOR2_X1 U617 ( .A1(n604), .A2(n556), .ZN(n496) );
  NAND2_X1 U618 ( .A1(n494), .A2(G221), .ZN(n495) );
  XOR2_X1 U619 ( .A(n495), .B(KEYINPUT21), .Z(n670) );
  NAND2_X1 U620 ( .A1(n496), .A2(n670), .ZN(n498) );
  XNOR2_X1 U621 ( .A(n498), .B(n497), .ZN(n580) );
  NOR2_X1 U622 ( .A1(n674), .A2(n580), .ZN(n500) );
  XNOR2_X1 U623 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n499) );
  XNOR2_X1 U624 ( .A(n500), .B(n499), .ZN(n508) );
  XNOR2_X1 U625 ( .A(n736), .B(n507), .ZN(n705) );
  XNOR2_X1 U626 ( .A(n510), .B(n509), .ZN(n520) );
  XOR2_X1 U627 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n515) );
  NAND2_X1 U628 ( .A1(G224), .A2(n741), .ZN(n514) );
  XNOR2_X1 U629 ( .A(n515), .B(n514), .ZN(n517) );
  XNOR2_X1 U630 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U631 ( .A(n519), .B(n520), .ZN(n640) );
  XNOR2_X1 U632 ( .A(n522), .B(KEYINPUT73), .ZN(n525) );
  NAND2_X1 U633 ( .A1(G210), .A2(n525), .ZN(n524) );
  NAND2_X1 U634 ( .A1(n525), .A2(G214), .ZN(n526) );
  INV_X1 U635 ( .A(n683), .ZN(n558) );
  XNOR2_X1 U636 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n527) );
  INV_X1 U637 ( .A(n656), .ZN(n652) );
  NAND2_X1 U638 ( .A1(n652), .A2(KEYINPUT47), .ZN(n528) );
  XNOR2_X1 U639 ( .A(n528), .B(KEYINPUT82), .ZN(n555) );
  XNOR2_X1 U640 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n541) );
  NAND2_X1 U641 ( .A1(G214), .A2(n529), .ZN(n530) );
  XNOR2_X1 U642 ( .A(n531), .B(n530), .ZN(n539) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(G122), .Z(n533) );
  XNOR2_X1 U644 ( .A(n533), .B(n532), .ZN(n537) );
  XOR2_X1 U645 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n535) );
  XNOR2_X1 U646 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U647 ( .A(n537), .B(n536), .Z(n538) );
  NOR2_X1 U648 ( .A1(G902), .A2(n714), .ZN(n540) );
  XNOR2_X1 U649 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U650 ( .A(G475), .B(n542), .ZN(n566) );
  XNOR2_X1 U651 ( .A(n544), .B(n543), .ZN(n549) );
  XOR2_X1 U652 ( .A(KEYINPUT100), .B(KEYINPUT102), .Z(n548) );
  XNOR2_X1 U653 ( .A(KEYINPUT101), .B(KEYINPUT103), .ZN(n545) );
  XNOR2_X1 U654 ( .A(n546), .B(n545), .ZN(n547) );
  NAND2_X1 U655 ( .A1(G217), .A2(n550), .ZN(n551) );
  NOR2_X1 U656 ( .A1(n716), .A2(G902), .ZN(n552) );
  XOR2_X1 U657 ( .A(n552), .B(G478), .Z(n563) );
  NAND2_X1 U658 ( .A1(n566), .A2(n563), .ZN(n662) );
  NAND2_X1 U659 ( .A1(n662), .A2(n659), .ZN(n553) );
  XOR2_X1 U660 ( .A(n553), .B(KEYINPUT105), .Z(n625) );
  INV_X1 U661 ( .A(n625), .ZN(n687) );
  NAND2_X1 U662 ( .A1(n687), .A2(KEYINPUT47), .ZN(n554) );
  INV_X1 U663 ( .A(n556), .ZN(n557) );
  XOR2_X1 U664 ( .A(KEYINPUT108), .B(n559), .Z(n560) );
  XNOR2_X1 U665 ( .A(KEYINPUT30), .B(n560), .ZN(n561) );
  INV_X1 U666 ( .A(n563), .ZN(n567) );
  NOR2_X1 U667 ( .A1(n567), .A2(n566), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n570), .A2(n601), .ZN(n564) );
  NOR2_X1 U669 ( .A1(n420), .A2(n564), .ZN(n655) );
  NAND2_X1 U670 ( .A1(n682), .A2(n683), .ZN(n565) );
  XNOR2_X1 U671 ( .A(n565), .B(KEYINPUT110), .ZN(n686) );
  NAND2_X1 U672 ( .A1(n567), .A2(n566), .ZN(n685) );
  NAND2_X1 U673 ( .A1(n570), .A2(n682), .ZN(n572) );
  XNOR2_X1 U674 ( .A(n575), .B(n574), .ZN(n578) );
  NAND2_X1 U675 ( .A1(n656), .A2(n625), .ZN(n576) );
  NOR2_X1 U676 ( .A1(n576), .A2(KEYINPUT47), .ZN(n577) );
  XOR2_X1 U677 ( .A(KEYINPUT87), .B(n599), .Z(n610) );
  NAND2_X1 U678 ( .A1(n683), .A2(n616), .ZN(n581) );
  NOR2_X1 U679 ( .A1(n581), .A2(n580), .ZN(n582) );
  INV_X1 U680 ( .A(n659), .ZN(n657) );
  NAND2_X1 U681 ( .A1(n582), .A2(n657), .ZN(n584) );
  NOR2_X1 U682 ( .A1(n420), .A2(n584), .ZN(n583) );
  XOR2_X1 U683 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n586) );
  OR2_X1 U684 ( .A1(n584), .A2(n608), .ZN(n585) );
  XNOR2_X1 U685 ( .A(n586), .B(n585), .ZN(n587) );
  NAND2_X1 U686 ( .A1(n420), .A2(n587), .ZN(n666) );
  OR2_X1 U687 ( .A1(n590), .A2(n662), .ZN(n591) );
  XOR2_X1 U688 ( .A(n591), .B(KEYINPUT111), .Z(n632) );
  INV_X1 U689 ( .A(n632), .ZN(n745) );
  NOR2_X1 U690 ( .A1(KEYINPUT80), .A2(n637), .ZN(n592) );
  NOR2_X1 U691 ( .A1(G898), .A2(n741), .ZN(n593) );
  XNOR2_X1 U692 ( .A(KEYINPUT91), .B(n593), .ZN(n725) );
  NOR2_X1 U693 ( .A1(n594), .A2(n725), .ZN(n595) );
  NOR2_X1 U694 ( .A1(n596), .A2(n595), .ZN(n597) );
  INV_X1 U695 ( .A(n618), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U697 ( .A(n603), .B(KEYINPUT35), .ZN(n746) );
  XNOR2_X1 U698 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n607) );
  INV_X1 U699 ( .A(n685), .ZN(n605) );
  NOR2_X1 U700 ( .A1(n746), .A2(n651), .ZN(n613) );
  NOR2_X1 U701 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U702 ( .A1(n671), .A2(n614), .ZN(n615) );
  NOR2_X1 U703 ( .A1(n616), .A2(n615), .ZN(n645) );
  NAND2_X1 U704 ( .A1(n679), .A2(n618), .ZN(n619) );
  NAND2_X1 U705 ( .A1(n674), .A2(n620), .ZN(n622) );
  NOR2_X1 U706 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U707 ( .A(n623), .B(KEYINPUT95), .ZN(n647) );
  XNOR2_X1 U708 ( .A(KEYINPUT96), .B(n624), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n629), .A2(n729), .ZN(n631) );
  INV_X1 U711 ( .A(KEYINPUT2), .ZN(n630) );
  OR2_X1 U712 ( .A1(KEYINPUT80), .A2(n745), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n632), .A2(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n633), .A2(KEYINPUT80), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U717 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n642) );
  XNOR2_X1 U718 ( .A(n640), .B(KEYINPUT55), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n644), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U720 ( .A(G101), .B(n645), .Z(G3) );
  NOR2_X1 U721 ( .A1(n659), .A2(n647), .ZN(n646) );
  XOR2_X1 U722 ( .A(G104), .B(n646), .Z(G6) );
  NOR2_X1 U723 ( .A1(n662), .A2(n647), .ZN(n649) );
  XNOR2_X1 U724 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n648) );
  XNOR2_X1 U725 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U726 ( .A(G107), .B(n650), .ZN(G9) );
  XOR2_X1 U727 ( .A(n651), .B(G110), .Z(G12) );
  XOR2_X1 U728 ( .A(G128), .B(KEYINPUT29), .Z(n654) );
  OR2_X1 U729 ( .A1(n662), .A2(n652), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n654), .B(n653), .ZN(G30) );
  XOR2_X1 U731 ( .A(G143), .B(n655), .Z(G45) );
  NAND2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U733 ( .A(n658), .B(G146), .ZN(G48) );
  NOR2_X1 U734 ( .A1(n659), .A2(n661), .ZN(n660) );
  XOR2_X1 U735 ( .A(G113), .B(n660), .Z(G15) );
  NOR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U737 ( .A(G116), .B(n663), .Z(G18) );
  XNOR2_X1 U738 ( .A(n353), .B(KEYINPUT112), .ZN(n664) );
  XNOR2_X1 U739 ( .A(n664), .B(KEYINPUT37), .ZN(n665) );
  XNOR2_X1 U740 ( .A(G125), .B(n665), .ZN(G27) );
  XNOR2_X1 U741 ( .A(G140), .B(n666), .ZN(G42) );
  XOR2_X1 U742 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n669) );
  NAND2_X1 U743 ( .A1(n599), .A2(n667), .ZN(n668) );
  XNOR2_X1 U744 ( .A(n669), .B(n668), .ZN(n677) );
  OR2_X1 U745 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n672), .B(KEYINPUT49), .ZN(n673) );
  XNOR2_X1 U747 ( .A(KEYINPUT113), .B(n673), .ZN(n675) );
  NAND2_X1 U748 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U751 ( .A(KEYINPUT51), .B(n680), .Z(n681) );
  NOR2_X1 U752 ( .A1(n700), .A2(n681), .ZN(n693) );
  NOR2_X1 U753 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U756 ( .A(KEYINPUT115), .B(n688), .Z(n689) );
  NOR2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U758 ( .A1(n691), .A2(n699), .ZN(n692) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n694), .B(KEYINPUT116), .ZN(n695) );
  XNOR2_X1 U761 ( .A(KEYINPUT52), .B(n695), .ZN(n696) );
  NOR2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n702) );
  NOR2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U764 ( .A(n704), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U765 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n707) );
  XNOR2_X1 U766 ( .A(n705), .B(KEYINPUT120), .ZN(n706) );
  XNOR2_X1 U767 ( .A(n707), .B(n706), .ZN(n709) );
  XNOR2_X1 U768 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n721), .A2(n710), .ZN(G54) );
  AND2_X1 U770 ( .A1(n711), .A2(G475), .ZN(n712) );
  XOR2_X1 U771 ( .A(KEYINPUT59), .B(KEYINPUT66), .Z(n713) );
  XOR2_X1 U772 ( .A(n717), .B(KEYINPUT123), .Z(n719) );
  XNOR2_X1 U773 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U774 ( .A1(n721), .A2(n720), .ZN(G66) );
  XNOR2_X1 U775 ( .A(n722), .B(n723), .ZN(n724) );
  NAND2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n733) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n726) );
  XNOR2_X1 U778 ( .A(KEYINPUT61), .B(n726), .ZN(n727) );
  NAND2_X1 U779 ( .A1(n727), .A2(G898), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n728), .B(KEYINPUT124), .ZN(n731) );
  NAND2_X1 U781 ( .A1(n729), .A2(n741), .ZN(n730) );
  NAND2_X1 U782 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U783 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U784 ( .A(KEYINPUT125), .B(n734), .ZN(G69) );
  XNOR2_X1 U785 ( .A(n736), .B(n735), .ZN(n740) );
  XNOR2_X1 U786 ( .A(G227), .B(n740), .ZN(n737) );
  NAND2_X1 U787 ( .A1(n737), .A2(G900), .ZN(n738) );
  NAND2_X1 U788 ( .A1(G953), .A2(n738), .ZN(n739) );
  XNOR2_X1 U789 ( .A(n739), .B(KEYINPUT126), .ZN(n744) );
  NAND2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n744), .A2(n743), .ZN(G72) );
  XOR2_X1 U792 ( .A(G134), .B(n745), .Z(G36) );
  XNOR2_X1 U793 ( .A(n746), .B(G122), .ZN(n747) );
  XNOR2_X1 U794 ( .A(n747), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U795 ( .A(n748), .B(G119), .ZN(G21) );
  XOR2_X1 U796 ( .A(n749), .B(G137), .Z(G39) );
  XOR2_X1 U797 ( .A(n750), .B(G131), .Z(G33) );
endmodule

