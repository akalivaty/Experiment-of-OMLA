//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT68), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(G137), .A3(new_n463), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n463), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  XNOR2_X1  g048(.A(new_n464), .B(KEYINPUT69), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n463), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n463), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n474), .A2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT70), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n480), .B1(G124), .B2(new_n482), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT71), .Z(G162));
  INV_X1    g059(.A(KEYINPUT74), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n486), .A2(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n464), .A2(new_n487), .A3(new_n463), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n464), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n491), .B(new_n492), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n490), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n463), .B1(new_n494), .B2(new_n495), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n486), .A2(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n488), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n485), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n464), .A2(new_n487), .A3(new_n463), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n508), .B2(new_n488), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(new_n496), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n509), .A2(KEYINPUT74), .A3(new_n490), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT75), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(new_n524), .ZN(new_n528));
  NAND3_X1  g103(.A1(KEYINPUT76), .A2(KEYINPUT5), .A3(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G88), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n526), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n530), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n517), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n535), .A2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND2_X1  g114(.A1(new_n525), .A2(G51), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n533), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G63), .A2(G651), .ZN(new_n543));
  OR3_X1    g118(.A1(new_n531), .A2(KEYINPUT77), .A3(new_n543), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT78), .B(KEYINPUT7), .Z(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n545), .B(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT77), .B1(new_n531), .B2(new_n543), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n542), .A2(new_n549), .ZN(G168));
  AOI22_X1  g125(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n517), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n525), .A2(G52), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n532), .A2(G90), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(G171));
  AOI22_X1  g131(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n517), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n525), .A2(G43), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n532), .A2(G81), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  AOI22_X1  g141(.A1(new_n530), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n517), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n532), .A2(G91), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n521), .A2(G53), .A3(G543), .A4(new_n522), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(KEYINPUT79), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(KEYINPUT79), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(KEYINPUT9), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n571), .A2(KEYINPUT79), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n570), .A2(new_n574), .A3(new_n576), .ZN(G299));
  XNOR2_X1  g152(.A(new_n555), .B(KEYINPUT80), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  NAND2_X1  g154(.A1(new_n532), .A2(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n525), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(G48), .A2(new_n525), .B1(new_n532), .B2(G86), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n530), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n517), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n586), .A2(KEYINPUT81), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n586), .A2(KEYINPUT81), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n532), .A2(G85), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  INV_X1    g166(.A(new_n523), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G543), .ZN(new_n593));
  XOR2_X1   g168(.A(KEYINPUT82), .B(G47), .Z(new_n594));
  OAI221_X1 g169(.A(new_n590), .B1(new_n517), .B2(new_n591), .C1(new_n593), .C2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(new_n532), .A2(G92), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT84), .B(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n531), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n603), .A2(G651), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n525), .A2(G54), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n598), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  MUX2_X1   g182(.A(new_n607), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g183(.A(new_n607), .B(G301), .S(G868), .Z(G321));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g185(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g186(.A(new_n607), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT86), .B(G559), .Z(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(G860), .B2(new_n613), .ZN(G148));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n476), .A2(G135), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT87), .Z(new_n620));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n621));
  NOR3_X1   g196(.A1(new_n621), .A2(new_n463), .A3(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n463), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(G123), .B2(new_n482), .ZN(new_n626));
  INV_X1    g201(.A(G2096), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n464), .A2(new_n470), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2100), .Z(new_n633));
  NAND3_X1  g208(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2443), .B(G2446), .Z(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(G14), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n645), .ZN(G401));
  XNOR2_X1  g226(.A(G2084), .B(G2090), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT90), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  AOI21_X1  g232(.A(KEYINPUT18), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(new_n627), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT20), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n665), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n665), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT91), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G229));
  NOR2_X1   g256(.A1(G16), .A2(G23), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT92), .ZN(new_n683));
  XNOR2_X1  g258(.A(G288), .B(KEYINPUT93), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT33), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n685), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1971), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n685), .A2(G6), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G305), .B2(G16), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT32), .B(G1981), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NOR4_X1   g272(.A1(new_n688), .A2(new_n691), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n482), .A2(G119), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(G107), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G2105), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n476), .B2(G131), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G25), .B2(G29), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  AND2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  MUX2_X1   g288(.A(G24), .B(G290), .S(G16), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1986), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n700), .A2(new_n701), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT36), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n482), .A2(G129), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT26), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n470), .A2(G105), .ZN(new_n722));
  AOI211_X1 g297(.A(new_n721), .B(new_n722), .C1(new_n476), .C2(G141), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n726), .B2(G32), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT27), .B(G1996), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT25), .Z(new_n733));
  AOI22_X1  g308(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  INV_X1    g309(.A(G139), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n733), .B1(new_n463), .B2(new_n734), .C1(new_n475), .C2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT96), .Z(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(new_n726), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n726), .B2(G33), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n730), .B(new_n731), .C1(new_n442), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(G162), .A2(G29), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G29), .B2(G35), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT29), .B(G2090), .Z(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n739), .A2(new_n442), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT97), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n740), .A2(new_n744), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n482), .A2(G128), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G116), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n476), .B2(G140), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT94), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n726), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT95), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT28), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2067), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n626), .A2(G29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n561), .A2(G16), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G16), .B2(G19), .ZN(new_n764));
  INV_X1    g339(.A(G1341), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n685), .A2(G21), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G168), .B2(new_n685), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n764), .A2(new_n765), .B1(new_n767), .B2(G1966), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n762), .B(new_n768), .C1(new_n765), .C2(new_n764), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n685), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n685), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1961), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n767), .A2(G1966), .ZN(new_n773));
  INV_X1    g348(.A(G160), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(G34), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n726), .B1(new_n775), .B2(G34), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n774), .A2(new_n726), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT31), .B(G11), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT98), .ZN(new_n783));
  INV_X1    g358(.A(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT30), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n784), .B2(KEYINPUT30), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n780), .A2(new_n781), .A3(new_n787), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n769), .A2(new_n772), .A3(new_n773), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n612), .A2(new_n685), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G4), .B2(new_n685), .ZN(new_n791));
  INV_X1    g366(.A(G1348), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n685), .A2(G20), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT23), .Z(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G299), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT99), .B(G1956), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n793), .A2(new_n794), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n726), .A2(G27), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G164), .B2(new_n726), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2078), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n798), .B2(new_n797), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n789), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n718), .A2(new_n748), .A3(new_n761), .A4(new_n805), .ZN(G311));
  INV_X1    g381(.A(G311), .ZN(G150));
  AOI22_X1  g382(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(new_n517), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n525), .A2(G55), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n532), .A2(G93), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n561), .B1(KEYINPUT100), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(KEYINPUT100), .B2(new_n812), .ZN(new_n814));
  INV_X1    g389(.A(new_n561), .ZN(new_n815));
  OR3_X1    g390(.A1(new_n815), .A2(KEYINPUT100), .A3(new_n812), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT38), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n612), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n821), .A2(new_n822), .A3(G860), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n812), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n825));
  XOR2_X1   g400(.A(new_n824), .B(new_n825), .Z(new_n826));
  OR2_X1    g401(.A1(new_n823), .A2(new_n826), .ZN(G145));
  NAND2_X1  g402(.A1(new_n482), .A2(G130), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT102), .Z(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n830));
  INV_X1    g405(.A(G118), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(G2105), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n476), .A2(G142), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n829), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n512), .A2(new_n501), .A3(new_n505), .A4(new_n490), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n749), .A2(new_n835), .A3(new_n753), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n835), .B1(new_n749), .B2(new_n753), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n724), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n838), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n840), .A2(new_n725), .A3(new_n836), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n841), .A3(new_n736), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n737), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n839), .B2(new_n841), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n834), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n839), .A2(new_n841), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n737), .ZN(new_n848));
  INV_X1    g423(.A(new_n834), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n849), .A3(new_n842), .ZN(new_n850));
  INV_X1    g425(.A(new_n631), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n846), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n846), .B2(new_n850), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n707), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n846), .A2(new_n850), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n631), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n857), .A2(new_n852), .A3(new_n708), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(G162), .B(new_n774), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(new_n626), .Z(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n855), .A2(new_n858), .A3(new_n859), .A4(new_n862), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g443(.A1(new_n607), .A2(G299), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n607), .A2(G299), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT104), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n817), .B(new_n615), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n869), .A2(KEYINPUT41), .A3(new_n870), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI22_X1  g454(.A1(new_n874), .A2(new_n875), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(new_n875), .B2(new_n874), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n684), .B(G303), .ZN(new_n882));
  XNOR2_X1  g457(.A(G305), .B(G290), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n882), .B(new_n883), .Z(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT42), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n881), .B(new_n885), .ZN(new_n886));
  MUX2_X1   g461(.A(new_n812), .B(new_n886), .S(G868), .Z(G295));
  MUX2_X1   g462(.A(new_n812), .B(new_n886), .S(G868), .Z(G331));
  NOR2_X1   g463(.A1(G301), .A2(G286), .ZN(new_n889));
  NOR2_X1   g464(.A1(G168), .A2(G171), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n817), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n816), .B(new_n814), .C1(new_n889), .C2(new_n890), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n877), .A2(new_n892), .A3(new_n878), .A4(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n893), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n894), .B(new_n895), .C1(new_n897), .C2(new_n871), .ZN(new_n898));
  INV_X1    g473(.A(new_n894), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT106), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n884), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n900), .A3(new_n884), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n865), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n872), .A2(new_n896), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n907), .A2(KEYINPUT107), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(KEYINPUT107), .A3(new_n894), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n884), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(new_n903), .A3(new_n911), .A4(new_n865), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(KEYINPUT44), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n903), .A2(new_n865), .ZN(new_n916));
  INV_X1    g491(.A(new_n910), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(KEYINPUT108), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(KEYINPUT108), .B2(new_n918), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n914), .B1(new_n920), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g496(.A(KEYINPUT126), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n499), .A2(new_n500), .ZN(new_n923));
  AOI22_X1  g498(.A1(new_n489), .A2(new_n923), .B1(new_n511), .B2(new_n496), .ZN(new_n924));
  AOI21_X1  g499(.A(G1384), .B1(new_n924), .B2(new_n509), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n465), .A2(new_n467), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(G2105), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n927), .A2(G40), .A3(new_n471), .A4(new_n469), .ZN(new_n928));
  XNOR2_X1  g503(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n925), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n754), .B(G2067), .Z(new_n932));
  INV_X1    g507(.A(G1996), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n724), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n707), .B(new_n711), .Z(new_n936));
  OAI21_X1  g511(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(G290), .A2(G1986), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G290), .A2(G1986), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(KEYINPUT110), .A3(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n941), .B(new_n931), .C1(KEYINPUT110), .C2(new_n940), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G40), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n468), .A2(new_n472), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n925), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(G8), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1976), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n684), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G288), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(G1976), .ZN(new_n952));
  OR3_X1    g527(.A1(new_n950), .A2(KEYINPUT52), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1981), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n584), .B(new_n954), .C1(new_n587), .C2(new_n588), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n584), .A2(new_n586), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n955), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n947), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n958), .B2(new_n957), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n950), .B2(KEYINPUT52), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n950), .A2(new_n961), .A3(KEYINPUT52), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n953), .B(new_n960), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(G303), .A2(G8), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT55), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n835), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n945), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n514), .A2(new_n969), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(new_n929), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT111), .B(G1971), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n507), .B2(new_n513), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G2090), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n928), .B1(new_n970), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n976), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n968), .B1(new_n985), .B2(G8), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n945), .B1(new_n970), .B2(new_n982), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n980), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n988), .B1(new_n976), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n968), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n965), .A2(new_n987), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT62), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n514), .A2(new_n969), .A3(new_n930), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT45), .B1(new_n835), .B2(new_n969), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n999), .B2(new_n928), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT114), .B(new_n945), .C1(new_n925), .C2(KEYINPUT45), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1966), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n928), .B1(new_n925), .B2(new_n981), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(KEYINPUT115), .A3(new_n779), .A4(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1006), .B(new_n779), .C1(new_n977), .C2(new_n978), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1004), .A2(new_n1007), .A3(new_n1010), .A4(G168), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1004), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(G286), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n996), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1011), .A2(G8), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(KEYINPUT51), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n995), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1014), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT51), .B1(new_n1019), .B2(new_n1016), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1012), .A2(new_n996), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(KEYINPUT62), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n994), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n974), .B2(new_n443), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n990), .A2(G1961), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n997), .A2(new_n1000), .A3(new_n443), .A4(new_n1001), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1026), .A2(KEYINPUT121), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT53), .B1(new_n1026), .B2(KEYINPUT121), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT122), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n928), .B1(new_n970), .B2(new_n971), .ZN(new_n1032));
  AOI22_X1  g607(.A1(KEYINPUT114), .A2(new_n1032), .B1(new_n977), .B2(new_n930), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n443), .A4(new_n1000), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1026), .A2(KEYINPUT121), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(KEYINPUT53), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(KEYINPUT122), .A3(new_n1025), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1024), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT123), .B1(new_n1039), .B2(G301), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1024), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1037), .A2(KEYINPUT122), .A3(new_n1025), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT122), .B1(new_n1037), .B2(new_n1025), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n1045));
  INV_X1    g620(.A(G301), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1040), .A2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1023), .A2(new_n1048), .A3(KEYINPUT124), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT124), .B1(new_n1023), .B2(new_n1048), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n964), .A2(new_n993), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n960), .A2(new_n949), .A3(new_n951), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n947), .B1(new_n1052), .B2(new_n955), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT116), .B(KEYINPUT63), .Z(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n993), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1057), .A2(new_n964), .A3(new_n986), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1013), .A2(G8), .A3(G168), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1056), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT63), .B1(new_n992), .B2(new_n968), .ZN(new_n1062));
  NOR4_X1   g637(.A1(new_n1057), .A2(new_n1062), .A3(new_n964), .A4(new_n1059), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1054), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1049), .A2(new_n1050), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n994), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT53), .B(new_n443), .C1(new_n925), .C2(new_n930), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1041), .B(new_n1025), .C1(new_n972), .C2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G171), .ZN(new_n1069));
  OAI211_X1 g644(.A(KEYINPUT54), .B(new_n1069), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n1072));
  NOR2_X1   g647(.A1(new_n1068), .A2(new_n1046), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n1048), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n946), .A2(G2067), .ZN(new_n1075));
  XOR2_X1   g650(.A(new_n1075), .B(KEYINPUT117), .Z(new_n1076));
  OR2_X1    g651(.A1(new_n990), .A2(G1348), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(new_n612), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n607), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT60), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n607), .A2(KEYINPUT60), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n974), .A2(new_n933), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n974), .A2(KEYINPUT118), .A3(new_n933), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT58), .B(G1341), .Z(new_n1088));
  NAND2_X1  g663(.A1(new_n946), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1090), .A2(new_n1091), .A3(new_n561), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1090), .B2(new_n561), .ZN(new_n1093));
  INV_X1    g668(.A(new_n574), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n568), .A2(new_n569), .A3(new_n576), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT57), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n570), .A2(new_n574), .A3(new_n1097), .A4(new_n576), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1101), .B(new_n972), .C1(new_n929), .C2(new_n973), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1956), .B1(new_n979), .B2(new_n983), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1099), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1103), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n974), .A2(new_n1100), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1099), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1092), .A2(new_n1093), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1090), .A2(new_n561), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT59), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1090), .A2(new_n1091), .A3(new_n561), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1112), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1110), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(KEYINPUT119), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1083), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1080), .A2(new_n1108), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1124), .A2(new_n1104), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1071), .B(new_n1074), .C1(new_n1123), .C2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n943), .B1(new_n1065), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n932), .A2(new_n725), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n931), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n931), .A2(new_n933), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT46), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT47), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n708), .A2(new_n711), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n935), .A2(new_n1135), .B1(G2067), .B2(new_n754), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n938), .A2(new_n931), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT48), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n931), .A2(new_n1136), .B1(new_n937), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT125), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n922), .B1(new_n1128), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n943), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1070), .B(new_n1066), .C1(new_n1123), .C2(new_n1126), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1072), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1040), .A2(new_n1047), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1073), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1023), .A2(new_n1048), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1064), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1023), .A2(new_n1048), .A3(KEYINPUT124), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1143), .B1(new_n1149), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1141), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(KEYINPUT126), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1142), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g734(.A1(new_n461), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1161));
  AOI21_X1  g735(.A(new_n1161), .B1(new_n906), .B2(new_n912), .ZN(new_n1162));
  AND3_X1   g736(.A1(new_n867), .A2(KEYINPUT127), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g737(.A(KEYINPUT127), .B1(new_n867), .B2(new_n1162), .ZN(new_n1164));
  NOR2_X1   g738(.A1(new_n1163), .A2(new_n1164), .ZN(G308));
  NAND2_X1  g739(.A1(new_n867), .A2(new_n1162), .ZN(G225));
endmodule


