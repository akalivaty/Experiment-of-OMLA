//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT81), .ZN(new_n204));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT75), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n209), .B(new_n205), .C1(new_n212), .C2(KEYINPUT75), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT29), .ZN(new_n217));
  AND2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G141gat), .B(G148gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(G155gat), .B2(G162gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G141gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G141gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G155gat), .B(G162gat), .ZN(new_n230));
  INV_X1    g029(.A(G155gat), .ZN(new_n231));
  INV_X1    g030(.A(G162gat), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT2), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n224), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n216), .B1(new_n217), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n224), .A2(new_n234), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n213), .A2(new_n209), .A3(new_n205), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n210), .A2(new_n212), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(new_n217), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n238), .B1(new_n241), .B2(new_n235), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n204), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n224), .A2(new_n234), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT29), .B1(new_n214), .B2(new_n215), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g045(.A(new_n216), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n236), .A2(new_n217), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n203), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n246), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G22gat), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n243), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n243), .B2(new_n251), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT82), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G78gat), .B(G106gat), .Z(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT31), .ZN(new_n257));
  INV_X1    g056(.A(G50gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n243), .A2(new_n251), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(new_n252), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n255), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT83), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT83), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n255), .A2(new_n262), .A3(new_n265), .A4(new_n259), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n253), .A2(new_n254), .ZN(new_n268));
  INV_X1    g067(.A(new_n259), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G227gat), .ZN(new_n273));
  INV_X1    g072(.A(G233gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276));
  AND2_X1   g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n276), .B1(new_n277), .B2(KEYINPUT24), .ZN(new_n278));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT24), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT64), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(KEYINPUT64), .A3(new_n280), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n278), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT66), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(G169gat), .A3(G176gat), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n286), .A2(new_n288), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT65), .B(G176gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n286), .A2(G169gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G176gat), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n281), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n290), .A2(new_n292), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n286), .ZN(new_n306));
  AND4_X1   g105(.A1(new_n301), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n291), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n289), .A2(KEYINPUT66), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n314));
  NOR3_X1   g113(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT68), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n305), .A2(new_n317), .A3(new_n310), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G190gat), .ZN(new_n320));
  AND2_X1   g119(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g124(.A(KEYINPUT28), .B(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n277), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n319), .A2(KEYINPUT69), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT69), .B1(new_n319), .B2(new_n327), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n309), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G113gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT70), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT70), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G113gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n334), .A3(G120gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(G113gat), .B2(G120gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(G127gat), .A2(G134gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(G127gat), .A2(G134gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(G113gat), .A2(G120gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n339), .B(new_n340), .C1(new_n337), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT69), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n305), .A2(new_n317), .A3(new_n310), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n317), .B1(new_n305), .B2(new_n310), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT26), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n287), .A2(KEYINPUT68), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT68), .B1(new_n287), .B2(new_n351), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT27), .B(G183gat), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT28), .B1(new_n356), .B2(new_n320), .ZN(new_n357));
  INV_X1    g156(.A(new_n326), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n279), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n348), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n319), .A2(KEYINPUT69), .A3(new_n327), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n345), .A3(new_n309), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n275), .B1(new_n347), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT72), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n366));
  NOR3_X1   g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n275), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n345), .B1(new_n362), .B2(new_n309), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n307), .B1(new_n297), .B2(new_n298), .ZN(new_n370));
  AOI211_X1 g169(.A(new_n346), .B(new_n370), .C1(new_n360), .C2(new_n361), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n366), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT72), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n347), .A2(new_n275), .A3(new_n363), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377));
  XNOR2_X1  g176(.A(G15gat), .B(G43gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(G71gat), .ZN(new_n379));
  INV_X1    g178(.A(G99gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n376), .B(KEYINPUT32), .C1(new_n377), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n376), .A2(KEYINPUT32), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n376), .A2(new_n377), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n381), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT34), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n364), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n375), .A2(new_n383), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n383), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n365), .B1(new_n364), .B2(new_n366), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n372), .A2(KEYINPUT72), .A3(new_n373), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n388), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(KEYINPUT73), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n390), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n272), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n342), .A2(new_n224), .A3(new_n234), .A4(new_n344), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT78), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT4), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n400), .B2(KEYINPUT4), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n408), .A2(new_n345), .A3(new_n236), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n399), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n405), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n400), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n412), .B(new_n413), .C1(new_n414), .C2(new_n400), .ZN(new_n415));
  OR3_X1    g214(.A1(new_n415), .A2(new_n399), .A3(new_n409), .ZN(new_n416));
  INV_X1    g215(.A(new_n413), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n345), .A2(new_n244), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n400), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n419), .B2(new_n399), .ZN(new_n420));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT0), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(G57gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G85gat), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n410), .A2(new_n416), .A3(new_n420), .A4(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n425), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT79), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n400), .A2(KEYINPUT4), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT78), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n346), .A2(new_n238), .A3(new_n411), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n402), .ZN(new_n433));
  INV_X1    g232(.A(new_n409), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT5), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n415), .A2(new_n399), .A3(new_n409), .ZN(new_n436));
  INV_X1    g235(.A(new_n420), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n429), .B1(new_n438), .B2(new_n424), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n410), .A2(new_n416), .A3(new_n420), .ZN(new_n440));
  INV_X1    g239(.A(new_n424), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(KEYINPUT79), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n442), .A3(new_n426), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n428), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n439), .A2(new_n442), .A3(KEYINPUT80), .A4(new_n426), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n427), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G226gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(new_n274), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(KEYINPUT29), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n349), .A2(new_n350), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n359), .B1(new_n451), .B2(new_n316), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n452), .B2(new_n370), .ZN(new_n453));
  INV_X1    g252(.A(new_n449), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n453), .B(new_n216), .C1(new_n330), .C2(new_n454), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n452), .A2(new_n370), .A3(new_n454), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n456), .B1(new_n330), .B2(new_n450), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n457), .B2(new_n216), .ZN(new_n458));
  XNOR2_X1  g257(.A(G8gat), .B(G36gat), .ZN(new_n459));
  INV_X1    g258(.A(G64gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(G92gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(KEYINPUT30), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n458), .B2(new_n462), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT76), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT76), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n463), .B(new_n466), .C1(new_n458), .C2(new_n462), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT30), .B1(new_n458), .B2(new_n462), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n447), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n202), .B1(new_n398), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n427), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n438), .A2(KEYINPUT85), .A3(new_n424), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n425), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n473), .B1(new_n477), .B2(new_n443), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n464), .A2(new_n468), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT88), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n390), .A2(new_n393), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n390), .A2(new_n393), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n271), .A2(new_n202), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT88), .B1(new_n478), .B2(new_n479), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n469), .B(new_n463), .C1(new_n458), .C2(new_n462), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n413), .B1(new_n433), .B2(new_n434), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n419), .A2(new_n417), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n489), .A2(new_n490), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n492), .A2(new_n493), .A3(new_n424), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n494), .A2(KEYINPUT40), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n476), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(KEYINPUT40), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n488), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n496), .A2(new_n426), .A3(new_n442), .A4(new_n439), .ZN(new_n499));
  XOR2_X1   g298(.A(KEYINPUT87), .B(KEYINPUT38), .Z(new_n500));
  OAI21_X1  g299(.A(KEYINPUT86), .B1(new_n457), .B2(new_n247), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n453), .B(new_n247), .C1(new_n330), .C2(new_n454), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503));
  INV_X1    g302(.A(new_n450), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n362), .B2(new_n309), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n503), .B(new_n216), .C1(new_n505), .C2(new_n456), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT37), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n462), .B1(new_n458), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n500), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n455), .B(KEYINPUT37), .C1(new_n457), .C2(new_n216), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n510), .A2(new_n500), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n473), .B(new_n499), .C1(new_n511), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n458), .A2(new_n462), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n271), .B(new_n498), .C1(new_n514), .C2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT84), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n267), .A2(new_n518), .A3(new_n270), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n267), .B2(new_n270), .ZN(new_n520));
  OAI22_X1  g319(.A1(new_n447), .A2(new_n470), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n395), .B2(new_n397), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(new_n389), .B2(new_n394), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  OAI22_X1  g327(.A1(new_n472), .A2(new_n487), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G43gat), .B(G50gat), .Z(new_n530));
  INV_X1    g329(.A(KEYINPUT89), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G43gat), .B(G50gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT89), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(KEYINPUT15), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT15), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT90), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n537), .B2(new_n538), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n536), .A2(new_n530), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n535), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(G29gat), .A2(G36gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT14), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(new_n539), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n544), .A2(new_n546), .B1(new_n547), .B2(new_n535), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT17), .ZN(new_n549));
  INV_X1    g348(.A(G8gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(G15gat), .B(G22gat), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n551), .A2(G1gat), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n552), .B2(KEYINPUT91), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT16), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n551), .B1(new_n554), .B2(G1gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n556), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n549), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n548), .ZN(new_n562));
  NAND2_X1  g361(.A1(G229gat), .A2(G233gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT18), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n559), .B(new_n548), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n563), .B(KEYINPUT13), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n571), .A2(new_n573), .B1(new_n565), .B2(new_n566), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(G197gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT11), .ZN(new_n578));
  INV_X1    g377(.A(G169gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT12), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n570), .A2(new_n583), .A3(new_n574), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n529), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT7), .B1(new_n587), .B2(KEYINPUT94), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(KEYINPUT94), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G106gat), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n380), .A2(new_n591), .A3(KEYINPUT95), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT95), .B1(new_n380), .B2(new_n591), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(KEYINPUT8), .A3(new_n593), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n590), .B(new_n594), .C1(G85gat), .C2(G92gat), .ZN(new_n595));
  XOR2_X1   g394(.A(G99gat), .B(G106gat), .Z(new_n596));
  OR2_X1    g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(KEYINPUT96), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT96), .B1(new_n597), .B2(new_n598), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n549), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n598), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n548), .A3(new_n599), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G190gat), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n602), .A2(new_n607), .A3(new_n320), .A4(new_n603), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n208), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n609), .A2(G218gat), .A3(new_n610), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(KEYINPUT93), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT97), .ZN(new_n616));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n612), .A2(KEYINPUT93), .A3(new_n613), .A4(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G57gat), .B(G64gat), .Z(new_n623));
  INV_X1    g422(.A(G71gat), .ZN(new_n624));
  INV_X1    g423(.A(G78gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n623), .B1(KEYINPUT9), .B2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G71gat), .B(G78gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G127gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n629), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n559), .B1(KEYINPUT21), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n632), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n636));
  XNOR2_X1  g435(.A(G155gat), .B(G183gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n635), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n207), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n639), .B(new_n641), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n622), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(G230gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n274), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n597), .A2(new_n629), .A3(new_n598), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n629), .B1(new_n597), .B2(new_n598), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n633), .A4(new_n599), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n645), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n649), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(new_n645), .A3(new_n647), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n300), .ZN(new_n658));
  INV_X1    g457(.A(G204gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n656), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n643), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n586), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n447), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT98), .B(G1gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1324gat));
  XNOR2_X1  g467(.A(KEYINPUT16), .B(G8gat), .ZN(new_n669));
  NOR2_X1   g468(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n664), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n488), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n671), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n673), .B(KEYINPUT99), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(G8gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(G1325gat));
  INV_X1    g478(.A(G15gat), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n395), .A2(new_n397), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT36), .ZN(new_n683));
  INV_X1    g482(.A(new_n527), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n524), .A2(KEYINPUT101), .A3(new_n527), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n664), .A2(new_n680), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n483), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n680), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n519), .A2(new_n520), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n664), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  INV_X1    g494(.A(new_n622), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n642), .A2(new_n662), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT102), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n698), .A2(KEYINPUT102), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n586), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(G29gat), .A3(new_n665), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT45), .Z(new_n703));
  AND3_X1   g502(.A1(new_n529), .A2(KEYINPUT44), .A3(new_n696), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n683), .A2(new_n681), .A3(new_n684), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT101), .B1(new_n524), .B2(new_n527), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n522), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n472), .A2(new_n487), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n696), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n704), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n582), .A2(KEYINPUT103), .A3(new_n584), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n583), .B1(new_n570), .B2(new_n574), .ZN(new_n714));
  INV_X1    g513(.A(new_n574), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n581), .B(new_n715), .C1(new_n568), .C2(new_n569), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n711), .A2(new_n697), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n665), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n720), .ZN(G1328gat));
  NOR3_X1   g520(.A1(new_n701), .A2(G36gat), .A3(new_n479), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  OAI21_X1  g522(.A(G36gat), .B1(new_n719), .B2(new_n479), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1329gat));
  NAND2_X1  g524(.A1(new_n687), .A2(G43gat), .ZN(new_n726));
  INV_X1    g525(.A(new_n483), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n701), .A2(new_n727), .ZN(new_n728));
  OAI22_X1  g527(.A1(new_n719), .A2(new_n726), .B1(G43gat), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g529(.A(G50gat), .B1(new_n719), .B2(new_n271), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n701), .B(KEYINPUT104), .ZN(new_n732));
  INV_X1    g531(.A(new_n692), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n258), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT105), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n731), .B(KEYINPUT48), .C1(new_n732), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n732), .A2(new_n735), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n719), .A2(new_n692), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(G50gat), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(new_n739), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g539(.A1(new_n517), .A2(new_n521), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n685), .B2(new_n686), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n398), .A2(new_n471), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT35), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n643), .A2(new_n718), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n748), .A3(new_n662), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n747), .A2(new_n748), .A3(new_n751), .A4(new_n662), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n447), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT107), .B(G57gat), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1332gat));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n488), .B1(new_n757), .B2(new_n460), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT108), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n760), .A2(KEYINPUT109), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(KEYINPUT109), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n757), .A2(new_n460), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n761), .A2(new_n757), .A3(new_n460), .A4(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1333gat));
  XNOR2_X1  g566(.A(new_n483), .B(KEYINPUT111), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n624), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n750), .A2(G71gat), .A3(new_n687), .A4(new_n752), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(KEYINPUT110), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(KEYINPUT110), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT50), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n770), .B(new_n776), .C1(new_n772), .C2(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1334gat));
  NAND2_X1  g577(.A1(new_n753), .A2(new_n733), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g579(.A1(new_n529), .A2(KEYINPUT44), .A3(new_n696), .ZN(new_n781));
  INV_X1    g580(.A(new_n662), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n718), .A2(new_n642), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n622), .B1(new_n742), .B2(new_n746), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n781), .B(new_n783), .C1(new_n784), .C2(KEYINPUT44), .ZN(new_n785));
  OAI21_X1  g584(.A(G85gat), .B1(new_n785), .B2(new_n665), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n718), .A2(new_n642), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n696), .B(new_n787), .C1(new_n708), .C2(new_n709), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT112), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n784), .A2(KEYINPUT51), .A3(new_n787), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n788), .A2(new_n793), .A3(new_n789), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n796), .A2(G85gat), .A3(new_n665), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n786), .B1(new_n797), .B2(new_n782), .ZN(G1336gat));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  NOR2_X1   g599(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n788), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n801), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n747), .A2(new_n696), .A3(new_n787), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n782), .A2(G92gat), .A3(new_n479), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT114), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809));
  AOI211_X1 g608(.A(new_n809), .B(new_n806), .C1(new_n802), .C2(new_n804), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G92gat), .B1(new_n785), .B2(new_n479), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n800), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(new_n795), .B2(new_n807), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n711), .A2(new_n815), .A3(new_n488), .A4(new_n783), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT115), .B1(new_n785), .B2(new_n479), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(G92gat), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n799), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n788), .B(new_n803), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n809), .B1(new_n821), .B2(new_n806), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n805), .A2(KEYINPUT114), .A3(new_n807), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n812), .A3(new_n823), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n824), .A2(KEYINPUT52), .B1(new_n814), .B2(new_n818), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT116), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n820), .A2(new_n826), .ZN(G1337gat));
  OAI21_X1  g626(.A(G99gat), .B1(new_n785), .B2(new_n688), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n795), .A2(new_n380), .A3(new_n483), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(new_n782), .ZN(G1338gat));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831));
  OAI21_X1  g630(.A(G106gat), .B1(new_n785), .B2(new_n271), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n272), .A2(new_n662), .A3(new_n591), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n831), .B(new_n832), .C1(new_n796), .C2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G106gat), .B1(new_n785), .B2(new_n692), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n821), .B2(new_n833), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT53), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(G1339gat));
  NOR2_X1   g637(.A1(new_n665), .A2(new_n488), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n642), .ZN(new_n841));
  INV_X1    g640(.A(new_n652), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n650), .A2(new_n651), .A3(new_n645), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(KEYINPUT54), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n661), .B1(new_n652), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(KEYINPUT55), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n656), .A2(new_n661), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT55), .B1(new_n844), .B2(new_n846), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n712), .A3(new_n717), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n563), .B1(new_n561), .B2(new_n562), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n571), .A2(new_n573), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n580), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n662), .A2(new_n584), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n696), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n584), .A2(new_n855), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n851), .A2(new_n620), .A3(new_n621), .A4(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n841), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n712), .A2(new_n717), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(new_n642), .A3(new_n622), .A4(new_n782), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n840), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n692), .A3(new_n483), .ZN(new_n866));
  INV_X1    g665(.A(new_n585), .ZN(new_n867));
  OAI21_X1  g666(.A(G113gat), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n398), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n863), .B1(new_n332), .B2(new_n334), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT117), .ZN(G1340gat));
  OR3_X1    g673(.A1(new_n869), .A2(G120gat), .A3(new_n782), .ZN(new_n875));
  OAI21_X1  g674(.A(G120gat), .B1(new_n866), .B2(new_n782), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1341gat));
  NOR2_X1   g676(.A1(new_n866), .A2(new_n841), .ZN(new_n878));
  INV_X1    g677(.A(G127gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n870), .A2(new_n881), .A3(new_n642), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT118), .B1(new_n869), .B2(new_n841), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n880), .B1(new_n884), .B2(new_n879), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n885), .B(new_n886), .ZN(G1342gat));
  NOR3_X1   g686(.A1(new_n869), .A2(G134gat), .A3(new_n622), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT56), .ZN(new_n889));
  OAI21_X1  g688(.A(G134gat), .B1(new_n866), .B2(new_n622), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1343gat));
  NOR2_X1   g690(.A1(new_n687), .A2(new_n840), .ZN(new_n892));
  XNOR2_X1  g691(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n652), .A2(new_n845), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n660), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n652), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n714), .B2(new_n716), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n856), .B1(new_n899), .B2(new_n849), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n622), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n642), .B1(new_n901), .B2(new_n860), .ZN(new_n902));
  INV_X1    g701(.A(new_n864), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT57), .B(new_n733), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n622), .A2(new_n858), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n907), .A2(new_n851), .B1(new_n900), .B2(new_n622), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n864), .B1(new_n908), .B2(new_n642), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n909), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n733), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n271), .B1(new_n862), .B2(new_n864), .ZN(new_n912));
  XNOR2_X1  g711(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n892), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G141gat), .B1(new_n915), .B2(new_n867), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  INV_X1    g716(.A(new_n912), .ZN(new_n918));
  INV_X1    g717(.A(new_n892), .ZN(new_n919));
  NOR4_X1   g718(.A1(new_n918), .A2(G141gat), .A3(new_n867), .A4(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n916), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n718), .B(new_n892), .C1(new_n911), .C2(new_n914), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G141gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n921), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n923), .B1(new_n926), .B2(KEYINPUT58), .ZN(new_n927));
  AOI211_X1 g726(.A(KEYINPUT123), .B(new_n917), .C1(new_n925), .C2(new_n921), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(G1344gat));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n913), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n643), .A2(new_n585), .A3(new_n662), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n733), .B1(new_n902), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n782), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n227), .B1(new_n935), .B2(new_n892), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(KEYINPUT125), .A3(KEYINPUT59), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT59), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n940), .B(G148gat), .C1(new_n915), .C2(new_n782), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n918), .A2(new_n919), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n227), .A3(new_n662), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT124), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n946), .ZN(G1345gat));
  NOR3_X1   g746(.A1(new_n915), .A2(new_n231), .A3(new_n841), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n918), .A2(new_n841), .A3(new_n919), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n949), .A2(KEYINPUT126), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(KEYINPUT126), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n952), .B2(new_n231), .ZN(G1346gat));
  OAI21_X1  g752(.A(G162gat), .B1(new_n915), .B2(new_n622), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n944), .A2(new_n232), .A3(new_n696), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1347gat));
  NOR2_X1   g755(.A1(new_n447), .A2(new_n479), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n958), .B1(new_n862), .B2(new_n864), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(new_n398), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n579), .A3(new_n718), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n692), .A3(new_n768), .ZN(new_n962));
  OAI21_X1  g761(.A(G169gat), .B1(new_n962), .B2(new_n867), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1348gat));
  AOI21_X1  g763(.A(G176gat), .B1(new_n960), .B2(new_n662), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n962), .A2(new_n294), .A3(new_n782), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(G1349gat));
  NAND3_X1  g766(.A1(new_n960), .A2(new_n356), .A3(new_n642), .ZN(new_n968));
  OAI21_X1  g767(.A(G183gat), .B1(new_n962), .B2(new_n841), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g770(.A1(KEYINPUT127), .A2(KEYINPUT61), .ZN(new_n972));
  OAI211_X1 g771(.A(G190gat), .B(new_n972), .C1(new_n962), .C2(new_n622), .ZN(new_n973));
  NOR2_X1   g772(.A1(KEYINPUT127), .A2(KEYINPUT61), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n320), .A3(new_n696), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n974), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(G1351gat));
  NOR2_X1   g777(.A1(new_n687), .A2(new_n958), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n918), .A2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(G197gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n981), .A2(new_n982), .A3(new_n718), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n980), .B1(new_n930), .B2(new_n934), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n984), .A2(new_n585), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n983), .B1(new_n985), .B2(new_n982), .ZN(G1352gat));
  NAND3_X1  g785(.A1(new_n981), .A2(new_n659), .A3(new_n662), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n659), .B1(new_n935), .B2(new_n979), .ZN(new_n990));
  OR3_X1    g789(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(G1353gat));
  NAND3_X1  g790(.A1(new_n981), .A2(new_n207), .A3(new_n642), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n984), .A2(new_n642), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n993), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n994));
  AOI21_X1  g793(.A(KEYINPUT63), .B1(new_n993), .B2(G211gat), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(G1354gat));
  AOI21_X1  g795(.A(G218gat), .B1(new_n981), .B2(new_n696), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n622), .A2(new_n208), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n997), .B1(new_n984), .B2(new_n998), .ZN(G1355gat));
endmodule


