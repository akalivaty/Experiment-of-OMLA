//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n203), .B1(new_n204), .B2(G13), .ZN(new_n205));
  INV_X1    g0005(.A(G13), .ZN(new_n206));
  NAND4_X1  g0006(.A1(new_n206), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT66), .Z(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G116), .ZN(new_n215));
  INV_X1    g0015(.A(G270), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G68), .B2(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT65), .B(G244), .Z(new_n224));
  AOI211_X1 g0024(.A(new_n212), .B(new_n223), .C1(G77), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(G1), .B2(G20), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G58), .ZN(new_n231));
  INV_X1    g0031(.A(G68), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n210), .B(new_n227), .C1(new_n230), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n216), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n229), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n219), .A2(new_n231), .A3(new_n232), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n254), .A2(G150), .B1(new_n255), .B2(G20), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n231), .A2(KEYINPUT8), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  MUX2_X1   g0058(.A(new_n257), .B(new_n258), .S(KEYINPUT69), .Z(new_n259));
  NAND2_X1  g0059(.A1(new_n229), .A2(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n228), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n262), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G20), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n261), .A2(new_n267), .B1(new_n269), .B2(G50), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n219), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT9), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n252), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G222), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G223), .A2(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G77), .B2(new_n280), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  OAI211_X1 g0087(.A(G1), .B(G13), .C1(new_n252), .C2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n284), .B(new_n290), .C1(G77), .C2(new_n280), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n286), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n288), .A2(new_n293), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(G226), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G200), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n270), .A2(KEYINPUT9), .A3(new_n273), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n292), .A2(G190), .A3(new_n297), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n276), .A2(new_n299), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n300), .A2(new_n301), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(new_n276), .A4(new_n299), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n232), .A2(G20), .ZN(new_n308));
  INV_X1    g0108(.A(G77), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n308), .B1(new_n260), .B2(new_n309), .C1(new_n219), .C2(new_n253), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n267), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n311), .B(KEYINPUT72), .Z(new_n312));
  OR2_X1    g0112(.A1(new_n312), .A2(KEYINPUT11), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n308), .A2(G1), .A3(new_n206), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(KEYINPUT12), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n314), .A2(KEYINPUT12), .ZN(new_n316));
  AOI211_X1 g0116(.A(new_n315), .B(new_n316), .C1(new_n269), .C2(G68), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(KEYINPUT11), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n313), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT71), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n280), .A2(G226), .A3(new_n281), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n280), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n322), .A2(new_n323), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n295), .B1(new_n326), .B2(new_n289), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n296), .A2(G238), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n328), .B1(new_n327), .B2(new_n329), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n319), .B1(G190), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(G200), .B1(new_n330), .B2(new_n331), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n298), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n292), .A2(new_n338), .A3(new_n297), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n274), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n258), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n254), .B1(G20), .B2(G77), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT15), .B(G87), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n260), .B2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n267), .B1(new_n269), .B2(G77), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n272), .A2(new_n309), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT70), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n281), .A2(G232), .ZN(new_n350));
  INV_X1    g0150(.A(G238), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n280), .B(new_n350), .C1(new_n351), .C2(new_n281), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(new_n289), .C1(G107), .C2(new_n280), .ZN(new_n353));
  INV_X1    g0153(.A(new_n295), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n296), .A2(new_n224), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G200), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n345), .A2(KEYINPUT70), .A3(new_n346), .ZN(new_n358));
  INV_X1    g0158(.A(G190), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n349), .A2(new_n357), .A3(new_n358), .A4(new_n360), .ZN(new_n361));
  AND4_X1   g0161(.A1(new_n307), .A2(new_n335), .A3(new_n340), .A4(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(G169), .B1(new_n330), .B2(new_n331), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT14), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n332), .A2(G179), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n366), .B(G169), .C1(new_n330), .C2(new_n331), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n319), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n356), .A2(new_n336), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n347), .B(new_n370), .C1(G179), .C2(new_n356), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  OR2_X1    g0173(.A1(G223), .A2(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n220), .A2(G1698), .ZN(new_n375));
  AND2_X1   g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NOR2_X1   g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n374), .B(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT73), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(new_n382), .A3(new_n379), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n289), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n288), .A2(G232), .A3(new_n293), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT74), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n288), .A2(new_n387), .A3(G232), .A4(new_n293), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n295), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n384), .A2(G179), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n336), .B1(new_n384), .B2(new_n389), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT75), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n378), .A2(new_n382), .A3(new_n379), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n382), .B1(new_n378), .B2(new_n379), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n393), .A2(new_n394), .A3(new_n288), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n386), .A2(new_n388), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n354), .ZN(new_n397));
  OAI21_X1  g0197(.A(G169), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT75), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n384), .A2(G179), .A3(new_n389), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n278), .A2(new_n229), .A3(new_n279), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n279), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G68), .ZN(new_n408));
  INV_X1    g0208(.A(G159), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n253), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G58), .A2(G68), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n229), .B1(new_n233), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n413), .B1(new_n407), .B2(G68), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(KEYINPUT16), .A3(new_n411), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n267), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n259), .A2(new_n272), .ZN(new_n421));
  INV_X1    g0221(.A(new_n267), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(G1), .B2(new_n229), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n423), .B2(new_n259), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n402), .A2(KEYINPUT18), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT18), .B1(new_n402), .B2(new_n426), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n384), .A2(G190), .A3(new_n389), .ZN(new_n430));
  OAI21_X1  g0230(.A(G200), .B1(new_n395), .B2(new_n397), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n420), .A2(new_n430), .A3(new_n431), .A4(new_n425), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n433), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n362), .A2(new_n373), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n271), .A2(new_n215), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n268), .A2(G33), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n265), .A2(new_n266), .A3(new_n271), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n443), .B2(new_n215), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n262), .A2(new_n228), .B1(G20), .B2(new_n215), .ZN(new_n445));
  NAND2_X1  g0245(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G283), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(new_n229), .C1(G33), .C2(new_n221), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n445), .B2(new_n448), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n449), .A2(new_n450), .B1(KEYINPUT83), .B2(KEYINPUT20), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n268), .A2(G45), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT78), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT5), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G41), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT78), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n457), .A2(new_n458), .A3(new_n268), .A4(G45), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n294), .B1(KEYINPUT5), .B2(new_n287), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n455), .A2(new_n459), .A3(new_n288), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n268), .A3(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n456), .A2(G41), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n288), .B(G270), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n461), .A2(new_n464), .A3(KEYINPUT82), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G264), .A2(G1698), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n280), .B(new_n470), .C1(new_n222), .C2(G1698), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(new_n289), .C1(G303), .C2(new_n280), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n452), .A2(new_n469), .A3(G179), .A4(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n461), .A2(KEYINPUT82), .A3(new_n464), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT82), .B1(new_n461), .B2(new_n464), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G200), .ZN(new_n477));
  INV_X1    g0277(.A(new_n452), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n477), .B(new_n478), .C1(new_n359), .C2(new_n476), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT21), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n336), .B1(new_n469), .B2(new_n472), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n452), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n476), .A2(new_n452), .A3(new_n480), .A4(G169), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n473), .B(new_n479), .C1(new_n482), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT84), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n476), .A2(new_n452), .A3(G169), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT21), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n483), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT84), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n473), .A4(new_n479), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT81), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n271), .A2(G97), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n443), .B2(G97), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT76), .B1(new_n407), .B2(G107), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT76), .ZN(new_n497));
  INV_X1    g0297(.A(G107), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n497), .B(new_n498), .C1(new_n405), .C2(new_n406), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n500), .A2(new_n221), .A3(G107), .ZN(new_n501));
  XNOR2_X1  g0301(.A(G97), .B(G107), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n503), .A2(new_n229), .B1(new_n309), .B2(new_n253), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n496), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n495), .B1(new_n505), .B2(new_n422), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n288), .B(G257), .C1(new_n462), .C2(new_n463), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(G244), .B(new_n281), .C1(new_n376), .C2(new_n377), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT77), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n510), .A2(KEYINPUT4), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n280), .A2(G244), .A3(new_n281), .A4(new_n511), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n447), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n508), .B1(new_n516), .B2(new_n289), .ZN(new_n517));
  AOI21_X1  g0317(.A(G169), .B1(new_n517), .B2(new_n461), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n338), .A3(new_n461), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n506), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n495), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n407), .A2(G107), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n497), .ZN(new_n524));
  INV_X1    g0324(.A(new_n504), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n407), .A2(KEYINPUT76), .A3(G107), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n522), .B1(new_n527), .B2(new_n267), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n517), .A2(new_n461), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G200), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n517), .A2(G190), .A3(new_n461), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n521), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n351), .A2(new_n281), .ZN(new_n534));
  INV_X1    g0334(.A(G244), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G1698), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n534), .B(new_n536), .C1(new_n376), .C2(new_n377), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n289), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n454), .A2(new_n214), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n268), .A2(new_n294), .A3(G45), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n288), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT79), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n288), .B1(new_n537), .B2(new_n538), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT79), .B1(new_n547), .B2(new_n543), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G190), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT80), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n213), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n323), .A2(new_n229), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(KEYINPUT19), .A3(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n229), .B(G68), .C1(new_n376), .C2(new_n377), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n323), .A2(G20), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n556), .B(new_n557), .C1(KEYINPUT19), .C2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(new_n267), .B1(new_n272), .B2(new_n343), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n443), .A2(G87), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n545), .B1(new_n540), .B2(new_n544), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n547), .A2(new_n543), .A3(KEYINPUT79), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n562), .B1(new_n565), .B2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n549), .A2(KEYINPUT80), .A3(G190), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n552), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n338), .B1(new_n563), .B2(new_n564), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n560), .B1(new_n343), .B2(new_n442), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n570), .C1(G169), .C2(new_n549), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n493), .B1(new_n533), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n288), .B(G264), .C1(new_n462), .C2(new_n463), .ZN(new_n574));
  INV_X1    g0374(.A(G294), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n252), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n278), .A2(new_n279), .B1(new_n222), .B2(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n214), .A2(new_n281), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n461), .B(new_n574), .C1(new_n579), .C2(new_n288), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(G179), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n336), .B2(new_n580), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT23), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n229), .B2(G107), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n498), .A2(KEYINPUT23), .A3(G20), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n229), .B(G87), .C1(new_n376), .C2(new_n377), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT85), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT22), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n589), .A2(KEYINPUT22), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n588), .A2(new_n593), .A3(new_n590), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(KEYINPUT24), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  INV_X1    g0396(.A(new_n594), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(new_n591), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n267), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n443), .A2(G107), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n272), .B(new_n498), .C1(KEYINPUT86), .C2(KEYINPUT25), .ZN(new_n601));
  NAND2_X1  g0401(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n582), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n222), .A2(G1698), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n578), .B(new_n606), .C1(new_n376), .C2(new_n377), .ZN(new_n607));
  INV_X1    g0407(.A(new_n576), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n289), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(new_n359), .A3(new_n461), .A4(new_n574), .ZN(new_n611));
  INV_X1    g0411(.A(G200), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n611), .A2(KEYINPUT87), .B1(new_n580), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n580), .A2(KEYINPUT87), .A3(new_n612), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n605), .B1(new_n604), .B2(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n521), .A2(new_n568), .A3(new_n532), .A4(new_n571), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n617), .B2(KEYINPUT81), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n439), .A2(new_n492), .A3(new_n573), .A4(new_n618), .ZN(G372));
  OAI211_X1 g0419(.A(new_n473), .B(new_n605), .C1(new_n482), .C2(new_n484), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n527), .A2(new_n267), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n518), .B1(new_n621), .B2(new_n495), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n516), .A2(new_n289), .ZN(new_n623));
  AND4_X1   g0423(.A1(G190), .A2(new_n623), .A3(new_n461), .A4(new_n507), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n612), .B1(new_n517), .B2(new_n461), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n622), .A2(new_n520), .B1(new_n626), .B2(new_n528), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n615), .A2(new_n604), .ZN(new_n628));
  OAI21_X1  g0428(.A(G200), .B1(new_n547), .B2(new_n543), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n560), .A2(new_n561), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n550), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n547), .A2(new_n543), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n336), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n569), .A2(new_n570), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n628), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n620), .A2(new_n627), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT26), .B1(new_n572), .B2(new_n521), .ZN(new_n639));
  INV_X1    g0439(.A(new_n635), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n506), .A2(new_n631), .A3(new_n519), .A4(new_n520), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n439), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n432), .B(KEYINPUT17), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n372), .A2(new_n646), .A3(new_n335), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n398), .A2(new_n400), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n426), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT18), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT18), .B1(new_n426), .B2(new_n648), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n307), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n645), .A2(new_n340), .A3(new_n655), .ZN(G369));
  NAND3_X1  g0456(.A1(new_n268), .A2(new_n229), .A3(G13), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n486), .A2(new_n491), .B1(new_n452), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n489), .A2(new_n473), .ZN(new_n664));
  INV_X1    g0464(.A(new_n662), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n664), .A2(new_n478), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n604), .A2(new_n662), .ZN(new_n670));
  OAI22_X1  g0470(.A1(new_n616), .A2(new_n670), .B1(new_n605), .B2(new_n665), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OR3_X1    g0472(.A1(new_n664), .A2(new_n616), .A3(new_n662), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n662), .B(KEYINPUT88), .Z(new_n674));
  NAND3_X1  g0474(.A1(new_n582), .A2(new_n604), .A3(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0478(.A(new_n208), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n553), .A2(new_n213), .A3(new_n215), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n680), .A2(new_n268), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n235), .B2(new_n680), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT28), .Z(new_n684));
  INV_X1    g0484(.A(new_n521), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n685), .A2(new_n642), .A3(new_n571), .A4(new_n568), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n686), .B(new_n635), .C1(new_n642), .C2(new_n641), .ZN(new_n687));
  INV_X1    g0487(.A(new_n638), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n665), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT94), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT29), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n618), .A2(new_n492), .A3(new_n573), .A4(new_n674), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n549), .A2(G179), .A3(new_n517), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n476), .A2(new_n580), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT30), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(KEYINPUT30), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n695), .A2(new_n696), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n580), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n469), .A2(new_n472), .A3(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n697), .B(KEYINPUT30), .C1(new_n703), .C2(new_n694), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n633), .A2(KEYINPUT90), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT90), .ZN(new_n707));
  AOI21_X1  g0507(.A(G179), .B1(new_n632), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n476), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT91), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT91), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n476), .A2(new_n706), .A3(new_n711), .A4(new_n708), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n710), .A2(new_n529), .A3(new_n580), .A4(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n705), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n712), .A2(new_n529), .A3(new_n580), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT93), .B1(new_n716), .B2(new_n710), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n662), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n705), .A2(new_n713), .ZN(new_n721));
  INV_X1    g0521(.A(new_n674), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n693), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n644), .A2(new_n674), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT94), .B1(new_n726), .B2(new_n691), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n691), .B2(new_n689), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n692), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n684), .B1(new_n730), .B2(G1), .ZN(G364));
  AOI21_X1  g0531(.A(new_n228), .B1(G20), .B2(new_n336), .ZN(new_n732));
  INV_X1    g0532(.A(new_n280), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n229), .A2(new_n359), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n338), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G322), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n359), .A2(G179), .A3(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n229), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n338), .A2(new_n612), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G326), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n740), .A2(new_n575), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT98), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(KEYINPUT98), .ZN(new_n746));
  INV_X1    g0546(.A(G311), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n229), .A2(G190), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n735), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n745), .B(new_n746), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT99), .Z(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(new_n338), .A3(new_n612), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT96), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n738), .B(new_n751), .C1(G329), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n741), .A2(new_n748), .ZN(new_n759));
  INV_X1    g0559(.A(G317), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(KEYINPUT33), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(KEYINPUT33), .B2(new_n760), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n612), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n748), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n758), .B(new_n762), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n734), .A2(new_n764), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n766), .B1(G303), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n740), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n771), .B1(new_n231), .B2(new_n736), .C1(new_n219), .C2(new_n742), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n765), .A2(new_n498), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n759), .A2(new_n232), .ZN(new_n774));
  NOR4_X1   g0574(.A1(new_n772), .A2(new_n733), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n757), .A2(KEYINPUT32), .A3(G159), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT32), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n756), .B2(new_n409), .ZN(new_n778));
  INV_X1    g0578(.A(new_n749), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n776), .A2(new_n778), .B1(G77), .B2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n775), .B(new_n780), .C1(new_n213), .C2(new_n767), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT97), .Z(new_n782));
  OAI21_X1  g0582(.A(new_n732), .B1(new_n769), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n206), .A2(G20), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n268), .B1(new_n784), .B2(G45), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n680), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n667), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n679), .A2(new_n733), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G355), .ZN(new_n793));
  INV_X1    g0593(.A(G45), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n247), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n679), .A2(new_n280), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G45), .B2(new_n234), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n793), .B1(G116), .B2(new_n208), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n790), .A2(new_n732), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT95), .Z(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n783), .A2(new_n787), .A3(new_n791), .A4(new_n801), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n663), .A2(new_n666), .A3(G330), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n669), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n787), .B2(new_n804), .ZN(G396));
  NOR2_X1   g0605(.A1(new_n371), .A2(new_n662), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n347), .A2(new_n662), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n361), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n806), .B1(new_n808), .B2(new_n371), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n726), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n644), .A2(new_n674), .A3(new_n809), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n725), .B(new_n813), .Z(new_n814));
  INV_X1    g0614(.A(new_n787), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n732), .ZN(new_n817));
  INV_X1    g0617(.A(new_n736), .ZN(new_n818));
  INV_X1    g0618(.A(new_n759), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G143), .A2(new_n818), .B1(new_n819), .B2(G150), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n821), .B2(new_n742), .C1(new_n409), .C2(new_n749), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT34), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n823), .A2(KEYINPUT34), .B1(G58), .B2(new_n770), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n733), .B1(new_n757), .B2(G132), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n767), .A2(new_n219), .B1(new_n765), .B2(new_n232), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT100), .Z(new_n828));
  NAND4_X1  g0628(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n771), .B1(new_n498), .B2(new_n767), .C1(new_n756), .C2(new_n747), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G283), .B2(new_n819), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n765), .A2(new_n213), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n742), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G303), .A2(new_n834), .B1(new_n818), .B2(G294), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n280), .B1(new_n779), .B2(G116), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n831), .A2(new_n833), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n817), .B1(new_n829), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n732), .A2(new_n788), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n815), .B(new_n838), .C1(new_n309), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n789), .B2(new_n809), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n816), .A2(new_n841), .ZN(G384));
  AOI21_X1  g0642(.A(new_n438), .B1(new_n728), .B2(new_n692), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n655), .A2(new_n340), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT39), .ZN(new_n846));
  INV_X1    g0646(.A(new_n660), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT16), .B1(new_n418), .B2(new_n411), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n232), .B1(new_n405), .B2(new_n406), .ZN(new_n849));
  NOR4_X1   g0649(.A1(new_n849), .A2(new_n416), .A3(new_n410), .A4(new_n413), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n848), .A2(new_n850), .A3(new_n422), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n847), .B1(new_n851), .B2(new_n424), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT75), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n399), .B1(new_n398), .B2(new_n400), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n426), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n650), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n402), .A2(KEYINPUT18), .A3(new_n426), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n852), .B1(new_n858), .B2(new_n646), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n649), .A2(new_n432), .A3(new_n852), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n852), .A2(new_n432), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT37), .B1(new_n402), .B2(new_n426), .ZN(new_n863));
  AOI22_X1  g0663(.A1(KEYINPUT37), .A2(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n859), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n434), .B(new_n435), .C1(new_n651), .C2(new_n652), .ZN(new_n866));
  INV_X1    g0666(.A(new_n852), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n862), .A2(new_n863), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT38), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n846), .B1(new_n865), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n368), .A2(new_n319), .A3(new_n665), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n860), .B1(new_n859), .B2(new_n864), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n867), .B1(new_n429), .B2(new_n436), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n871), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT39), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n873), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n876), .A2(new_n878), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n319), .A2(new_n882), .A3(new_n662), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n319), .A2(new_n662), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n369), .A2(new_n335), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n368), .A2(new_n319), .A3(new_n662), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT103), .ZN(new_n889));
  INV_X1    g0689(.A(new_n806), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n812), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n889), .B1(new_n812), .B2(new_n890), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n881), .B(new_n888), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n653), .A2(new_n847), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n880), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n845), .B(new_n895), .ZN(new_n896));
  XOR2_X1   g0696(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n897));
  OAI211_X1 g0697(.A(KEYINPUT31), .B(new_n662), .C1(new_n715), .C2(new_n717), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n693), .A2(new_n720), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n810), .B1(new_n886), .B2(new_n887), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n877), .B2(new_n871), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n865), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n897), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n864), .B1(new_n867), .B2(new_n866), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n878), .B1(new_n905), .B2(KEYINPUT38), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n906), .A2(KEYINPUT40), .A3(new_n899), .A4(new_n900), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n904), .A2(new_n439), .A3(new_n899), .A4(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n904), .A2(G330), .A3(new_n907), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n899), .A2(G330), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n438), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n908), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n896), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n268), .B2(new_n784), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT35), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n503), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G116), .A3(new_n230), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT101), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n916), .B2(new_n503), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT36), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n235), .A2(G77), .A3(new_n412), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT102), .Z(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(G50), .B2(new_n232), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n206), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n915), .A2(new_n921), .A3(new_n925), .ZN(G367));
  INV_X1    g0726(.A(G150), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n280), .B1(new_n736), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n765), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(G77), .ZN(new_n930));
  INV_X1    g0730(.A(G143), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(new_n931), .B2(new_n742), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(G58), .B2(new_n768), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n759), .A2(new_n409), .B1(new_n749), .B2(new_n219), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT107), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(new_n232), .C2(new_n740), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n928), .B(new_n936), .C1(G137), .C2(new_n757), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT108), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n767), .A2(new_n215), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT46), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n742), .A2(new_n747), .B1(new_n749), .B2(new_n763), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n733), .B1(new_n765), .B2(new_n221), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(G303), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n736), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n940), .B(new_n945), .C1(G107), .C2(new_n770), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n575), .B2(new_n759), .C1(new_n760), .C2(new_n756), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n938), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n732), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n562), .A2(new_n662), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n640), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT106), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n953), .B(new_n954), .C1(new_n636), .C2(new_n952), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n953), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n790), .ZN(new_n957));
  INV_X1    g0757(.A(new_n796), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n799), .B1(new_n208), .B2(new_n343), .C1(new_n243), .C2(new_n958), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n950), .A2(new_n787), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n627), .B1(new_n528), .B2(new_n674), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n685), .A2(new_n722), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n676), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT44), .B1(new_n676), .B2(new_n963), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n676), .A2(KEYINPUT44), .A3(new_n963), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n966), .A2(new_n672), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n964), .A2(new_n965), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT45), .B1(new_n676), .B2(new_n963), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n967), .B(new_n968), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n672), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n671), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n664), .B2(new_n662), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(new_n673), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n669), .B(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n729), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n969), .A2(new_n974), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n730), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n680), .B(KEYINPUT41), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n786), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n963), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n984), .A2(new_n673), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n521), .B1(new_n961), .B2(new_n605), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n674), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT43), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n956), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n956), .A2(new_n990), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n992), .A2(new_n994), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n996), .A2(new_n997), .B1(new_n672), .B2(new_n984), .ZN(new_n998));
  INV_X1    g0798(.A(new_n997), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n672), .A2(new_n984), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n1000), .A3(new_n995), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n960), .B1(new_n983), .B2(new_n1002), .ZN(G387));
  NOR2_X1   g0803(.A1(new_n259), .A2(new_n759), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G68), .A2(new_n779), .B1(new_n929), .B2(G97), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n219), .B2(new_n736), .C1(new_n409), .C2(new_n742), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(G150), .C2(new_n757), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n768), .A2(G77), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n740), .A2(new_n343), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1007), .A2(new_n280), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G311), .A2(new_n819), .B1(new_n818), .B2(G317), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n944), .B2(new_n749), .C1(new_n737), .C2(new_n742), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT48), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n763), .B2(new_n740), .C1(new_n575), .C2(new_n767), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT49), .Z(new_n1015));
  OAI221_X1 g0815(.A(new_n733), .B1(new_n215), .B2(new_n765), .C1(new_n756), .C2(new_n743), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1010), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n815), .B1(new_n1017), .B2(new_n732), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n958), .B1(new_n240), .B2(G45), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n681), .B2(new_n792), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n341), .A2(new_n219), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n794), .B1(new_n232), .B2(new_n309), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1022), .A2(new_n681), .A3(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1020), .A2(new_n1024), .B1(G107), .B2(new_n208), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n800), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n790), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1018), .B(new_n1026), .C1(new_n671), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n978), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n680), .B1(new_n730), .B2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1028), .B1(new_n785), .B2(new_n978), .C1(new_n1030), .C2(new_n979), .ZN(G393));
  OAI221_X1 g0831(.A(new_n799), .B1(new_n221), .B2(new_n208), .C1(new_n958), .C2(new_n250), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n833), .B1(new_n258), .B2(new_n749), .C1(new_n309), .C2(new_n740), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n280), .B1(new_n767), .B2(new_n232), .C1(new_n219), .C2(new_n759), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n742), .A2(new_n927), .B1(new_n736), .B2(new_n409), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1036), .B(new_n1037), .Z(new_n1038));
  OAI211_X1 g0838(.A(new_n1035), .B(new_n1038), .C1(new_n931), .C2(new_n756), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n742), .A2(new_n760), .B1(new_n736), .B2(new_n747), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT52), .Z(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G116), .B2(new_n770), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n779), .A2(G294), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n757), .A2(G322), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n280), .B(new_n773), .C1(G283), .C2(new_n768), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n759), .A2(new_n944), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1039), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n815), .B1(new_n1048), .B2(new_n732), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1032), .B(new_n1049), .C1(new_n963), .C2(new_n1027), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n969), .A2(new_n974), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1050), .B1(new_n1051), .B2(new_n785), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n680), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n979), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1052), .B1(new_n980), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(G390));
  OAI21_X1  g0857(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1058), .A2(new_n874), .B1(new_n873), .B2(new_n879), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n808), .A2(new_n371), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n665), .B(new_n1060), .C1(new_n687), .C2(new_n688), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1061), .A2(new_n890), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n888), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n906), .B(new_n874), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n724), .A2(new_n888), .A3(G330), .A4(new_n809), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1059), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n899), .A2(G330), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n900), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n873), .A2(new_n879), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n812), .A2(new_n890), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT103), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n812), .A2(new_n889), .A3(new_n890), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1063), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1071), .B1(new_n1075), .B2(new_n875), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1070), .B1(new_n1076), .B2(new_n1064), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1068), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n786), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT113), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT113), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1078), .A2(new_n1081), .A3(new_n786), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1071), .A2(new_n788), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n259), .A2(new_n839), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n740), .A2(new_n309), .B1(new_n736), .B2(new_n215), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT115), .Z(new_n1087));
  NAND2_X1  g0887(.A1(new_n757), .A2(G294), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n834), .A2(G283), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n213), .A2(new_n767), .B1(new_n759), .B2(new_n498), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n232), .A2(new_n765), .B1(new_n749), .B2(new_n221), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1090), .A2(new_n1091), .A3(new_n280), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n768), .A2(G150), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  INV_X1    g0895(.A(G125), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n756), .A2(new_n1096), .B1(new_n409), .B2(new_n740), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n280), .B1(new_n765), .B2(new_n219), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT114), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n819), .A2(G137), .ZN(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT54), .B(G143), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1100), .B1(new_n1101), .B2(new_n742), .C1(new_n749), .C2(new_n1102), .ZN(new_n1103));
  OR4_X1    g0903(.A1(new_n1095), .A2(new_n1097), .A3(new_n1099), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(G132), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n736), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1093), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n815), .B1(new_n1107), .B2(new_n732), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1084), .A2(new_n1085), .A3(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1083), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT112), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1070), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1076), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n843), .A2(new_n844), .A3(new_n912), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n899), .A2(G330), .A3(new_n809), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1063), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n724), .A2(G330), .A3(new_n809), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1069), .A2(new_n900), .B1(new_n1119), .B2(new_n1063), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n891), .A2(new_n892), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n680), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(KEYINPUT110), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT110), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1123), .A2(new_n1126), .A3(new_n680), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1122), .A2(new_n1115), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT111), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1068), .B2(new_n1077), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1113), .A2(new_n1114), .A3(KEYINPUT111), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1111), .B1(new_n1128), .B2(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1123), .A2(new_n1126), .A3(new_n680), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1126), .B1(new_n1123), .B2(new_n680), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1111), .B(new_n1134), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1110), .B1(new_n1135), .B2(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1115), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1078), .B2(new_n1129), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT119), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n895), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT55), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n307), .A2(new_n1148), .A3(new_n340), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n307), .B2(new_n340), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n274), .A2(new_n847), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n274), .B(new_n847), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1147), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1147), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n909), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n909), .A2(new_n1158), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1146), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n909), .A2(new_n1158), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1157), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1163), .A2(new_n1155), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1164), .A2(new_n904), .A3(G330), .A4(new_n907), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1162), .A2(new_n1165), .A3(new_n1145), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1141), .B1(new_n1143), .B2(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n880), .A2(new_n893), .A3(new_n894), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1162), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1123), .A2(new_n1115), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(KEYINPUT57), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1168), .A2(new_n1174), .A3(new_n680), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1167), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n786), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1164), .A2(new_n788), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n219), .B1(new_n376), .B2(G41), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n740), .A2(new_n927), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n1101), .A2(new_n736), .B1(new_n767), .B2(new_n1102), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT117), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n1096), .B2(new_n742), .C1(new_n821), .C2(new_n749), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1180), .B(new_n1183), .C1(G132), .C2(new_n819), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT59), .ZN(new_n1185));
  AOI21_X1  g0985(.A(G33), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(G41), .B1(new_n757), .B2(G124), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n409), .C2(new_n765), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1179), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n834), .A2(G116), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n929), .A2(G58), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1191), .A2(new_n1008), .A3(new_n1192), .A4(new_n733), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n759), .A2(new_n221), .B1(new_n749), .B2(new_n343), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT116), .Z(new_n1195));
  AOI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(G107), .C2(new_n818), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G41), .B1(new_n770), .B2(G68), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n763), .C2(new_n756), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT58), .Z(new_n1199));
  OAI21_X1  g0999(.A(new_n732), .B1(new_n1190), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n815), .B1(new_n219), .B2(new_n839), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1178), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1175), .A2(new_n1177), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT120), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1175), .A2(new_n1177), .A3(new_n1203), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT120), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1208), .ZN(G375));
  NAND2_X1  g1009(.A1(new_n1063), .A2(new_n788), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1192), .B1(new_n759), .B2(new_n1102), .C1(new_n756), .C2(new_n1101), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n740), .A2(new_n219), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n742), .A2(new_n1105), .B1(new_n736), .B2(new_n821), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1211), .A2(new_n733), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n927), .B2(new_n749), .C1(new_n409), .C2(new_n767), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n930), .B1(new_n221), .B2(new_n767), .C1(new_n215), .C2(new_n759), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n280), .B(new_n1216), .C1(G303), .C2(new_n757), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1009), .B1(new_n763), .B2(new_n736), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT121), .Z(new_n1219));
  NAND2_X1  g1019(.A1(new_n779), .A2(G107), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n834), .A2(G294), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1217), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n817), .B1(new_n1215), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n815), .B(new_n1223), .C1(new_n232), .C2(new_n839), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1122), .A2(new_n786), .B1(new_n1210), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1122), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1142), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n982), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1225), .B1(new_n1228), .B2(new_n1129), .ZN(G381));
  NAND2_X1  g1029(.A1(new_n1083), .A2(new_n1109), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1134), .B2(new_n1128), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(G375), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1056), .B(new_n960), .C1(new_n983), .C2(new_n1002), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1234), .A2(G396), .A3(G393), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(G381), .A2(G384), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT122), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1237), .A2(KEYINPUT122), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1233), .A2(new_n1238), .A3(new_n1239), .ZN(G407));
  INV_X1    g1040(.A(G213), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1233), .B2(new_n661), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(G407), .ZN(G409));
  XOR2_X1   g1043(.A(G393), .B(G396), .Z(new_n1244));
  NAND2_X1  g1044(.A1(G387), .A2(G390), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1234), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(KEYINPUT125), .A3(new_n1234), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1244), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1244), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1176), .A2(new_n982), .A3(new_n1173), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1202), .B1(new_n1172), .B2(new_n786), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1110), .A2(new_n1254), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1254), .A2(KEYINPUT112), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1230), .B1(new_n1259), .B2(new_n1138), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1260), .B2(new_n1206), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1241), .A2(G343), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1053), .B1(new_n1227), .B2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1265), .B(new_n1130), .C1(new_n1264), .C2(new_n1227), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(G384), .A3(new_n1225), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(G384), .B1(new_n1266), .B2(new_n1225), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1261), .A2(new_n1263), .A3(new_n1270), .ZN(new_n1271));
  OR2_X1    g1071(.A1(new_n1271), .A2(KEYINPUT62), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(KEYINPUT62), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G378), .A2(new_n1204), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1262), .B1(new_n1276), .B2(new_n1258), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1262), .A2(G2897), .ZN(new_n1278));
  XOR2_X1   g1078(.A(new_n1278), .B(KEYINPUT123), .Z(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1269), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1267), .A3(new_n1279), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1277), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1253), .B1(new_n1275), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT124), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n1277), .B2(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1289), .A2(KEYINPUT124), .A3(new_n1283), .A4(new_n1281), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1273), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1271), .A2(KEYINPUT63), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1261), .A2(new_n1294), .A3(new_n1270), .A4(new_n1263), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1292), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1291), .A2(new_n1296), .A3(KEYINPUT126), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT126), .B1(new_n1291), .B2(new_n1296), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1286), .B1(new_n1297), .B2(new_n1298), .ZN(G405));
  NAND2_X1  g1099(.A1(G375), .A2(new_n1231), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1270), .B1(new_n1300), .B2(new_n1276), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1232), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1276), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1270), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1302), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT127), .B1(new_n1301), .B2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1300), .A2(new_n1276), .A3(new_n1270), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT127), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1304), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1306), .A2(new_n1253), .A3(new_n1310), .ZN(new_n1311));
  OAI221_X1 g1111(.A(KEYINPUT127), .B1(new_n1250), .B2(new_n1252), .C1(new_n1301), .C2(new_n1305), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(G402));
endmodule


