//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n219), .B1(new_n201), .B2(new_n220), .C1(new_n205), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n212), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n212), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n210), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n230), .A2(G50), .A3(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n224), .B(new_n227), .C1(new_n229), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G222), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n256), .B1(new_n257), .B2(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n250), .C2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G274), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n268), .B1(G226), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(G200), .B2(new_n273), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n228), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT66), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n210), .B2(G1), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n209), .A2(KEYINPUT66), .A3(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n280), .A2(G50), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G58), .A2(G68), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n210), .B1(new_n286), .B2(new_n214), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n210), .A2(new_n250), .ZN(new_n288));
  INV_X1    g0088(.A(G150), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g0090(.A(KEYINPUT8), .B(G58), .Z(new_n291));
  NOR2_X1   g0091(.A1(new_n250), .A2(G20), .ZN(new_n292));
  AOI211_X1 g0092(.A(new_n287), .B(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n278), .A2(new_n228), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n285), .B1(G50), .B2(new_n277), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n296), .A2(new_n297), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(KEYINPUT67), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n276), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(KEYINPUT67), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(KEYINPUT67), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n276), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n273), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n296), .C1(G179), .C2(new_n273), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n304), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n277), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n202), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT12), .ZN(new_n314));
  NOR2_X1   g0114(.A1(G20), .A2(G33), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n316));
  INV_X1    g0116(.A(new_n292), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n257), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(KEYINPUT11), .A3(new_n294), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n280), .A2(G68), .A3(new_n284), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n314), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT11), .B1(new_n318), .B2(new_n294), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT14), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT13), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n264), .A2(G238), .A3(new_n269), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n267), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT68), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n267), .A2(new_n327), .A3(KEYINPUT68), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n251), .A2(new_n253), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n333), .A2(new_n215), .A3(G1698), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n251), .A2(new_n253), .A3(G232), .A4(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n261), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n326), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n267), .A2(new_n327), .A3(KEYINPUT68), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT68), .B1(new_n267), .B2(new_n327), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n338), .B(new_n326), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n325), .B(G169), .C1(new_n339), .C2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT13), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(G179), .A3(new_n342), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n342), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n325), .B1(new_n349), .B2(G169), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n324), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(G200), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(new_n323), .C1(new_n274), .C2(new_n349), .ZN(new_n353));
  INV_X1    g0153(.A(new_n291), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n354), .A2(new_n288), .B1(new_n210), .B2(new_n257), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(new_n317), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n294), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n257), .B1(new_n282), .B2(new_n283), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n280), .A2(new_n359), .B1(new_n257), .B2(new_n312), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G238), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n258), .A2(new_n362), .B1(new_n206), .B2(new_n254), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n333), .A2(new_n220), .A3(G1698), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n261), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n268), .B1(G244), .B2(new_n271), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n361), .B1(new_n368), .B2(G169), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n367), .A2(G179), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n361), .B1(new_n368), .B2(G190), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n311), .A2(new_n351), .A3(new_n353), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n291), .A2(new_n284), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n378), .A2(new_n279), .B1(new_n277), .B2(new_n291), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n252), .A2(KEYINPUT70), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT70), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT3), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n382), .A3(G33), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT69), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n250), .ZN(new_n385));
  NAND2_X1  g0185(.A1(KEYINPUT69), .A2(G33), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(KEYINPUT3), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(G20), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n202), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n383), .A2(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n210), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT7), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT71), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G58), .A2(G68), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n210), .B1(new_n203), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G159), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n288), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n395), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n396), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n286), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n315), .A2(G159), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(KEYINPUT71), .A3(new_n403), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n400), .A2(KEYINPUT16), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n295), .B1(new_n394), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n389), .A2(G20), .ZN(new_n408));
  AOI21_X1  g0208(.A(G33), .B1(new_n380), .B2(new_n382), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT3), .B1(new_n385), .B2(new_n386), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n389), .B1(new_n254), .B2(G20), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n202), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n402), .A2(new_n403), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n407), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n379), .B1(new_n406), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT72), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n259), .A2(new_n255), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n215), .A2(G1698), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n418), .B1(new_n391), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n261), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n267), .B1(new_n270), .B2(new_n220), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n274), .A3(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n383), .A2(new_n387), .A3(new_n419), .A4(new_n420), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n264), .B1(new_n427), .B2(new_n418), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n372), .B1(new_n428), .B2(new_n424), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT74), .B1(new_n416), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n391), .A2(new_n389), .A3(new_n210), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G68), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n388), .A2(new_n389), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n405), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n415), .A2(new_n435), .A3(new_n294), .ZN(new_n436));
  INV_X1    g0236(.A(new_n379), .ZN(new_n437));
  AND4_X1   g0237(.A1(KEYINPUT74), .A2(new_n436), .A3(new_n437), .A4(new_n430), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT17), .B1(new_n431), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(G169), .B1(new_n423), .B2(new_n425), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n428), .A2(G179), .A3(new_n424), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT73), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G179), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n423), .A2(new_n443), .A3(new_n425), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT73), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n307), .B1(new_n428), .B2(new_n424), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT18), .B1(new_n448), .B2(new_n416), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n436), .A2(new_n437), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT17), .B1(new_n416), .B2(new_n430), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n439), .A2(new_n449), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n377), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR4_X1   g0260(.A1(new_n333), .A2(KEYINPUT22), .A3(G20), .A4(new_n216), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n383), .A2(new_n387), .A3(new_n210), .A4(G87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT84), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT22), .B1(new_n463), .B2(KEYINPUT84), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g0267(.A1(KEYINPUT78), .A2(G116), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT78), .A2(G116), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n385), .A2(new_n386), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OR3_X1    g0272(.A1(new_n472), .A2(KEYINPUT86), .A3(G20), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT86), .B1(new_n472), .B2(G20), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT87), .B1(new_n206), .B2(G20), .ZN(new_n475));
  XOR2_X1   g0275(.A(new_n475), .B(KEYINPUT23), .Z(new_n476));
  AND3_X1   g0276(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g0277(.A(KEYINPUT85), .B(KEYINPUT24), .Z(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n467), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n467), .B2(new_n477), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n294), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT76), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n250), .B2(G1), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n209), .A2(KEYINPUT76), .A3(G33), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n279), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT25), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n277), .B2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n312), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n487), .A2(G107), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n482), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT88), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n265), .A2(G1), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  NOR2_X1   g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n264), .ZN(new_n498));
  INV_X1    g0298(.A(G264), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(KEYINPUT88), .A3(G264), .A4(new_n264), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n471), .A2(G294), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n221), .A2(G1698), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(G250), .B2(G1698), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n391), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n261), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT5), .B(G41), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(new_n264), .A3(G274), .A4(new_n494), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n502), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G169), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n502), .A2(new_n507), .A3(G179), .A4(new_n509), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n511), .A2(KEYINPUT89), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT89), .B1(new_n511), .B2(new_n512), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n492), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n510), .A2(G190), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n510), .A2(new_n372), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n482), .B(new_n491), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT77), .ZN(new_n521));
  INV_X1    g0321(.A(new_n408), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n380), .A2(new_n382), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n250), .ZN(new_n524));
  INV_X1    g0324(.A(new_n386), .ZN(new_n525));
  NOR2_X1   g0325(.A1(KEYINPUT69), .A2(G33), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n252), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n522), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT7), .B1(new_n333), .B2(new_n210), .ZN(new_n529));
  OAI21_X1  g0329(.A(G107), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g0330(.A(G97), .B(G107), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g0333(.A(KEYINPUT75), .B(G97), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n532), .A2(G107), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(G20), .B1(G77), .B2(new_n315), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n295), .B1(new_n530), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n277), .A2(G97), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n487), .B2(G97), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n521), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n537), .A2(G20), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n315), .A2(G77), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n206), .B1(new_n411), .B2(new_n412), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n294), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(KEYINPUT77), .A3(new_n541), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT4), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n255), .A2(G244), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n391), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G244), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n555), .A2(new_n255), .A3(new_n251), .A4(new_n253), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G283), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n251), .A2(new_n253), .A3(G250), .A4(G1698), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n264), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n509), .B1(new_n498), .B2(new_n221), .ZN(new_n561));
  OAI21_X1  g0361(.A(G169), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n561), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n383), .A2(new_n387), .A3(G244), .A4(new_n255), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n551), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n563), .B(G179), .C1(new_n566), .C2(new_n264), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n550), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(G200), .B1(new_n560), .B2(new_n561), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n563), .B(G190), .C1(new_n566), .C2(new_n264), .ZN(new_n571));
  AND4_X1   g0371(.A1(new_n548), .A2(new_n570), .A3(new_n541), .A4(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G238), .A2(G1698), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n554), .B2(G1698), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n383), .A2(new_n575), .A3(new_n387), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n472), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n261), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n494), .A2(new_n217), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n264), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n264), .A2(G274), .ZN(new_n581));
  INV_X1    g0381(.A(new_n494), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n578), .A2(G190), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n264), .B1(new_n576), .B2(new_n472), .ZN(new_n586));
  OAI21_X1  g0386(.A(G200), .B1(new_n586), .B2(new_n583), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n210), .B1(new_n336), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT79), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(KEYINPUT79), .B(new_n210), .C1(new_n336), .C2(new_n589), .ZN(new_n593));
  XNOR2_X1  g0393(.A(KEYINPUT80), .B(G87), .ZN(new_n594));
  OR2_X1    g0394(.A1(KEYINPUT75), .A2(G97), .ZN(new_n595));
  NAND2_X1  g0395(.A1(KEYINPUT75), .A2(G97), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n206), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n383), .A2(new_n387), .A3(new_n210), .A4(G68), .ZN(new_n599));
  XOR2_X1   g0399(.A(KEYINPUT75), .B(G97), .Z(new_n600));
  OAI21_X1  g0400(.A(new_n589), .B1(new_n600), .B2(new_n317), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n294), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n356), .A2(new_n312), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n487), .A2(G87), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n578), .A2(G179), .A3(new_n584), .ZN(new_n607));
  OAI21_X1  g0407(.A(G169), .B1(new_n586), .B2(new_n583), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n356), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT81), .B1(new_n487), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT81), .ZN(new_n612));
  NOR4_X1   g0412(.A1(new_n279), .A2(new_n486), .A3(new_n612), .A4(new_n356), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n603), .A2(new_n614), .A3(new_n604), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n588), .A2(new_n606), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n569), .A2(new_n573), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n557), .A2(new_n210), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n600), .B2(G33), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT20), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(KEYINPUT83), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n468), .A2(new_n469), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G20), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(KEYINPUT83), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n294), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n620), .A2(new_n622), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n294), .B(new_n625), .C1(new_n470), .C2(new_n210), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n618), .B1(new_n534), .B2(new_n250), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n628), .A2(new_n629), .B1(KEYINPUT83), .B2(new_n621), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n487), .A2(G116), .B1(new_n312), .B2(new_n623), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(G257), .A2(G1698), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n499), .B2(G1698), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n383), .A2(new_n636), .A3(new_n387), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n333), .A2(G303), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(KEYINPUT82), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT82), .B1(new_n637), .B2(new_n638), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n261), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n497), .A2(G270), .A3(new_n264), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n509), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n642), .A2(G190), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n641), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n639), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n648), .B2(new_n261), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n634), .B(new_n646), .C1(new_n649), .C2(new_n372), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT21), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n633), .A2(G169), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n642), .A2(new_n645), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n654), .A2(KEYINPUT21), .A3(G169), .A4(new_n633), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n644), .A2(new_n443), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n633), .A2(new_n642), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n650), .A2(new_n653), .A3(new_n655), .A4(new_n657), .ZN(new_n658));
  NOR4_X1   g0458(.A1(new_n460), .A2(new_n520), .A3(new_n617), .A4(new_n658), .ZN(G372));
  AND2_X1   g0459(.A1(new_n455), .A2(new_n449), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n436), .A2(new_n430), .A3(new_n437), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT74), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n416), .A2(KEYINPUT74), .A3(new_n430), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n456), .B1(new_n665), .B2(KEYINPUT17), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n348), .A2(new_n350), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n668), .A2(new_n324), .B1(new_n353), .B2(new_n371), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n660), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n304), .A3(new_n306), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n609), .A2(new_n615), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n602), .A2(new_n294), .B1(new_n312), .B2(new_n356), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n585), .A3(new_n605), .A4(new_n587), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n569), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n548), .A2(new_n541), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n672), .A2(new_n568), .A3(new_n674), .A4(new_n677), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n676), .B(new_n672), .C1(KEYINPUT26), .C2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT90), .ZN(new_n680));
  INV_X1    g0480(.A(new_n491), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT22), .ZN(new_n682));
  INV_X1    g0482(.A(new_n463), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT84), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n461), .B1(new_n685), .B2(new_n464), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n478), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n467), .A2(new_n477), .A3(new_n479), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n681), .B1(new_n690), .B2(new_n294), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n511), .A2(new_n512), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n680), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n653), .A2(new_n655), .A3(new_n657), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n492), .A2(KEYINPUT90), .A3(new_n692), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n543), .A2(new_n549), .B1(new_n562), .B2(new_n567), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n699), .A2(new_n572), .A3(new_n675), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n519), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n679), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n309), .B(new_n671), .C1(new_n460), .C2(new_n703), .ZN(G369));
  NAND3_X1  g0504(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(G213), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n634), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n695), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n658), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n516), .A2(new_n519), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n691), .B2(new_n711), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n492), .A2(new_n515), .A3(new_n710), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n694), .A2(new_n697), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n711), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n696), .A2(new_n710), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n720), .A2(new_n722), .A3(new_n724), .ZN(G399));
  INV_X1    g0525(.A(new_n225), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OR3_X1    g0528(.A1(new_n597), .A2(new_n594), .A3(G116), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(G1), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(new_n232), .B2(new_n728), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  OR3_X1    g0533(.A1(new_n703), .A2(KEYINPUT29), .A3(new_n710), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n586), .A2(new_n583), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G179), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n737), .B(new_n510), .C1(new_n560), .C2(new_n561), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n649), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT91), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n560), .A2(new_n561), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n642), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n736), .A2(new_n507), .A3(new_n502), .A4(new_n656), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n740), .B(KEYINPUT30), .C1(new_n742), .C2(new_n743), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n739), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n735), .B1(new_n748), .B2(new_n711), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n711), .A2(new_n735), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n700), .A2(new_n696), .A3(new_n650), .A4(new_n711), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n749), .B1(new_n748), .B2(new_n751), .C1(new_n752), .C2(new_n520), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT26), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n699), .A2(new_n755), .A3(new_n616), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n678), .A2(KEYINPUT26), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n756), .A2(new_n672), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n695), .B1(new_n492), .B2(new_n515), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n701), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n711), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(KEYINPUT29), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n734), .A2(new_n754), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n733), .B1(new_n764), .B2(G1), .ZN(G364));
  AND2_X1   g0565(.A1(new_n210), .A2(G13), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n209), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n727), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n714), .B2(G330), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G330), .B2(new_n714), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n769), .B(KEYINPUT92), .Z(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n228), .B1(G20), .B2(new_n307), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n225), .A2(new_n254), .ZN(new_n779));
  INV_X1    g0579(.A(G355), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n780), .B1(G116), .B2(new_n225), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n225), .A2(new_n391), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n265), .B2(new_n233), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n245), .A2(new_n265), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n772), .B1(new_n778), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n210), .A2(new_n274), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n443), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n210), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G58), .A2(new_n790), .B1(new_n793), .B2(G77), .ZN(new_n794));
  NAND3_X1  g0594(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n274), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n794), .B1(new_n214), .B2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT93), .Z(new_n799));
  NOR2_X1   g0599(.A1(G179), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n791), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G159), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT32), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n372), .A2(G179), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n787), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n333), .B1(new_n807), .B2(new_n594), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n791), .A2(new_n805), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n206), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n795), .A2(G190), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n202), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n210), .B1(new_n800), .B2(G190), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n205), .ZN(new_n815));
  NOR4_X1   g0615(.A1(new_n804), .A2(new_n810), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n799), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G303), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n333), .B1(new_n806), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n814), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(G294), .B2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G322), .A2(new_n790), .B1(new_n802), .B2(G329), .ZN(new_n822));
  INV_X1    g0622(.A(new_n809), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G283), .A2(new_n823), .B1(new_n793), .B2(G311), .ZN(new_n824));
  XNOR2_X1  g0624(.A(KEYINPUT33), .B(G317), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n811), .A2(new_n825), .B1(new_n796), .B2(G326), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n821), .A2(new_n822), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n817), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n786), .B1(new_n776), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n775), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n714), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n771), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  NOR3_X1   g0633(.A1(new_n369), .A2(new_n370), .A3(new_n710), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n374), .A2(new_n375), .B1(new_n361), .B2(new_n710), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n371), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n703), .B2(new_n710), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n376), .A2(new_n711), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n703), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n769), .B1(new_n840), .B2(new_n754), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n754), .B2(new_n840), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n776), .A2(new_n773), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT94), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n772), .B1(G77), .B2(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G68), .A2(new_n823), .B1(new_n802), .B2(G132), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n214), .B2(new_n806), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n391), .B(new_n847), .C1(G58), .C2(new_n820), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G143), .A2(new_n790), .B1(new_n793), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n797), .B2(new_n850), .C1(new_n289), .C2(new_n812), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n848), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(G311), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n809), .A2(new_n216), .B1(new_n801), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT95), .Z(new_n858));
  INV_X1    g0658(.A(G294), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n206), .A2(new_n806), .B1(new_n789), .B2(new_n859), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n254), .B(new_n860), .C1(new_n470), .C2(new_n793), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n796), .A2(G303), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n815), .B1(new_n811), .B2(G283), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n855), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n845), .B1(new_n865), .B2(new_n776), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n361), .A2(new_n710), .ZN(new_n867));
  INV_X1    g0667(.A(new_n375), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(new_n373), .ZN(new_n869));
  INV_X1    g0669(.A(new_n371), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n834), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n866), .B1(new_n871), .B2(new_n774), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT96), .Z(new_n873));
  NAND2_X1  g0673(.A1(new_n842), .A2(new_n873), .ZN(G384));
  OR2_X1    g0674(.A1(new_n537), .A2(KEYINPUT35), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n537), .A2(KEYINPUT35), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(G116), .A3(new_n229), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT36), .Z(new_n878));
  NAND3_X1  g0678(.A1(new_n233), .A2(G77), .A3(new_n396), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n214), .A2(G68), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n209), .B(G13), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n668), .A2(new_n324), .A3(new_n711), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n400), .B(new_n404), .C1(new_n433), .C2(new_n434), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n407), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n379), .B1(new_n885), .B2(new_n406), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(new_n708), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n458), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n448), .B2(new_n708), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n665), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT37), .B1(new_n452), .B2(new_n454), .ZN(new_n891));
  INV_X1    g0691(.A(new_n708), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n454), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n891), .A2(new_n663), .A3(new_n664), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n431), .A2(new_n438), .ZN(new_n900));
  INV_X1    g0700(.A(new_n886), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n452), .B2(new_n892), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n454), .A2(new_n442), .A3(new_n447), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(new_n899), .A3(new_n893), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(new_n665), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT38), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n887), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n666), .B2(new_n660), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n907), .A2(new_n909), .A3(KEYINPUT97), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT97), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n897), .B1(new_n890), .B2(new_n894), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n911), .B1(new_n888), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n898), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT39), .ZN(new_n915));
  INV_X1    g0715(.A(new_n893), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n458), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n904), .A2(new_n661), .A3(new_n893), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n894), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n907), .A2(new_n909), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT39), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n883), .B1(new_n915), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n835), .B1(new_n703), .B2(new_n839), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n323), .A2(new_n711), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n351), .A2(new_n353), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n351), .B2(new_n353), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT97), .B1(new_n907), .B2(new_n909), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n888), .A2(new_n912), .A3(new_n911), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n934), .A2(new_n935), .B1(new_n897), .B2(new_n896), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n933), .A2(new_n936), .B1(new_n660), .B2(new_n892), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT98), .B1(new_n925), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n883), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n934), .A2(new_n935), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n940), .B1(new_n941), .B2(new_n898), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n939), .B1(new_n942), .B2(new_n923), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n660), .A2(new_n892), .ZN(new_n944));
  INV_X1    g0744(.A(new_n933), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n944), .B1(new_n945), .B2(new_n914), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT98), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n938), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n671), .A2(new_n309), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n734), .A2(new_n762), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n459), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n949), .B(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(G330), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n351), .A2(new_n353), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n927), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n351), .A2(new_n353), .A3(new_n928), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n837), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT40), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n749), .B1(new_n752), .B2(new_n520), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT99), .B1(new_n748), .B2(new_n751), .ZN(new_n961));
  INV_X1    g0761(.A(new_n747), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n502), .A2(new_n656), .A3(new_n507), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n963), .A2(new_n741), .A3(new_n736), .A4(new_n642), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT30), .B1(new_n964), .B2(new_n740), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n962), .A2(new_n965), .B1(new_n649), .B2(new_n738), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT99), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n966), .A2(new_n967), .A3(new_n750), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n958), .B(new_n959), .C1(new_n960), .C2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n941), .B2(new_n898), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n893), .B1(new_n666), .B2(new_n660), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n894), .A2(new_n919), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n897), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n888), .A2(new_n912), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n871), .B1(new_n929), .B2(new_n930), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n617), .A2(new_n658), .A3(new_n710), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n966), .A2(new_n710), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n716), .A2(new_n978), .B1(new_n979), .B2(new_n735), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n961), .A2(new_n968), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n959), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n971), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n960), .A2(new_n969), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n460), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n954), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n986), .B2(new_n984), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n953), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n209), .B2(new_n766), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n953), .A2(new_n988), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n882), .B1(new_n990), .B2(new_n991), .ZN(G367));
  OAI221_X1 g0792(.A(new_n777), .B1(new_n225), .B2(new_n356), .C1(new_n782), .C2(new_n241), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n772), .A2(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G283), .A2(new_n793), .B1(new_n802), .B2(G317), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n807), .A2(KEYINPUT46), .A3(G116), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n391), .B1(new_n818), .B2(new_n789), .C1(new_n600), .C2(new_n809), .ZN(new_n998));
  XNOR2_X1  g0798(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n623), .B2(new_n806), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n206), .B2(new_n814), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n812), .A2(new_n859), .B1(new_n797), .B2(new_n856), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n820), .A2(G68), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1004), .B(new_n254), .C1(new_n201), .C2(new_n806), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n823), .A2(G77), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n289), .B2(new_n789), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n792), .A2(new_n214), .B1(new_n801), .B2(new_n850), .ZN(new_n1008));
  INV_X1    g0808(.A(G143), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n812), .A2(new_n398), .B1(new_n797), .B2(new_n1009), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1003), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  AOI21_X1  g0813(.A(new_n994), .B1(new_n1013), .B2(new_n776), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n606), .A2(new_n711), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1015), .A2(new_n609), .A3(new_n615), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n675), .B2(new_n1015), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(new_n830), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n717), .A2(new_n718), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n724), .B1(new_n1020), .B2(new_n723), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(new_n715), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1022), .A2(new_n763), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n677), .A2(new_n710), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n569), .A2(new_n573), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n568), .A2(new_n677), .A3(new_n710), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n722), .A2(new_n724), .A3(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT45), .Z(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n722), .B2(new_n724), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT44), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n719), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n720), .A3(new_n1031), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1023), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1035), .A2(KEYINPUT102), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(KEYINPUT102), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n764), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n727), .B(KEYINPUT41), .Z(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n768), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n716), .A2(new_n723), .A3(new_n1027), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT42), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1027), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n569), .B1(new_n1044), .B2(new_n516), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n711), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1042), .A2(KEYINPUT42), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1043), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n1048), .A2(KEYINPUT43), .A3(new_n1017), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1017), .B(KEYINPUT43), .Z(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n719), .A2(new_n1027), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT100), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1049), .B(new_n1051), .C1(new_n1053), .C2(KEYINPUT101), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(KEYINPUT101), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1054), .B(new_n1055), .Z(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1019), .B1(new_n1041), .B2(new_n1057), .ZN(G387));
  NOR2_X1   g0858(.A1(new_n1022), .A2(new_n767), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n717), .A2(new_n718), .A3(new_n775), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n238), .A2(new_n265), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1061), .A2(new_n782), .B1(new_n730), .B2(new_n779), .ZN(new_n1062));
  OR3_X1    g0862(.A1(new_n354), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT50), .B1(new_n354), .B2(G50), .ZN(new_n1064));
  AOI21_X1  g0864(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1063), .A2(new_n730), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1062), .A2(new_n1066), .B1(new_n206), .B2(new_n726), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n772), .B1(new_n1067), .B2(new_n778), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G317), .A2(new_n790), .B1(new_n793), .B2(G303), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT106), .B(G322), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1069), .B1(new_n797), .B2(new_n1070), .C1(new_n856), .C2(new_n812), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n807), .A2(G294), .B1(new_n820), .B2(G283), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT49), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n470), .A2(new_n823), .B1(new_n802), .B2(G326), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1078), .A2(new_n391), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n809), .A2(new_n205), .B1(new_n801), .B2(new_n289), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n806), .A2(new_n257), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1082), .A2(new_n1083), .A3(new_n391), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT104), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n814), .A2(new_n356), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G50), .B2(new_n790), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT105), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n291), .A2(new_n811), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n793), .A2(G68), .B1(G159), .B2(new_n796), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1081), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1068), .B1(new_n1092), .B2(new_n776), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1059), .B1(new_n1060), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT107), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1022), .B2(new_n763), .ZN(new_n1096));
  OR3_X1    g0896(.A1(new_n1096), .A2(new_n1023), .A3(new_n728), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1022), .A2(new_n1095), .A3(new_n763), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1094), .B1(new_n1097), .B2(new_n1098), .ZN(G393));
  NAND2_X1  g0899(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1023), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n728), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(KEYINPUT113), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT113), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1105), .B(new_n1102), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1100), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1044), .A2(new_n775), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT108), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n777), .B1(new_n225), .B2(new_n600), .C1(new_n782), .C2(new_n248), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n772), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT109), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n790), .A2(G311), .B1(G317), .B2(new_n796), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT52), .Z(new_n1115));
  OAI22_X1  g0915(.A1(new_n792), .A2(new_n859), .B1(new_n801), .B2(new_n1070), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G283), .B2(new_n807), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n333), .B1(new_n809), .B2(new_n206), .C1(new_n812), .C2(new_n818), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n470), .B2(new_n820), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT112), .Z(new_n1121));
  AOI22_X1  g0921(.A1(new_n790), .A2(G159), .B1(G150), .B2(new_n796), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT110), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(KEYINPUT51), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(KEYINPUT51), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n806), .A2(new_n202), .B1(new_n801), .B2(new_n1009), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT111), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n354), .A2(new_n792), .B1(new_n216), .B2(new_n809), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n812), .A2(new_n214), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n814), .A2(new_n257), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1128), .A2(new_n391), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1125), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1121), .B1(new_n1124), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1113), .B1(new_n776), .B2(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1108), .A2(new_n768), .B1(new_n1110), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1107), .A2(new_n1135), .ZN(G390));
  OAI21_X1  g0936(.A(new_n772), .B1(new_n291), .B2(new_n844), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n254), .B(new_n1130), .C1(G68), .C2(new_n823), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G87), .A2(new_n807), .B1(new_n790), .B2(G116), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n534), .A2(new_n793), .B1(new_n802), .B2(G294), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G107), .A2(new_n811), .B1(new_n796), .B2(G283), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n254), .B1(new_n809), .B2(new_n214), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G125), .B2(new_n802), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT117), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n807), .A2(G150), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1146), .A2(KEYINPUT53), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1146), .A2(KEYINPUT53), .B1(new_n796), .B2(G128), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n790), .A2(G132), .B1(new_n793), .B2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n820), .A2(G159), .B1(G137), .B2(new_n811), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1142), .B1(new_n1145), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1137), .B1(new_n776), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n923), .B1(KEYINPUT39), .B2(new_n914), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n1157), .B2(new_n774), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n933), .A2(new_n883), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n915), .A3(new_n924), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT114), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n883), .B1(new_n921), .B2(new_n922), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n869), .A2(new_n870), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n760), .A2(new_n711), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n931), .B1(new_n1164), .B2(new_n835), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1161), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n835), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n932), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n939), .B1(new_n974), .B2(new_n975), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(KEYINPUT114), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n753), .A2(new_n932), .A3(G330), .A4(new_n871), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1160), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1156), .A2(new_n1159), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n985), .A2(new_n954), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n958), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1173), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1158), .B1(new_n1177), .B2(new_n767), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT116), .ZN(new_n1179));
  OAI211_X1 g0979(.A(G330), .B(new_n871), .C1(new_n960), .C2(new_n969), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(KEYINPUT115), .A3(new_n931), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1167), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n1182), .A3(new_n1172), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT115), .B1(new_n1180), .B2(new_n931), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1179), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1182), .A2(new_n1172), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1184), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1186), .A2(new_n1187), .A3(KEYINPUT116), .A4(new_n1181), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n931), .B1(new_n754), .B2(new_n837), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1176), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n926), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n459), .A2(new_n1175), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n952), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n728), .B1(new_n1197), .B2(new_n1177), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1177), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1178), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(G378));
  OAI21_X1  g1002(.A(G330), .B1(new_n971), .B2(new_n983), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n296), .A2(new_n892), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT55), .Z(new_n1205));
  XNOR2_X1  g1005(.A(new_n310), .B(new_n1205), .ZN(new_n1206));
  XOR2_X1   g1006(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1206), .B(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1203), .A2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1209), .B(G330), .C1(new_n983), .C2(new_n971), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n925), .A2(KEYINPUT98), .A3(new_n937), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n947), .B1(new_n943), .B2(new_n946), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1213), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n938), .A2(new_n948), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1185), .A2(new_n1188), .B1(new_n926), .B2(new_n1191), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1196), .B1(new_n1177), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT57), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n728), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1218), .A2(new_n1220), .A3(KEYINPUT57), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT121), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1218), .A2(new_n1220), .A3(KEYINPUT121), .A4(KEYINPUT57), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n820), .A2(G150), .B1(G125), .B2(new_n796), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT119), .Z(new_n1230));
  INV_X1    g1030(.A(G128), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n789), .A2(new_n1231), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n806), .A2(new_n1149), .B1(new_n792), .B2(new_n850), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(G132), .C2(new_n811), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1230), .A2(new_n1234), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n802), .A2(G124), .ZN(new_n1238));
  AOI211_X1 g1038(.A(G33), .B(G41), .C1(new_n823), .C2(G159), .ZN(new_n1239));
  AND4_X1   g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n796), .A2(G116), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1004), .B(new_n1241), .C1(new_n205), .C2(new_n812), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n789), .A2(new_n206), .B1(new_n792), .B2(new_n356), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n809), .A2(new_n201), .ZN(new_n1244));
  INV_X1    g1044(.A(G283), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n801), .A2(new_n1245), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n391), .A2(new_n263), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT118), .B1(new_n1248), .B2(new_n1083), .ZN(new_n1249));
  OR3_X1    g1049(.A1(new_n1248), .A2(KEYINPUT118), .A3(new_n1083), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1247), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT58), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G50), .B1(new_n250), .B2(new_n263), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1251), .A2(new_n1252), .B1(new_n1248), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1252), .B2(new_n1251), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n776), .B1(new_n1240), .B2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(new_n769), .C1(G50), .C2(new_n844), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1209), .B2(new_n773), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1218), .B2(new_n768), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1228), .A2(new_n1259), .ZN(G375));
  NAND2_X1  g1060(.A1(new_n1219), .A2(new_n1195), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1197), .A2(new_n1040), .A3(new_n1261), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n767), .B(KEYINPUT122), .Z(new_n1263));
  NAND2_X1  g1063(.A1(new_n1193), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n772), .B1(G68), .B2(new_n844), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(G97), .A2(new_n807), .B1(new_n802), .B2(G303), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1266), .B1(new_n206), .B2(new_n792), .C1(new_n1245), .C2(new_n789), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n623), .A2(new_n812), .B1(new_n797), .B2(new_n859), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1006), .A2(new_n333), .ZN(new_n1269));
  NOR4_X1   g1069(.A1(new_n1267), .A2(new_n1086), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OR2_X1    g1071(.A1(new_n1271), .A2(KEYINPUT123), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n391), .B(new_n1244), .C1(G137), .C2(new_n790), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1150), .A2(new_n811), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n820), .A2(G50), .B1(G132), .B2(new_n796), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n792), .A2(new_n289), .B1(new_n801), .B2(new_n1231), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(G159), .B2(new_n807), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1271), .A2(KEYINPUT123), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1272), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1265), .B1(new_n1280), .B2(new_n776), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n932), .B2(new_n774), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1262), .A2(new_n1264), .A3(new_n1282), .ZN(G381));
  OAI211_X1 g1083(.A(new_n832), .B(new_n1094), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1284));
  NOR4_X1   g1084(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(G387), .A2(G378), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n1228), .A3(new_n1259), .A4(new_n1286), .ZN(G407));
  NAND2_X1  g1087(.A1(new_n709), .A2(G213), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1228), .A2(new_n1201), .A3(new_n1259), .A4(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(G407), .A2(G213), .A3(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(KEYINPUT124), .ZN(G409));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1228), .A2(G378), .A3(new_n1259), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1258), .B1(new_n1218), .B2(new_n1263), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1039), .B2(new_n1221), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1201), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1288), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1264), .B(new_n1282), .C1(new_n1300), .C2(G384), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1261), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1219), .A2(KEYINPUT60), .A3(new_n1195), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1304), .A2(new_n1197), .A3(new_n727), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G384), .A2(new_n1300), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1302), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1307), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1293), .B1(new_n1299), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1310), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1313), .A2(G2897), .A3(new_n1289), .A4(new_n1308), .ZN(new_n1314));
  INV_X1    g1114(.A(G2897), .ZN(new_n1315));
  OAI22_X1  g1115(.A1(new_n1309), .A2(new_n1310), .B1(new_n1315), .B2(new_n1288), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT61), .B1(new_n1299), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT126), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT102), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1108), .A2(new_n1320), .A3(new_n1023), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1035), .A2(KEYINPUT102), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n763), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n767), .B1(new_n1323), .B2(new_n1039), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1056), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1319), .B1(new_n1325), .B2(new_n1019), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1019), .ZN(new_n1327));
  AOI211_X1 g1127(.A(KEYINPUT126), .B(new_n1327), .C1(new_n1324), .C2(new_n1056), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G393), .A2(G396), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1284), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1107), .A2(new_n1135), .A3(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1330), .B1(new_n1107), .B2(new_n1135), .ZN(new_n1332));
  OAI22_X1  g1132(.A1(new_n1326), .A2(new_n1328), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1330), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G390), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(G387), .A2(KEYINPUT126), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1325), .A2(new_n1319), .A3(new_n1019), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1107), .A2(new_n1135), .A3(new_n1330), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1335), .A2(new_n1336), .A3(new_n1337), .A4(new_n1338), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1333), .A2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1289), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1311), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(KEYINPUT63), .A3(new_n1342), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1312), .A2(new_n1318), .A3(new_n1340), .A4(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT62), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1341), .A2(new_n1345), .A3(new_n1342), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT61), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1347), .B1(new_n1341), .B2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1345), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1346), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1344), .B1(new_n1351), .B2(new_n1340), .ZN(G405));
  INV_X1    g1152(.A(new_n1294), .ZN(new_n1353));
  AOI21_X1  g1153(.A(G378), .B1(new_n1228), .B2(new_n1259), .ZN(new_n1354));
  OAI21_X1  g1154(.A(KEYINPUT127), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(G375), .A2(new_n1201), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT127), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1356), .A2(new_n1357), .A3(new_n1294), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1355), .A2(new_n1358), .A3(new_n1311), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1356), .A2(new_n1342), .A3(new_n1357), .A4(new_n1294), .ZN(new_n1360));
  AND3_X1   g1160(.A1(new_n1359), .A2(new_n1340), .A3(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1340), .B1(new_n1360), .B2(new_n1359), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1361), .A2(new_n1362), .ZN(G402));
endmodule


