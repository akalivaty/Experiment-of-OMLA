

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(G2104), .A2(n522), .ZN(n887) );
  INV_X1 U553 ( .A(KEYINPUT92), .ZN(n660) );
  INV_X1 U554 ( .A(n646), .ZN(n681) );
  OR2_X1 U555 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U556 ( .A1(n634), .A2(n633), .ZN(n646) );
  BUF_X1 U557 ( .A(n646), .Z(n696) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n634) );
  NOR2_X1 U559 ( .A1(G651), .A2(n586), .ZN(n774) );
  OR2_X1 U560 ( .A1(n535), .A2(n534), .ZN(n536) );
  AND2_X1 U561 ( .A1(n528), .A2(n527), .ZN(G160) );
  AND2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n886) );
  NAND2_X1 U563 ( .A1(n886), .A2(G113), .ZN(n521) );
  INV_X1 U564 ( .A(G2105), .ZN(n522) );
  AND2_X1 U565 ( .A1(G2104), .A2(n522), .ZN(n518) );
  XNOR2_X2 U566 ( .A(n518), .B(KEYINPUT64), .ZN(n891) );
  NAND2_X1 U567 ( .A1(n891), .A2(G101), .ZN(n519) );
  XOR2_X1 U568 ( .A(n519), .B(KEYINPUT23), .Z(n520) );
  AND2_X1 U569 ( .A1(n521), .A2(n520), .ZN(n528) );
  NAND2_X1 U570 ( .A1(G125), .A2(n887), .ZN(n526) );
  XNOR2_X1 U571 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n524) );
  NOR2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XNOR2_X2 U573 ( .A(n524), .B(n523), .ZN(n890) );
  NAND2_X1 U574 ( .A1(G137), .A2(n890), .ZN(n525) );
  AND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U576 ( .A1(G114), .A2(n886), .ZN(n530) );
  NAND2_X1 U577 ( .A1(G126), .A2(n887), .ZN(n529) );
  NAND2_X1 U578 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U579 ( .A(KEYINPUT84), .B(n531), .ZN(n535) );
  NAND2_X1 U580 ( .A1(n890), .A2(G138), .ZN(n533) );
  NAND2_X1 U581 ( .A1(G102), .A2(n891), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U583 ( .A(KEYINPUT85), .B(n536), .ZN(G164) );
  INV_X1 U584 ( .A(G651), .ZN(n540) );
  NOR2_X1 U585 ( .A1(G543), .A2(n540), .ZN(n537) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n537), .Z(n775) );
  NAND2_X1 U587 ( .A1(G64), .A2(n775), .ZN(n539) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n586) );
  NAND2_X1 U589 ( .A1(G52), .A2(n774), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n539), .A2(n538), .ZN(n545) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n779) );
  NAND2_X1 U592 ( .A1(G90), .A2(n779), .ZN(n542) );
  NOR2_X1 U593 ( .A1(n586), .A2(n540), .ZN(n776) );
  NAND2_X1 U594 ( .A1(G77), .A2(n776), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U596 ( .A(KEYINPUT9), .B(n543), .Z(n544) );
  NOR2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U598 ( .A(KEYINPUT66), .B(n546), .ZN(G171) );
  INV_X1 U599 ( .A(G171), .ZN(G301) );
  NAND2_X1 U600 ( .A1(G85), .A2(n779), .ZN(n548) );
  NAND2_X1 U601 ( .A1(G72), .A2(n776), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U603 ( .A1(G60), .A2(n775), .ZN(n550) );
  NAND2_X1 U604 ( .A1(G47), .A2(n774), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n551) );
  OR2_X1 U606 ( .A1(n552), .A2(n551), .ZN(G290) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U608 ( .A1(G65), .A2(n775), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G53), .A2(n774), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U611 ( .A1(G91), .A2(n779), .ZN(n556) );
  NAND2_X1 U612 ( .A1(G78), .A2(n776), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n773) );
  INV_X1 U615 ( .A(n773), .ZN(G299) );
  INV_X1 U616 ( .A(G120), .ZN(G236) );
  INV_X1 U617 ( .A(G69), .ZN(G235) );
  INV_X1 U618 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U619 ( .A(KEYINPUT7), .B(KEYINPUT72), .ZN(n571) );
  NAND2_X1 U620 ( .A1(n779), .A2(G89), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U622 ( .A1(G76), .A2(n776), .ZN(n560) );
  NAND2_X1 U623 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n562), .B(KEYINPUT5), .ZN(n569) );
  XNOR2_X1 U625 ( .A(KEYINPUT71), .B(KEYINPUT6), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n775), .A2(G63), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(KEYINPUT70), .ZN(n565) );
  NAND2_X1 U628 ( .A1(G51), .A2(n774), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U632 ( .A(n571), .B(n570), .ZN(G168) );
  XOR2_X1 U633 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U634 ( .A1(G61), .A2(n775), .ZN(n573) );
  NAND2_X1 U635 ( .A1(G86), .A2(n779), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n776), .A2(G73), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT2), .B(n574), .Z(n575) );
  NOR2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n774), .A2(G48), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(G305) );
  NAND2_X1 U642 ( .A1(G88), .A2(n779), .ZN(n580) );
  NAND2_X1 U643 ( .A1(G75), .A2(n776), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT78), .B(n581), .Z(n585) );
  NAND2_X1 U646 ( .A1(G62), .A2(n775), .ZN(n583) );
  NAND2_X1 U647 ( .A1(G50), .A2(n774), .ZN(n582) );
  AND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(G303) );
  NAND2_X1 U650 ( .A1(G87), .A2(n586), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G74), .A2(G651), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U653 ( .A1(n775), .A2(n589), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G49), .A2(n774), .ZN(n590) );
  XOR2_X1 U655 ( .A(KEYINPUT77), .B(n590), .Z(n591) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(G288) );
  INV_X1 U657 ( .A(KEYINPUT40), .ZN(n749) );
  NAND2_X1 U658 ( .A1(G160), .A2(G40), .ZN(n632) );
  NOR2_X1 U659 ( .A1(n634), .A2(n632), .ZN(n739) );
  NAND2_X1 U660 ( .A1(G105), .A2(n891), .ZN(n593) );
  XNOR2_X1 U661 ( .A(n593), .B(KEYINPUT38), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G117), .A2(n886), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U664 ( .A1(G129), .A2(n887), .ZN(n596) );
  XNOR2_X1 U665 ( .A(KEYINPUT89), .B(n596), .ZN(n597) );
  NOR2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U667 ( .A(n599), .B(KEYINPUT90), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G141), .A2(n890), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n601), .A2(n600), .ZN(n876) );
  NOR2_X1 U670 ( .A1(G1996), .A2(n876), .ZN(n1007) );
  NAND2_X1 U671 ( .A1(G107), .A2(n886), .ZN(n603) );
  NAND2_X1 U672 ( .A1(G95), .A2(n891), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U674 ( .A1(G119), .A2(n887), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G131), .A2(n890), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  OR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n877) );
  XNOR2_X1 U678 ( .A(KEYINPUT88), .B(G1991), .ZN(n944) );
  NOR2_X1 U679 ( .A1(n877), .A2(n944), .ZN(n1000) );
  NOR2_X1 U680 ( .A1(G1986), .A2(G290), .ZN(n608) );
  XOR2_X1 U681 ( .A(n608), .B(KEYINPUT97), .Z(n609) );
  NOR2_X1 U682 ( .A1(n1000), .A2(n609), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n877), .A2(n944), .ZN(n611) );
  NAND2_X1 U684 ( .A1(G1996), .A2(n876), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n1005) );
  NOR2_X1 U686 ( .A1(n612), .A2(n1005), .ZN(n613) );
  NOR2_X1 U687 ( .A1(n1007), .A2(n613), .ZN(n614) );
  XNOR2_X1 U688 ( .A(KEYINPUT39), .B(n614), .ZN(n626) );
  XNOR2_X1 U689 ( .A(KEYINPUT37), .B(G2067), .ZN(n627) );
  NAND2_X1 U690 ( .A1(G104), .A2(n891), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(KEYINPUT86), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G140), .A2(n890), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n619) );
  XOR2_X1 U694 ( .A(KEYINPUT87), .B(KEYINPUT34), .Z(n618) );
  XNOR2_X1 U695 ( .A(n619), .B(n618), .ZN(n624) );
  NAND2_X1 U696 ( .A1(G116), .A2(n886), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G128), .A2(n887), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U699 ( .A(KEYINPUT35), .B(n622), .Z(n623) );
  NOR2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U701 ( .A(KEYINPUT36), .B(n625), .ZN(n873) );
  NOR2_X1 U702 ( .A1(n627), .A2(n873), .ZN(n1013) );
  NAND2_X1 U703 ( .A1(n739), .A2(n1013), .ZN(n741) );
  NAND2_X1 U704 ( .A1(n626), .A2(n741), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n873), .A2(n627), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT98), .ZN(n997) );
  NAND2_X1 U707 ( .A1(n629), .A2(n997), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n739), .A2(n630), .ZN(n631) );
  XNOR2_X1 U709 ( .A(KEYINPUT99), .B(n631), .ZN(n747) );
  INV_X1 U710 ( .A(n632), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G8), .A2(n696), .ZN(n732) );
  NOR2_X1 U712 ( .A1(G1981), .A2(G305), .ZN(n635) );
  XOR2_X1 U713 ( .A(n635), .B(KEYINPUT24), .Z(n636) );
  NOR2_X1 U714 ( .A1(n732), .A2(n636), .ZN(n737) );
  NAND2_X1 U715 ( .A1(G56), .A2(n775), .ZN(n637) );
  XOR2_X1 U716 ( .A(KEYINPUT14), .B(n637), .Z(n643) );
  NAND2_X1 U717 ( .A1(n779), .A2(G81), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n638), .B(KEYINPUT12), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G68), .A2(n776), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U721 ( .A(KEYINPUT13), .B(n641), .Z(n642) );
  NOR2_X1 U722 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n774), .A2(G43), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n920) );
  NAND2_X1 U725 ( .A1(G1996), .A2(n681), .ZN(n647) );
  XOR2_X1 U726 ( .A(n647), .B(KEYINPUT26), .Z(n648) );
  NOR2_X1 U727 ( .A1(n920), .A2(n648), .ZN(n650) );
  NAND2_X1 U728 ( .A1(G1341), .A2(n696), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n666) );
  NAND2_X1 U730 ( .A1(G54), .A2(n774), .ZN(n657) );
  NAND2_X1 U731 ( .A1(G66), .A2(n775), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G79), .A2(n776), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n779), .A2(G92), .ZN(n653) );
  XOR2_X1 U735 ( .A(KEYINPUT68), .B(n653), .Z(n654) );
  NOR2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n658), .B(KEYINPUT15), .ZN(n659) );
  XNOR2_X1 U739 ( .A(KEYINPUT69), .B(n659), .ZN(n918) );
  NOR2_X1 U740 ( .A1(n666), .A2(n918), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n661), .B(n660), .ZN(n665) );
  NAND2_X1 U742 ( .A1(G1348), .A2(n696), .ZN(n663) );
  XOR2_X2 U743 ( .A(n681), .B(KEYINPUT91), .Z(n679) );
  NAND2_X1 U744 ( .A1(G2067), .A2(n679), .ZN(n662) );
  NAND2_X1 U745 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U746 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n666), .A2(n918), .ZN(n667) );
  NAND2_X1 U748 ( .A1(n668), .A2(n667), .ZN(n673) );
  NAND2_X1 U749 ( .A1(n679), .A2(G2072), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(KEYINPUT27), .ZN(n671) );
  INV_X1 U751 ( .A(G1956), .ZN(n971) );
  NOR2_X1 U752 ( .A1(n971), .A2(n679), .ZN(n670) );
  NOR2_X1 U753 ( .A1(n671), .A2(n670), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n773), .A2(n674), .ZN(n672) );
  NAND2_X1 U755 ( .A1(n673), .A2(n672), .ZN(n677) );
  NOR2_X1 U756 ( .A1(n773), .A2(n674), .ZN(n675) );
  XOR2_X1 U757 ( .A(n675), .B(KEYINPUT28), .Z(n676) );
  NAND2_X1 U758 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U759 ( .A(n678), .B(KEYINPUT29), .ZN(n685) );
  XOR2_X1 U760 ( .A(G2078), .B(KEYINPUT25), .Z(n940) );
  INV_X1 U761 ( .A(n679), .ZN(n680) );
  NOR2_X1 U762 ( .A1(n940), .A2(n680), .ZN(n683) );
  NOR2_X1 U763 ( .A1(n681), .A2(G1961), .ZN(n682) );
  NOR2_X1 U764 ( .A1(n683), .A2(n682), .ZN(n687) );
  NOR2_X1 U765 ( .A1(G301), .A2(n687), .ZN(n684) );
  NOR2_X1 U766 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U767 ( .A(n686), .B(KEYINPUT93), .ZN(n709) );
  NAND2_X1 U768 ( .A1(G301), .A2(n687), .ZN(n688) );
  XNOR2_X1 U769 ( .A(KEYINPUT95), .B(n688), .ZN(n694) );
  NOR2_X1 U770 ( .A1(G1966), .A2(n732), .ZN(n711) );
  NOR2_X1 U771 ( .A1(G2084), .A2(n696), .ZN(n710) );
  NOR2_X1 U772 ( .A1(n711), .A2(n710), .ZN(n689) );
  NAND2_X1 U773 ( .A1(G8), .A2(n689), .ZN(n690) );
  XNOR2_X1 U774 ( .A(KEYINPUT30), .B(n690), .ZN(n691) );
  NOR2_X1 U775 ( .A1(G168), .A2(n691), .ZN(n692) );
  XNOR2_X1 U776 ( .A(n692), .B(KEYINPUT94), .ZN(n693) );
  NOR2_X1 U777 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U778 ( .A(KEYINPUT31), .B(n695), .Z(n708) );
  INV_X1 U779 ( .A(G8), .ZN(n701) );
  NOR2_X1 U780 ( .A1(G1971), .A2(n732), .ZN(n698) );
  NOR2_X1 U781 ( .A1(G2090), .A2(n696), .ZN(n697) );
  NOR2_X1 U782 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U783 ( .A1(n699), .A2(G303), .ZN(n700) );
  OR2_X1 U784 ( .A1(n701), .A2(n700), .ZN(n703) );
  AND2_X1 U785 ( .A1(n708), .A2(n703), .ZN(n702) );
  NAND2_X1 U786 ( .A1(n709), .A2(n702), .ZN(n706) );
  INV_X1 U787 ( .A(n703), .ZN(n704) );
  OR2_X1 U788 ( .A1(n704), .A2(G286), .ZN(n705) );
  NAND2_X1 U789 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U790 ( .A(n707), .B(KEYINPUT32), .ZN(n716) );
  AND2_X1 U791 ( .A1(n709), .A2(n708), .ZN(n714) );
  AND2_X1 U792 ( .A1(G8), .A2(n710), .ZN(n712) );
  OR2_X1 U793 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U794 ( .A1(n716), .A2(n715), .ZN(n731) );
  NOR2_X1 U795 ( .A1(G1976), .A2(G288), .ZN(n722) );
  NOR2_X1 U796 ( .A1(G1971), .A2(G303), .ZN(n717) );
  NOR2_X1 U797 ( .A1(n722), .A2(n717), .ZN(n933) );
  INV_X1 U798 ( .A(KEYINPUT33), .ZN(n718) );
  AND2_X1 U799 ( .A1(n933), .A2(n718), .ZN(n719) );
  NAND2_X1 U800 ( .A1(n731), .A2(n719), .ZN(n727) );
  INV_X1 U801 ( .A(n732), .ZN(n720) );
  NAND2_X1 U802 ( .A1(G1976), .A2(G288), .ZN(n929) );
  AND2_X1 U803 ( .A1(n720), .A2(n929), .ZN(n721) );
  NOR2_X1 U804 ( .A1(KEYINPUT33), .A2(n721), .ZN(n725) );
  NAND2_X1 U805 ( .A1(n722), .A2(KEYINPUT33), .ZN(n723) );
  NOR2_X1 U806 ( .A1(n732), .A2(n723), .ZN(n724) );
  NOR2_X1 U807 ( .A1(n725), .A2(n724), .ZN(n726) );
  AND2_X1 U808 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U809 ( .A(G1981), .B(G305), .Z(n915) );
  NAND2_X1 U810 ( .A1(n728), .A2(n915), .ZN(n735) );
  NOR2_X1 U811 ( .A1(G2090), .A2(G303), .ZN(n729) );
  NAND2_X1 U812 ( .A1(G8), .A2(n729), .ZN(n730) );
  NAND2_X1 U813 ( .A1(n731), .A2(n730), .ZN(n733) );
  NAND2_X1 U814 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U815 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U816 ( .A1(n737), .A2(n736), .ZN(n744) );
  XOR2_X1 U817 ( .A(G1986), .B(G290), .Z(n930) );
  INV_X1 U818 ( .A(n1005), .ZN(n738) );
  NAND2_X1 U819 ( .A1(n930), .A2(n738), .ZN(n740) );
  NAND2_X1 U820 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U821 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U822 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U823 ( .A(n745), .B(KEYINPUT96), .ZN(n746) );
  NOR2_X1 U824 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U825 ( .A(n749), .B(n748), .ZN(G329) );
  NAND2_X1 U826 ( .A1(G7), .A2(G661), .ZN(n750) );
  XNOR2_X1 U827 ( .A(n750), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U828 ( .A(G223), .ZN(n814) );
  NAND2_X1 U829 ( .A1(n814), .A2(G567), .ZN(n751) );
  XNOR2_X1 U830 ( .A(n751), .B(KEYINPUT67), .ZN(n752) );
  XNOR2_X1 U831 ( .A(KEYINPUT11), .B(n752), .ZN(G234) );
  INV_X1 U832 ( .A(G860), .ZN(n757) );
  OR2_X1 U833 ( .A1(n920), .A2(n757), .ZN(G153) );
  NAND2_X1 U834 ( .A1(G301), .A2(G868), .ZN(n754) );
  INV_X1 U835 ( .A(G868), .ZN(n795) );
  NAND2_X1 U836 ( .A1(n918), .A2(n795), .ZN(n753) );
  NAND2_X1 U837 ( .A1(n754), .A2(n753), .ZN(G284) );
  NAND2_X1 U838 ( .A1(G868), .A2(G286), .ZN(n756) );
  NAND2_X1 U839 ( .A1(G299), .A2(n795), .ZN(n755) );
  NAND2_X1 U840 ( .A1(n756), .A2(n755), .ZN(G297) );
  NAND2_X1 U841 ( .A1(n757), .A2(G559), .ZN(n758) );
  INV_X1 U842 ( .A(n918), .ZN(n792) );
  NAND2_X1 U843 ( .A1(n758), .A2(n792), .ZN(n759) );
  XNOR2_X1 U844 ( .A(n759), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U845 ( .A1(G868), .A2(n920), .ZN(n762) );
  NAND2_X1 U846 ( .A1(G868), .A2(n792), .ZN(n760) );
  NOR2_X1 U847 ( .A1(G559), .A2(n760), .ZN(n761) );
  NOR2_X1 U848 ( .A1(n762), .A2(n761), .ZN(G282) );
  NAND2_X1 U849 ( .A1(G111), .A2(n886), .ZN(n764) );
  NAND2_X1 U850 ( .A1(G99), .A2(n891), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n770) );
  NAND2_X1 U852 ( .A1(n887), .A2(G123), .ZN(n765) );
  XNOR2_X1 U853 ( .A(n765), .B(KEYINPUT18), .ZN(n767) );
  NAND2_X1 U854 ( .A1(G135), .A2(n890), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U856 ( .A(KEYINPUT73), .B(n768), .Z(n769) );
  NOR2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n999) );
  XNOR2_X1 U858 ( .A(n999), .B(G2096), .ZN(n772) );
  INV_X1 U859 ( .A(G2100), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(G156) );
  INV_X1 U861 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U862 ( .A(n773), .B(G288), .ZN(n791) );
  NAND2_X1 U863 ( .A1(G55), .A2(n774), .ZN(n784) );
  NAND2_X1 U864 ( .A1(G67), .A2(n775), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G80), .A2(n776), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G93), .A2(n779), .ZN(n780) );
  XNOR2_X1 U868 ( .A(KEYINPUT75), .B(n780), .ZN(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U871 ( .A(n785), .B(KEYINPUT76), .ZN(n824) );
  XNOR2_X1 U872 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n787) );
  XNOR2_X1 U873 ( .A(G290), .B(G166), .ZN(n786) );
  XNOR2_X1 U874 ( .A(n787), .B(n786), .ZN(n788) );
  XNOR2_X1 U875 ( .A(n824), .B(n788), .ZN(n789) );
  XNOR2_X1 U876 ( .A(n789), .B(G305), .ZN(n790) );
  XNOR2_X1 U877 ( .A(n791), .B(n790), .ZN(n901) );
  NAND2_X1 U878 ( .A1(G559), .A2(n792), .ZN(n793) );
  XOR2_X1 U879 ( .A(n920), .B(n793), .Z(n821) );
  XOR2_X1 U880 ( .A(n901), .B(n821), .Z(n794) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n797) );
  NOR2_X1 U882 ( .A1(n824), .A2(G868), .ZN(n796) );
  NOR2_X1 U883 ( .A1(n797), .A2(n796), .ZN(G295) );
  NAND2_X1 U884 ( .A1(G2078), .A2(G2084), .ZN(n798) );
  XOR2_X1 U885 ( .A(KEYINPUT20), .B(n798), .Z(n799) );
  NAND2_X1 U886 ( .A1(G2090), .A2(n799), .ZN(n801) );
  XNOR2_X1 U887 ( .A(KEYINPUT80), .B(KEYINPUT21), .ZN(n800) );
  XNOR2_X1 U888 ( .A(n801), .B(n800), .ZN(n802) );
  NAND2_X1 U889 ( .A1(G2072), .A2(n802), .ZN(G158) );
  XNOR2_X1 U890 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U891 ( .A1(G235), .A2(G236), .ZN(n803) );
  XNOR2_X1 U892 ( .A(n803), .B(KEYINPUT83), .ZN(n804) );
  NOR2_X1 U893 ( .A1(G237), .A2(n804), .ZN(n805) );
  NAND2_X1 U894 ( .A1(G108), .A2(n805), .ZN(n825) );
  NAND2_X1 U895 ( .A1(G567), .A2(n825), .ZN(n812) );
  XOR2_X1 U896 ( .A(KEYINPUT22), .B(KEYINPUT81), .Z(n807) );
  NAND2_X1 U897 ( .A1(G132), .A2(G82), .ZN(n806) );
  XNOR2_X1 U898 ( .A(n807), .B(n806), .ZN(n808) );
  NOR2_X1 U899 ( .A1(n808), .A2(G218), .ZN(n809) );
  XNOR2_X1 U900 ( .A(KEYINPUT82), .B(n809), .ZN(n810) );
  NAND2_X1 U901 ( .A1(n810), .A2(G96), .ZN(n826) );
  NAND2_X1 U902 ( .A1(G2106), .A2(n826), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n907) );
  NAND2_X1 U904 ( .A1(G661), .A2(G483), .ZN(n813) );
  NOR2_X1 U905 ( .A1(n907), .A2(n813), .ZN(n818) );
  NAND2_X1 U906 ( .A1(n818), .A2(G36), .ZN(G176) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n814), .ZN(G217) );
  INV_X1 U908 ( .A(G661), .ZN(n816) );
  NAND2_X1 U909 ( .A1(G2), .A2(G15), .ZN(n815) );
  NOR2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U911 ( .A(KEYINPUT102), .B(n817), .Z(G259) );
  NAND2_X1 U912 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U914 ( .A(KEYINPUT103), .B(n820), .Z(G188) );
  XOR2_X1 U915 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  XOR2_X1 U917 ( .A(n821), .B(KEYINPUT74), .Z(n822) );
  NOR2_X1 U918 ( .A1(G860), .A2(n822), .ZN(n823) );
  XOR2_X1 U919 ( .A(n824), .B(n823), .Z(G145) );
  INV_X1 U920 ( .A(G132), .ZN(G219) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  INV_X1 U922 ( .A(G82), .ZN(G220) );
  NOR2_X1 U923 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U925 ( .A(G2454), .B(G2446), .ZN(n835) );
  XNOR2_X1 U926 ( .A(G2430), .B(G2443), .ZN(n833) );
  XOR2_X1 U927 ( .A(G2435), .B(KEYINPUT100), .Z(n828) );
  XNOR2_X1 U928 ( .A(G2451), .B(G2438), .ZN(n827) );
  XNOR2_X1 U929 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U930 ( .A(n829), .B(G2427), .Z(n831) );
  XNOR2_X1 U931 ( .A(G1341), .B(G1348), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  NAND2_X1 U935 ( .A1(n836), .A2(G14), .ZN(n837) );
  XNOR2_X1 U936 ( .A(KEYINPUT101), .B(n837), .ZN(G401) );
  XOR2_X1 U937 ( .A(G2100), .B(G2678), .Z(n839) );
  XNOR2_X1 U938 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2090), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U944 ( .A(KEYINPUT105), .B(G2096), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n847) );
  XOR2_X1 U946 ( .A(G2078), .B(G2084), .Z(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1971), .B(G1961), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1966), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(G1981), .B(G1956), .Z(n851) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n857) );
  XOR2_X1 U957 ( .A(G1976), .B(G2474), .Z(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G136), .A2(n890), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n858), .B(KEYINPUT108), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G124), .A2(n887), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n859), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G112), .A2(n886), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G100), .A2(n891), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U968 ( .A1(n890), .A2(G139), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G103), .A2(n891), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G115), .A2(n886), .ZN(n869) );
  NAND2_X1 U972 ( .A1(G127), .A2(n887), .ZN(n868) );
  NAND2_X1 U973 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n870), .Z(n871) );
  NOR2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n992) );
  XNOR2_X1 U976 ( .A(n873), .B(n992), .ZN(n875) );
  XNOR2_X1 U977 ( .A(G164), .B(G160), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n880) );
  XNOR2_X1 U979 ( .A(G162), .B(n876), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U981 ( .A(n880), .B(n879), .Z(n885) );
  XOR2_X1 U982 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n882) );
  XNOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT111), .ZN(n881) );
  XNOR2_X1 U984 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U985 ( .A(KEYINPUT46), .B(n883), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n899) );
  NAND2_X1 U987 ( .A1(G118), .A2(n886), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G130), .A2(n887), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U990 ( .A1(n890), .A2(G142), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G106), .A2(n891), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U993 ( .A(KEYINPUT45), .B(n894), .Z(n895) );
  NOR2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n999), .B(n897), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U997 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U998 ( .A(n901), .B(G286), .ZN(n904) );
  XOR2_X1 U999 ( .A(KEYINPUT112), .B(n918), .Z(n902) );
  XNOR2_X1 U1000 ( .A(n920), .B(n902), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n905), .B(G301), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n906), .ZN(G397) );
  XOR2_X1 U1004 ( .A(KEYINPUT104), .B(n907), .Z(G319) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n908) );
  XOR2_X1 U1006 ( .A(KEYINPUT49), .B(n908), .Z(n909) );
  XNOR2_X1 U1007 ( .A(n909), .B(KEYINPUT113), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n910), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n911) );
  AND2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n913), .A2(G319), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1013 ( .A(G16), .B(KEYINPUT56), .Z(n938) );
  XOR2_X1 U1014 ( .A(G1966), .B(KEYINPUT123), .Z(n914) );
  XNOR2_X1 U1015 ( .A(G168), .B(n914), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n917), .B(KEYINPUT57), .ZN(n928) );
  XNOR2_X1 U1018 ( .A(G1348), .B(KEYINPUT124), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n919), .B(n918), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(G1341), .B(n920), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(G1971), .A2(G303), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(G1961), .B(G301), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n936) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(G1956), .B(G299), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n963) );
  XOR2_X1 U1033 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n959) );
  XNOR2_X1 U1034 ( .A(G2090), .B(G35), .ZN(n953) );
  XOR2_X1 U1035 ( .A(G2067), .B(G26), .Z(n939) );
  NAND2_X1 U1036 ( .A1(G28), .A2(n939), .ZN(n950) );
  XNOR2_X1 U1037 ( .A(G1996), .B(G32), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(n940), .B(G27), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1040 ( .A(KEYINPUT119), .B(n943), .Z(n948) );
  XNOR2_X1 U1041 ( .A(n944), .B(G25), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G2072), .B(G33), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT53), .B(n951), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n957) );
  XOR2_X1 U1048 ( .A(KEYINPUT120), .B(G34), .Z(n955) );
  XNOR2_X1 U1049 ( .A(G2084), .B(KEYINPUT54), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(n955), .B(n954), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(n959), .B(n958), .ZN(n960) );
  NOR2_X1 U1053 ( .A1(G29), .A2(n960), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(KEYINPUT122), .B(n961), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n964), .ZN(n990) );
  XNOR2_X1 U1057 ( .A(G1971), .B(G22), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G23), .B(G1976), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n968) );
  XOR2_X1 U1060 ( .A(G1986), .B(G24), .Z(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n970) );
  XOR2_X1 U1062 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n969) );
  XNOR2_X1 U1063 ( .A(n970), .B(n969), .ZN(n986) );
  XNOR2_X1 U1064 ( .A(G1961), .B(G5), .ZN(n984) );
  XNOR2_X1 U1065 ( .A(G20), .B(n971), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(G1341), .B(G19), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(G1981), .B(G6), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n978) );
  XOR2_X1 U1070 ( .A(KEYINPUT59), .B(G1348), .Z(n976) );
  XNOR2_X1 U1071 ( .A(G4), .B(n976), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1073 ( .A(KEYINPUT60), .B(n979), .Z(n981) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G21), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT125), .B(n982), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT61), .B(n987), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(G16), .A2(n988), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(n991), .B(KEYINPUT127), .ZN(n1022) );
  INV_X1 U1083 ( .A(G29), .ZN(n1020) );
  XOR2_X1 U1084 ( .A(G2072), .B(n992), .Z(n994) );
  XOR2_X1 U1085 ( .A(G164), .B(G2078), .Z(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n995), .B(KEYINPUT118), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(n996), .B(KEYINPUT50), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1016) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(G160), .B(G2084), .Z(n1001) );
  XNOR2_X1 U1092 ( .A(KEYINPUT115), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1011) );
  XOR2_X1 U1095 ( .A(G2090), .B(G162), .Z(n1006) );
  XNOR2_X1 U1096 ( .A(KEYINPUT116), .B(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(KEYINPUT51), .B(n1009), .Z(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(n1014), .B(KEYINPUT117), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(KEYINPUT52), .B(n1017), .Z(n1018) );
  NOR2_X1 U1104 ( .A1(KEYINPUT55), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .ZN(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

