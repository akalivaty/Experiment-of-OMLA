

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590;

  XOR2_X1 U318 ( .A(G176GAT), .B(G64GAT), .Z(n361) );
  XNOR2_X1 U319 ( .A(n404), .B(n359), .ZN(n360) );
  NOR2_X1 U320 ( .A1(n587), .A2(n453), .ZN(n456) );
  XOR2_X1 U321 ( .A(n365), .B(n364), .Z(n526) );
  XNOR2_X1 U322 ( .A(n405), .B(n391), .ZN(n523) );
  NOR2_X1 U323 ( .A1(n547), .A2(n481), .ZN(n286) );
  XOR2_X1 U324 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n287) );
  XNOR2_X1 U325 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U326 ( .A(n295), .B(n294), .ZN(n298) );
  NOR2_X1 U327 ( .A1(n535), .A2(n562), .ZN(n426) );
  XNOR2_X1 U328 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U329 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n473) );
  NOR2_X1 U330 ( .A1(n436), .A2(n435), .ZN(n492) );
  XNOR2_X1 U331 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U332 ( .A(KEYINPUT65), .B(KEYINPUT41), .ZN(n461) );
  XNOR2_X1 U333 ( .A(n474), .B(n473), .ZN(n536) );
  XNOR2_X1 U334 ( .A(n388), .B(n387), .ZN(n390) );
  NOR2_X1 U335 ( .A1(n523), .A2(n477), .ZN(n575) );
  XNOR2_X1 U336 ( .A(n462), .B(n461), .ZN(n511) );
  INV_X1 U337 ( .A(G190GAT), .ZN(n482) );
  INV_X1 U338 ( .A(G29GAT), .ZN(n485) );
  XNOR2_X1 U339 ( .A(n482), .B(KEYINPUT58), .ZN(n483) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n459) );
  XNOR2_X1 U341 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n460), .B(n459), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(n361), .B(G92GAT), .Z(n289) );
  XOR2_X1 U344 ( .A(KEYINPUT72), .B(G148GAT), .Z(n413) );
  XNOR2_X1 U345 ( .A(G204GAT), .B(n413), .ZN(n288) );
  XNOR2_X1 U346 ( .A(n289), .B(n288), .ZN(n295) );
  XOR2_X1 U347 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n291) );
  XNOR2_X1 U348 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n290) );
  XOR2_X1 U349 ( .A(n291), .B(n290), .Z(n293) );
  NAND2_X1 U350 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  INV_X1 U351 ( .A(n298), .ZN(n296) );
  NAND2_X1 U352 ( .A1(n296), .A2(KEYINPUT71), .ZN(n300) );
  INV_X1 U353 ( .A(KEYINPUT71), .ZN(n297) );
  NAND2_X1 U354 ( .A1(n298), .A2(n297), .ZN(n299) );
  NAND2_X1 U355 ( .A1(n300), .A2(n299), .ZN(n303) );
  XNOR2_X1 U356 ( .A(G99GAT), .B(G106GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n301), .B(G85GAT), .ZN(n348) );
  XNOR2_X1 U358 ( .A(n348), .B(KEYINPUT33), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U360 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n305) );
  XNOR2_X1 U361 ( .A(G71GAT), .B(G78GAT), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U363 ( .A(G57GAT), .B(n306), .ZN(n437) );
  XNOR2_X1 U364 ( .A(n307), .B(n437), .ZN(n462) );
  XOR2_X1 U365 ( .A(G1GAT), .B(KEYINPUT68), .Z(n438) );
  XOR2_X1 U366 ( .A(G141GAT), .B(G197GAT), .Z(n309) );
  XNOR2_X1 U367 ( .A(G50GAT), .B(G36GAT), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U369 ( .A(n438), .B(n310), .Z(n312) );
  NAND2_X1 U370 ( .A1(G229GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U372 ( .A(n313), .B(G8GAT), .Z(n320) );
  INV_X1 U373 ( .A(G43GAT), .ZN(n314) );
  NAND2_X1 U374 ( .A1(G29GAT), .A2(n314), .ZN(n316) );
  NAND2_X1 U375 ( .A1(n485), .A2(G43GAT), .ZN(n315) );
  NAND2_X1 U376 ( .A1(n316), .A2(n315), .ZN(n318) );
  XNOR2_X1 U377 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n331) );
  XNOR2_X1 U379 ( .A(n331), .B(KEYINPUT69), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U381 ( .A(G113GAT), .B(G15GAT), .Z(n322) );
  XNOR2_X1 U382 ( .A(G169GAT), .B(G22GAT), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U384 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n324) );
  XNOR2_X1 U385 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U387 ( .A(n326), .B(n325), .Z(n327) );
  XNOR2_X1 U388 ( .A(n328), .B(n327), .ZN(n576) );
  INV_X1 U389 ( .A(n576), .ZN(n539) );
  NAND2_X1 U390 ( .A1(n462), .A2(n539), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n329), .B(KEYINPUT74), .ZN(n494) );
  INV_X1 U392 ( .A(KEYINPUT9), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n332) );
  NAND2_X1 U394 ( .A1(G232GAT), .A2(G233GAT), .ZN(n333) );
  NAND2_X1 U395 ( .A1(n332), .A2(n333), .ZN(n337) );
  INV_X1 U396 ( .A(n332), .ZN(n335) );
  INV_X1 U397 ( .A(n333), .ZN(n334) );
  NAND2_X1 U398 ( .A1(n335), .A2(n334), .ZN(n336) );
  NAND2_X1 U399 ( .A1(n337), .A2(n336), .ZN(n339) );
  INV_X1 U400 ( .A(KEYINPUT76), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U402 ( .A(G50GAT), .B(G162GAT), .Z(n417) );
  XNOR2_X1 U403 ( .A(n417), .B(KEYINPUT77), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U405 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n343) );
  XNOR2_X1 U406 ( .A(G134GAT), .B(KEYINPUT75), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U408 ( .A(n345), .B(n344), .Z(n350) );
  XOR2_X1 U409 ( .A(G92GAT), .B(G218GAT), .Z(n347) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(G190GAT), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n348), .B(n358), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n559) );
  XNOR2_X1 U414 ( .A(n559), .B(KEYINPUT78), .ZN(n547) );
  XNOR2_X1 U415 ( .A(KEYINPUT36), .B(n547), .ZN(n587) );
  XNOR2_X1 U416 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n351), .B(G204GAT), .ZN(n421) );
  XOR2_X1 U418 ( .A(KEYINPUT79), .B(G211GAT), .Z(n353) );
  XNOR2_X1 U419 ( .A(G8GAT), .B(G183GAT), .ZN(n352) );
  XNOR2_X1 U420 ( .A(n353), .B(n352), .ZN(n441) );
  XNOR2_X1 U421 ( .A(n421), .B(n441), .ZN(n365) );
  XOR2_X1 U422 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n355) );
  XNOR2_X1 U423 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n354) );
  XNOR2_X1 U424 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U425 ( .A(G169GAT), .B(n356), .Z(n404) );
  XOR2_X1 U426 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n357) );
  XOR2_X1 U427 ( .A(n361), .B(n360), .Z(n363) );
  NAND2_X1 U428 ( .A1(G226GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n526), .B(KEYINPUT27), .ZN(n431) );
  XOR2_X1 U431 ( .A(KEYINPUT81), .B(G134GAT), .Z(n367) );
  XNOR2_X1 U432 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n366) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U434 ( .A(G113GAT), .B(n368), .ZN(n405) );
  XOR2_X1 U435 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n373) );
  XNOR2_X1 U436 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n287), .B(n369), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n370), .B(G141GAT), .ZN(n424) );
  INV_X1 U439 ( .A(n424), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n371), .B(KEYINPUT94), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U442 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n375) );
  XNOR2_X1 U443 ( .A(KEYINPUT6), .B(G57GAT), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U445 ( .A(n377), .B(n376), .Z(n388) );
  XOR2_X1 U446 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n379) );
  XNOR2_X1 U447 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U449 ( .A(G1GAT), .B(n380), .ZN(n386) );
  XOR2_X1 U450 ( .A(G155GAT), .B(G148GAT), .Z(n382) );
  XNOR2_X1 U451 ( .A(G127GAT), .B(G162GAT), .ZN(n381) );
  XNOR2_X1 U452 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U453 ( .A(G29GAT), .B(G85GAT), .Z(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n385) );
  NAND2_X1 U455 ( .A1(G225GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U456 ( .A(n390), .B(n389), .ZN(n391) );
  NAND2_X1 U457 ( .A1(n431), .A2(n523), .ZN(n535) );
  XOR2_X1 U458 ( .A(KEYINPUT82), .B(G190GAT), .Z(n393) );
  XNOR2_X1 U459 ( .A(G43GAT), .B(G99GAT), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U461 ( .A(G176GAT), .B(G183GAT), .Z(n395) );
  XNOR2_X1 U462 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U464 ( .A(n397), .B(n396), .Z(n402) );
  XOR2_X1 U465 ( .A(G15GAT), .B(G127GAT), .Z(n444) );
  XOR2_X1 U466 ( .A(n444), .B(KEYINPUT85), .Z(n399) );
  NAND2_X1 U467 ( .A1(G227GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U468 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U469 ( .A(G71GAT), .B(n400), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U471 ( .A(n404), .B(n403), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n406), .B(n405), .ZN(n562) );
  XOR2_X1 U473 ( .A(KEYINPUT87), .B(KEYINPUT90), .Z(n408) );
  XNOR2_X1 U474 ( .A(G218GAT), .B(G106GAT), .ZN(n407) );
  XNOR2_X1 U475 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U476 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n410) );
  XNOR2_X1 U477 ( .A(KEYINPUT22), .B(KEYINPUT86), .ZN(n409) );
  XNOR2_X1 U478 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U479 ( .A(n412), .B(n411), .Z(n419) );
  XOR2_X1 U480 ( .A(G22GAT), .B(G155GAT), .Z(n443) );
  XOR2_X1 U481 ( .A(n413), .B(n443), .Z(n415) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U486 ( .A(n420), .B(G78GAT), .Z(n423) );
  XNOR2_X1 U487 ( .A(n421), .B(G211GAT), .ZN(n422) );
  XNOR2_X1 U488 ( .A(n423), .B(n422), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n478) );
  XNOR2_X1 U490 ( .A(n478), .B(KEYINPUT28), .ZN(n503) );
  NAND2_X1 U491 ( .A1(n426), .A2(n503), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n427), .B(KEYINPUT99), .ZN(n436) );
  NAND2_X1 U493 ( .A1(n562), .A2(n526), .ZN(n428) );
  NAND2_X1 U494 ( .A1(n478), .A2(n428), .ZN(n429) );
  XNOR2_X1 U495 ( .A(n429), .B(KEYINPUT25), .ZN(n433) );
  NOR2_X1 U496 ( .A1(n478), .A2(n562), .ZN(n430) );
  XNOR2_X1 U497 ( .A(KEYINPUT26), .B(n430), .ZN(n574) );
  AND2_X1 U498 ( .A1(n431), .A2(n574), .ZN(n432) );
  NOR2_X1 U499 ( .A1(n433), .A2(n432), .ZN(n434) );
  NOR2_X1 U500 ( .A1(n523), .A2(n434), .ZN(n435) );
  XOR2_X1 U501 ( .A(KEYINPUT12), .B(G64GAT), .Z(n440) );
  XOR2_X1 U502 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U504 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U505 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U506 ( .A(n446), .B(n445), .ZN(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n448) );
  NAND2_X1 U508 ( .A1(G231GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U510 ( .A(KEYINPUT14), .B(n449), .Z(n450) );
  XNOR2_X1 U511 ( .A(n451), .B(n450), .ZN(n489) );
  NOR2_X1 U512 ( .A1(n492), .A2(n489), .ZN(n452) );
  XOR2_X1 U513 ( .A(KEYINPUT106), .B(n452), .Z(n453) );
  XOR2_X1 U514 ( .A(KEYINPUT108), .B(KEYINPUT37), .Z(n454) );
  XNOR2_X1 U515 ( .A(KEYINPUT107), .B(n454), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n456), .B(n455), .ZN(n522) );
  NOR2_X1 U517 ( .A1(n494), .A2(n522), .ZN(n458) );
  XOR2_X1 U518 ( .A(KEYINPUT38), .B(KEYINPUT109), .Z(n457) );
  XNOR2_X1 U519 ( .A(n458), .B(n457), .ZN(n509) );
  NAND2_X1 U520 ( .A1(n509), .A2(n562), .ZN(n460) );
  XOR2_X1 U521 ( .A(KEYINPUT117), .B(KEYINPUT47), .Z(n467) );
  NOR2_X1 U522 ( .A1(n511), .A2(n576), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n463), .B(KEYINPUT46), .ZN(n464) );
  XNOR2_X1 U524 ( .A(KEYINPUT116), .B(n489), .ZN(n570) );
  NOR2_X1 U525 ( .A1(n464), .A2(n570), .ZN(n465) );
  NAND2_X1 U526 ( .A1(n465), .A2(n559), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n467), .B(n466), .ZN(n472) );
  INV_X1 U528 ( .A(n489), .ZN(n584) );
  NOR2_X1 U529 ( .A1(n584), .A2(n587), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT45), .B(n468), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n469), .A2(n462), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n539), .A2(n470), .ZN(n471) );
  NOR2_X1 U533 ( .A1(n472), .A2(n471), .ZN(n474) );
  XOR2_X1 U534 ( .A(n526), .B(KEYINPUT120), .Z(n475) );
  NOR2_X1 U535 ( .A1(n536), .A2(n475), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT54), .B(n476), .Z(n477) );
  NAND2_X1 U537 ( .A1(n575), .A2(n478), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(n563) );
  INV_X1 U540 ( .A(n562), .ZN(n481) );
  AND2_X1 U541 ( .A1(n563), .A2(n286), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n523), .A2(n509), .ZN(n488) );
  XOR2_X1 U543 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n486) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n497) );
  NAND2_X1 U547 ( .A1(n489), .A2(n547), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT16), .B(n490), .ZN(n491) );
  NOR2_X1 U549 ( .A1(n492), .A2(n491), .ZN(n493) );
  XOR2_X1 U550 ( .A(KEYINPUT100), .B(n493), .Z(n512) );
  NOR2_X1 U551 ( .A1(n494), .A2(n512), .ZN(n495) );
  XOR2_X1 U552 ( .A(KEYINPUT101), .B(n495), .Z(n504) );
  NAND2_X1 U553 ( .A1(n504), .A2(n523), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U555 ( .A(G1GAT), .B(n498), .Z(G1324GAT) );
  NAND2_X1 U556 ( .A1(n526), .A2(n504), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n499), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n501) );
  NAND2_X1 U559 ( .A1(n504), .A2(n562), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U561 ( .A(G15GAT), .B(n502), .Z(G1326GAT) );
  INV_X1 U562 ( .A(n503), .ZN(n538) );
  NAND2_X1 U563 ( .A1(n504), .A2(n538), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n505), .B(KEYINPUT104), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G22GAT), .B(n506), .ZN(G1327GAT) );
  NAND2_X1 U566 ( .A1(n509), .A2(n526), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n507), .B(KEYINPUT110), .ZN(n508) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(n508), .ZN(G1329GAT) );
  NAND2_X1 U569 ( .A1(n538), .A2(n509), .ZN(n510) );
  XNOR2_X1 U570 ( .A(G50GAT), .B(n510), .ZN(G1331GAT) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n514) );
  INV_X1 U572 ( .A(n511), .ZN(n541) );
  NAND2_X1 U573 ( .A1(n576), .A2(n541), .ZN(n521) );
  NOR2_X1 U574 ( .A1(n512), .A2(n521), .ZN(n518) );
  NAND2_X1 U575 ( .A1(n523), .A2(n518), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  NAND2_X1 U577 ( .A1(n526), .A2(n518), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U579 ( .A(G71GAT), .B(KEYINPUT111), .Z(n517) );
  NAND2_X1 U580 ( .A1(n518), .A2(n562), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U583 ( .A1(n518), .A2(n538), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n525) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n531) );
  NAND2_X1 U587 ( .A1(n523), .A2(n531), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  XOR2_X1 U589 ( .A(G92GAT), .B(KEYINPUT113), .Z(n528) );
  NAND2_X1 U590 ( .A1(n531), .A2(n526), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n562), .A2(n531), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(KEYINPUT114), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n530), .ZN(G1338GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT44), .Z(n533) );
  NAND2_X1 U596 ( .A1(n531), .A2(n538), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n552) );
  NAND2_X1 U600 ( .A1(n552), .A2(n562), .ZN(n537) );
  NOR2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n539), .A2(n549), .ZN(n540) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U605 ( .A1(n549), .A2(n541), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n545) );
  NAND2_X1 U608 ( .A1(n549), .A2(n570), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U610 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  INV_X1 U612 ( .A(n547), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n552), .A2(n574), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n576), .A2(n558), .ZN(n553) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  NOR2_X1 U618 ( .A1(n511), .A2(n558), .ZN(n555) );
  XNOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n584), .A2(n558), .ZN(n557) );
  XOR2_X1 U623 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n569) );
  NOR2_X1 U628 ( .A1(n576), .A2(n569), .ZN(n564) );
  XOR2_X1 U629 ( .A(G169GAT), .B(n564), .Z(G1348GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n566) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n568) );
  NOR2_X1 U633 ( .A1(n511), .A2(n569), .ZN(n567) );
  XOR2_X1 U634 ( .A(n568), .B(n567), .Z(G1349GAT) );
  XOR2_X1 U635 ( .A(G183GAT), .B(KEYINPUT123), .Z(n573) );
  INV_X1 U636 ( .A(n569), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1350GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n576), .A2(n586), .ZN(n580) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(KEYINPUT60), .ZN(n578) );
  XNOR2_X1 U643 ( .A(KEYINPUT124), .B(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n462), .A2(n586), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n586), .ZN(n585) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n585), .Z(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(G218GAT), .B(n590), .Z(G1355GAT) );
endmodule

