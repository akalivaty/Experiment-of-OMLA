//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G116), .A2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT65), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n222), .B(new_n223), .C1(new_n219), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(KEYINPUT87), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT25), .ZN(new_n247));
  AOI211_X1 g0047(.A(G107), .B(new_n246), .C1(KEYINPUT86), .C2(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(KEYINPUT86), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n248), .A2(new_n249), .ZN(new_n252));
  INV_X1    g0052(.A(G107), .ZN(new_n253));
  INV_X1    g0053(.A(new_n246), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n212), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n203), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n251), .A2(new_n252), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n204), .B(G87), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT22), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT22), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(new_n204), .A4(G87), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT69), .B(G107), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT23), .B1(new_n273), .B2(new_n204), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n204), .A2(KEYINPUT23), .A3(G107), .ZN(new_n275));
  INV_X1    g0075(.A(G116), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT80), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT80), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G116), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n266), .A2(G20), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g0082(.A(KEYINPUT85), .B(KEYINPUT24), .Z(new_n283));
  NAND4_X1  g0083(.A1(new_n272), .A2(new_n274), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n284), .A2(new_n256), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n272), .A2(new_n274), .A3(new_n282), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n260), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n269), .A2(G257), .A3(G1698), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n269), .A2(G250), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G294), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT5), .B(G41), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n203), .A2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n212), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G41), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n297), .A2(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G264), .ZN(new_n303));
  OR2_X1    g0103(.A1(KEYINPUT5), .A2(G41), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT5), .A2(G41), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n298), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G274), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n300), .B2(new_n301), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n296), .A2(new_n303), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n294), .A2(new_n295), .B1(G264), .B2(new_n302), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(new_n309), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n245), .B1(new_n289), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n252), .ZN(new_n318));
  INV_X1    g0118(.A(new_n259), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n318), .A2(new_n250), .B1(new_n319), .B2(G107), .ZN(new_n320));
  INV_X1    g0120(.A(new_n288), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n284), .A2(new_n256), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n323), .A2(KEYINPUT87), .A3(new_n315), .A4(new_n312), .ZN(new_n324));
  INV_X1    g0124(.A(new_n310), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G190), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n310), .A2(G200), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n289), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n317), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT88), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT88), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n317), .A2(new_n324), .A3(new_n328), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  INV_X1    g0134(.A(G68), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT7), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n269), .B2(G20), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n261), .A2(new_n262), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n335), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G58), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n335), .ZN(new_n342));
  NOR2_X1   g0142(.A1(G58), .A2(G68), .ZN(new_n343));
  OAI21_X1  g0143(.A(G20), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(G20), .A2(G33), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G159), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n334), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n256), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n261), .B2(new_n262), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n267), .A2(KEYINPUT74), .A3(new_n268), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(new_n204), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n336), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n339), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G68), .ZN(new_n356));
  INV_X1    g0156(.A(new_n347), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n356), .A2(KEYINPUT75), .A3(KEYINPUT16), .A4(new_n357), .ZN(new_n358));
  NOR4_X1   g0158(.A1(new_n261), .A2(new_n262), .A3(new_n336), .A4(G20), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n353), .B2(new_n336), .ZN(new_n360));
  OAI211_X1 g0160(.A(KEYINPUT16), .B(new_n357), .C1(new_n360), .C2(new_n335), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT75), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n349), .B1(new_n358), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT67), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n301), .A2(G1), .A3(G13), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n203), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G232), .ZN(new_n371));
  INV_X1    g0171(.A(G226), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G1698), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G223), .B2(G1698), .ZN(new_n374));
  INV_X1    g0174(.A(G87), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n374), .A2(new_n338), .B1(new_n266), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n295), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n368), .A2(G274), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n365), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n371), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G190), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(G200), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT8), .B(G58), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT68), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n385), .B(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n246), .ZN(new_n389));
  INV_X1    g0189(.A(new_n256), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n203), .A2(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT17), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n383), .A2(new_n384), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT76), .B1(new_n364), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n349), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n361), .A2(new_n362), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n361), .A2(new_n362), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n383), .A2(new_n384), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT76), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n400), .A2(new_n402), .A3(new_n403), .A4(new_n394), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n389), .A2(new_n393), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n396), .A2(new_n404), .B1(new_n406), .B2(KEYINPUT17), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n381), .A2(new_n314), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n381), .A2(G169), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n405), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n410), .B1(new_n364), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT18), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n410), .C1(new_n364), .C2(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n407), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n379), .B1(new_n370), .B2(G238), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  OAI211_X1 g0219(.A(G232), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n420));
  OAI211_X1 g0220(.A(G226), .B(new_n291), .C1(new_n261), .C2(new_n262), .ZN(new_n421));
  INV_X1    g0221(.A(G97), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n420), .B(new_n421), .C1(new_n266), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n295), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n418), .A2(new_n419), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n419), .B1(new_n418), .B2(new_n424), .ZN(new_n426));
  OAI21_X1  g0226(.A(G169), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT14), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n418), .A2(new_n419), .A3(new_n424), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT73), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n418), .A2(new_n424), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT13), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n418), .A2(new_n424), .A3(KEYINPUT73), .A4(new_n419), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n431), .A2(new_n433), .A3(G179), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n436), .B(G169), .C1(new_n425), .C2(new_n426), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n428), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n281), .A2(G77), .B1(G20), .B2(new_n335), .ZN(new_n439));
  INV_X1    g0239(.A(G50), .ZN(new_n440));
  INV_X1    g0240(.A(new_n345), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n256), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT11), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n254), .A2(new_n335), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT12), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT71), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n257), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT71), .B1(new_n254), .B2(new_n256), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(G68), .A4(new_n391), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n442), .A2(KEYINPUT11), .A3(new_n256), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n445), .A2(new_n447), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n438), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n433), .A2(new_n429), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n455), .B2(G200), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n431), .A2(new_n433), .A3(G190), .A4(new_n434), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT10), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n338), .A2(new_n291), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G223), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n269), .A2(G222), .A3(new_n291), .ZN(new_n463));
  INV_X1    g0263(.A(new_n217), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n338), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n295), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n379), .B1(new_n370), .B2(G226), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(G190), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  INV_X1    g0270(.A(G200), .ZN(new_n471));
  OAI211_X1 g0271(.A(KEYINPUT72), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n387), .A2(new_n281), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n440), .A2(new_n341), .A3(new_n335), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n474), .A2(G20), .B1(G150), .B2(new_n345), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n390), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n254), .A2(new_n440), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n392), .B2(new_n440), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT9), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT9), .ZN(new_n480));
  INV_X1    g0280(.A(new_n478), .ZN(new_n481));
  INV_X1    g0281(.A(new_n475), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n387), .B2(new_n281), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n480), .B(new_n481), .C1(new_n483), .C2(new_n390), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n460), .B(new_n472), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n471), .B1(new_n467), .B2(new_n468), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(G190), .B2(new_n470), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n479), .A2(new_n484), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n489), .B(new_n490), .C1(KEYINPUT72), .C2(KEYINPUT10), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n461), .A2(G238), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n269), .A2(G232), .A3(new_n291), .ZN(new_n495));
  INV_X1    g0295(.A(new_n273), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n494), .B(new_n495), .C1(new_n269), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n295), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n379), .B1(new_n370), .B2(G244), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n311), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n385), .B(KEYINPUT70), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n441), .ZN(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT15), .B(G87), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n204), .A2(G33), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n204), .A2(new_n217), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n256), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n449), .A2(new_n450), .A3(G77), .A4(new_n391), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n217), .A2(new_n254), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n501), .B(new_n510), .C1(G179), .C2(new_n500), .ZN(new_n511));
  INV_X1    g0311(.A(new_n510), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n500), .B2(new_n382), .ZN(new_n513));
  INV_X1    g0313(.A(new_n500), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(new_n471), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n511), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n476), .A2(new_n478), .ZN(new_n517));
  INV_X1    g0317(.A(new_n470), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(new_n311), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n470), .A2(new_n314), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n417), .A2(new_n459), .A3(new_n493), .A4(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT4), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n338), .B2(new_n218), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n218), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n269), .A2(new_n291), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G283), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n269), .A2(G250), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n291), .B1(new_n532), .B2(KEYINPUT4), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n295), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n302), .A2(G257), .B1(new_n306), .B2(new_n308), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(G190), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT6), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n537), .A2(new_n422), .A3(G107), .ZN(new_n538));
  XNOR2_X1  g0338(.A(G97), .B(G107), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G77), .ZN(new_n541));
  OAI22_X1  g0341(.A1(new_n540), .A2(new_n204), .B1(new_n541), .B2(new_n441), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n496), .B1(new_n337), .B2(new_n339), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n256), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n246), .A2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n259), .B2(new_n422), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n536), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n302), .A2(G257), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n309), .ZN(new_n551));
  INV_X1    g0351(.A(G250), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n267), .B2(new_n268), .ZN(new_n553));
  OAI21_X1  g0353(.A(G1698), .B1(new_n553), .B2(new_n526), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n554), .A2(new_n529), .A3(new_n527), .A4(new_n530), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n555), .B2(new_n295), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n471), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT77), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n534), .A2(new_n535), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G200), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n441), .A2(new_n541), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n539), .A2(new_n537), .ZN(new_n562));
  INV_X1    g0362(.A(new_n538), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n561), .B1(new_n564), .B2(G20), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT7), .B1(new_n338), .B2(new_n204), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n273), .B1(new_n566), .B2(new_n359), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n390), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(new_n547), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT77), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n560), .A2(new_n569), .A3(new_n570), .A4(new_n536), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n558), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT78), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n559), .B2(G179), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n556), .A2(KEYINPUT78), .A3(new_n314), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n559), .A2(new_n311), .B1(new_n544), .B2(new_n548), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n204), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n375), .A2(new_n422), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n273), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n269), .A2(new_n204), .A3(G68), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n505), .B2(new_n422), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n256), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n504), .A2(new_n254), .ZN(new_n588));
  INV_X1    g0388(.A(new_n504), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n257), .A2(new_n258), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT81), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n586), .A2(new_n256), .B1(new_n254), .B2(new_n504), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT81), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(new_n590), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n269), .A2(G238), .A3(new_n291), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n269), .A2(G244), .A3(G1698), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n280), .A2(G33), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n295), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n295), .A2(new_n299), .A3(new_n552), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT79), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n378), .B2(new_n298), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n308), .A2(KEYINPUT79), .A3(new_n299), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n601), .A2(new_n606), .A3(new_n314), .ZN(new_n607));
  AOI21_X1  g0407(.A(G169), .B1(new_n601), .B2(new_n606), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n319), .A2(G87), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n593), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n471), .B1(new_n601), .B2(new_n606), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n601), .A2(new_n606), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G190), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n596), .A2(new_n609), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n572), .A2(new_n578), .A3(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n302), .A2(G270), .B1(new_n306), .B2(new_n308), .ZN(new_n619));
  OAI211_X1 g0419(.A(G264), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n620));
  OAI211_X1 g0420(.A(G257), .B(new_n291), .C1(new_n261), .C2(new_n262), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n267), .A2(G303), .A3(new_n268), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n295), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n619), .A2(KEYINPUT82), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT82), .B1(new_n619), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g0426(.A(G190), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n619), .A2(new_n624), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT82), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n619), .A2(new_n624), .A3(KEYINPUT82), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G200), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n277), .A2(new_n279), .A3(G20), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n530), .B(new_n204), .C1(G33), .C2(new_n422), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n256), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT20), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT20), .A4(new_n256), .ZN(new_n638));
  INV_X1    g0438(.A(new_n280), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n637), .A2(new_n638), .B1(new_n639), .B2(new_n254), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n449), .A2(new_n450), .A3(G116), .A4(new_n258), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n627), .A2(new_n632), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n311), .B1(new_n640), .B2(new_n641), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(KEYINPUT21), .A3(new_n630), .A4(new_n631), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT83), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n625), .A2(new_n626), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT83), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT21), .A4(new_n646), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n646), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT21), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n628), .A2(new_n314), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n653), .A2(new_n654), .B1(new_n642), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n645), .A2(new_n657), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n333), .A2(new_n525), .A3(new_n618), .A4(new_n658), .ZN(G372));
  INV_X1    g0459(.A(KEYINPUT89), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n492), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n487), .A2(KEYINPUT89), .A3(new_n491), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n511), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n458), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n407), .B1(new_n454), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(new_n416), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(new_n521), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n572), .A2(new_n328), .A3(new_n578), .A4(new_n617), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n289), .A2(new_n316), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n652), .A2(new_n656), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n596), .A2(new_n609), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n613), .A2(new_n616), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n674), .A2(new_n576), .A3(new_n675), .A4(new_n577), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI22_X1  g0478(.A1(new_n556), .A2(G169), .B1(new_n568), .B2(new_n547), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n574), .B2(new_n575), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT26), .B1(new_n680), .B2(new_n617), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n674), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n673), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n668), .B1(new_n524), .B2(new_n683), .ZN(G369));
  NAND3_X1  g0484(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(new_n687), .A3(G213), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n642), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT90), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n658), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n672), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n323), .A2(new_n690), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n333), .A2(new_n696), .B1(new_n670), .B2(new_n690), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n672), .A2(new_n690), .ZN(new_n700));
  INV_X1    g0500(.A(new_n690), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n333), .A2(new_n700), .B1(new_n670), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n207), .ZN(new_n704));
  OR3_X1    g0504(.A1(new_n704), .A2(KEYINPUT91), .A3(G41), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT91), .B1(new_n704), .B2(G41), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n273), .A2(G116), .A3(new_n581), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n210), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n701), .B1(new_n673), .B2(new_n682), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n317), .A2(new_n324), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n618), .B(new_n328), .C1(new_n714), .C2(new_n657), .ZN(new_n715));
  INV_X1    g0515(.A(new_n674), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n680), .A2(new_n617), .A3(KEYINPUT26), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n681), .B2(KEYINPUT92), .ZN(new_n718));
  OR3_X1    g0518(.A1(new_n676), .A2(KEYINPUT92), .A3(new_n677), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT93), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n715), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI211_X1 g0522(.A(KEYINPUT93), .B(new_n716), .C1(new_n718), .C2(new_n719), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n701), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n713), .B1(new_n724), .B2(KEYINPUT29), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n333), .A2(new_n618), .A3(new_n658), .A4(new_n701), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n615), .A2(new_n655), .A3(new_n556), .A4(new_n313), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n325), .A2(new_n615), .A3(G179), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n559), .A3(new_n649), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n727), .A2(new_n728), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n733), .B2(new_n690), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n726), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n725), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n711), .B1(new_n740), .B2(G1), .ZN(G364));
  INV_X1    g0541(.A(new_n707), .ZN(new_n742));
  INV_X1    g0542(.A(G13), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT94), .B1(new_n744), .B2(G45), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n203), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(KEYINPUT94), .A3(G45), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n742), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n694), .B2(G330), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G330), .B2(new_n694), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT95), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n704), .A2(new_n338), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G355), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G116), .B2(new_n207), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n351), .A2(new_n352), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n704), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G45), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(new_n760), .B2(new_n211), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n240), .A2(G45), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n756), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n212), .B1(G20), .B2(new_n311), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n749), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n471), .A2(G179), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(G20), .A3(G190), .ZN(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n338), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n204), .A2(new_n314), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n382), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n774), .B1(G326), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n382), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n204), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n776), .A2(G190), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G294), .A2(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n775), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n785), .A2(new_n382), .A3(G200), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n771), .A2(G20), .A3(new_n382), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n786), .A2(G322), .B1(G283), .B2(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n790));
  NOR4_X1   g0590(.A1(new_n204), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n790), .A2(G311), .B1(G329), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n778), .A2(new_n784), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n464), .A2(new_n790), .B1(new_n786), .B2(G58), .ZN(new_n794));
  INV_X1    g0594(.A(new_n782), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n335), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n780), .B(KEYINPUT98), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G97), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n800));
  INV_X1    g0600(.A(new_n791), .ZN(new_n801));
  INV_X1    g0601(.A(G159), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n801), .A2(new_n802), .A3(new_n800), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G50), .B2(new_n777), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n797), .A2(new_n799), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n787), .A2(new_n253), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n772), .A2(new_n375), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n807), .A2(new_n808), .A3(new_n338), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT97), .Z(new_n810));
  OAI21_X1  g0610(.A(new_n793), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT99), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n767), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n811), .B2(new_n812), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n770), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n766), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n694), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n753), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT100), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NOR2_X1   g0621(.A1(new_n511), .A2(new_n690), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n513), .A2(new_n515), .B1(new_n512), .B2(new_n701), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n511), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n712), .A2(new_n825), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n826), .A2(KEYINPUT102), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(KEYINPUT102), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n701), .B(new_n824), .C1(new_n673), .C2(new_n682), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n749), .B1(new_n830), .B2(new_n738), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n738), .B2(new_n830), .ZN(new_n832));
  INV_X1    g0632(.A(new_n749), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n767), .A2(new_n764), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n541), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G143), .A2(new_n786), .B1(new_n790), .B2(G159), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  INV_X1    g0637(.A(new_n777), .ZN(new_n838));
  INV_X1    g0638(.A(G150), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n836), .B1(new_n837), .B2(new_n838), .C1(new_n839), .C2(new_n795), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT34), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n757), .B1(new_n341), .B2(new_n780), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n801), .A2(new_n843), .B1(new_n440), .B2(new_n772), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n787), .A2(new_n335), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n280), .A2(new_n790), .B1(new_n782), .B2(G283), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n773), .B2(new_n838), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT101), .Z(new_n849));
  INV_X1    g0649(.A(G311), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n338), .B1(new_n801), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n772), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n786), .A2(G294), .B1(G107), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n375), .B2(new_n787), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n851), .B(new_n854), .C1(G97), .C2(new_n798), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n841), .A2(new_n846), .B1(new_n849), .B2(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n835), .B1(new_n814), .B2(new_n856), .C1(new_n824), .C2(new_n765), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n832), .A2(new_n857), .ZN(G384));
  NAND2_X1  g0658(.A1(new_n453), .A2(new_n690), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT106), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT106), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n453), .A2(new_n861), .A3(new_n690), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI221_X4 g0663(.A(new_n863), .B1(new_n457), .B2(new_n456), .C1(new_n438), .C2(new_n453), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n438), .A2(new_n453), .A3(new_n690), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n824), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n726), .B2(new_n736), .ZN(new_n867));
  INV_X1    g0667(.A(new_n688), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n364), .B2(new_n411), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n412), .A2(new_n406), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n357), .B1(new_n360), .B2(new_n335), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n390), .B1(new_n872), .B2(new_n334), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n398), .B2(new_n399), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n874), .A2(new_n405), .B1(new_n409), .B2(new_n408), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n688), .B1(new_n874), .B2(new_n405), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n364), .A2(new_n401), .A3(new_n411), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n871), .B1(new_n878), .B2(new_n870), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n876), .B1(new_n407), .B2(new_n416), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n867), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(KEYINPUT108), .B(KEYINPUT40), .Z(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT109), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT109), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(new_n869), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n407), .B2(new_n416), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n406), .A2(new_n412), .A3(new_n869), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n871), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n890), .B1(new_n896), .B2(KEYINPUT38), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(KEYINPUT40), .A3(new_n867), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n889), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n525), .A2(new_n737), .ZN(new_n901));
  OAI21_X1  g0701(.A(G330), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n901), .B2(new_n900), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n892), .B2(new_n895), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n881), .A2(new_n904), .A3(KEYINPUT39), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  AND4_X1   g0707(.A1(new_n870), .A2(new_n406), .A3(new_n412), .A4(new_n869), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n875), .A2(new_n877), .ZN(new_n909));
  INV_X1    g0709(.A(new_n876), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(new_n911), .B2(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n400), .A2(new_n405), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n414), .B1(new_n913), .B2(new_n410), .ZN(new_n914));
  INV_X1    g0714(.A(new_n415), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n404), .A2(new_n396), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n406), .A2(KEYINPUT17), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n910), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n907), .B1(new_n912), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n906), .B1(new_n921), .B2(new_n890), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT107), .B1(new_n905), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n454), .A2(new_n690), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT39), .B1(new_n881), .B2(new_n882), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n890), .B(new_n906), .C1(new_n896), .C2(KEYINPUT38), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT107), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n923), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n864), .A2(new_n865), .ZN(new_n930));
  INV_X1    g0730(.A(new_n822), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n829), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT105), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n829), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n930), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n921), .A2(new_n890), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n936), .A2(new_n937), .B1(new_n416), .B2(new_n688), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n929), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT29), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT92), .B1(new_n676), .B2(new_n677), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n678), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n676), .A2(KEYINPUT92), .A3(new_n677), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n674), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT93), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n720), .A2(new_n721), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(new_n715), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n940), .B1(new_n947), .B2(new_n701), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n525), .B1(new_n948), .B2(new_n713), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n668), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n939), .B(new_n950), .Z(new_n951));
  OR2_X1    g0751(.A1(new_n903), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n903), .A2(new_n951), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(new_n203), .C2(new_n744), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n211), .B1(new_n341), .B2(new_n335), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n955), .A2(new_n217), .B1(G50), .B2(new_n335), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(G1), .A3(new_n743), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT104), .Z(new_n958));
  OR2_X1    g0758(.A1(new_n564), .A2(KEYINPUT35), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n564), .A2(KEYINPUT35), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n959), .A2(G116), .A3(new_n213), .A4(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT36), .Z(new_n962));
  INV_X1    g0762(.A(KEYINPUT103), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n958), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n963), .B2(new_n962), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n954), .A2(new_n965), .ZN(G367));
  OAI211_X1 g0766(.A(new_n572), .B(new_n578), .C1(new_n569), .C2(new_n701), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n578), .B2(new_n701), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(new_n333), .A3(new_n700), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n970));
  INV_X1    g0770(.A(new_n714), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n578), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n969), .A2(KEYINPUT42), .B1(new_n701), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n611), .A2(new_n690), .ZN(new_n974));
  MUX2_X1   g0774(.A(new_n716), .B(new_n617), .S(new_n974), .Z(new_n975));
  AOI22_X1  g0775(.A1(new_n970), .A2(new_n973), .B1(KEYINPUT43), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n698), .A2(new_n968), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n707), .B(KEYINPUT41), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n702), .A2(new_n968), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n982), .A2(KEYINPUT111), .A3(KEYINPUT44), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(KEYINPUT44), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT110), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT111), .B1(new_n982), .B2(KEYINPUT44), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n982), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n983), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n702), .A2(new_n968), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT45), .Z(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n698), .ZN(new_n993));
  MUX2_X1   g0793(.A(new_n697), .B(new_n333), .S(new_n700), .Z(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(new_n695), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n739), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n989), .A2(new_n699), .A3(new_n991), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n993), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n981), .B1(new_n998), .B2(new_n740), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n748), .B(KEYINPUT112), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n980), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n768), .B1(new_n207), .B2(new_n504), .C1(new_n759), .C2(new_n236), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n749), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n269), .B1(new_n787), .B2(new_n217), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n786), .A2(G150), .B1(G137), .B2(new_n791), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n341), .B2(new_n772), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(G143), .C2(new_n777), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n790), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n1008), .A2(new_n440), .B1(new_n795), .B2(new_n802), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT113), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n798), .A2(G68), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1009), .A2(KEYINPUT113), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT46), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n772), .A2(new_n1014), .A3(new_n276), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G303), .B2(new_n786), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n757), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n791), .A2(G317), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n790), .A2(G283), .B1(G97), .B2(new_n788), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n273), .A2(new_n781), .B1(new_n777), .B2(G311), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1014), .B1(new_n639), .B2(new_n772), .ZN(new_n1022));
  INV_X1    g0822(.A(G294), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1021), .B(new_n1022), .C1(new_n1023), .C2(new_n795), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1013), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT47), .Z(new_n1026));
  OAI221_X1 g0826(.A(new_n1003), .B1(new_n817), .B2(new_n975), .C1(new_n1026), .C2(new_n814), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1001), .A2(new_n1027), .ZN(G387));
  INV_X1    g0828(.A(new_n708), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n754), .A2(new_n1029), .B1(new_n253), .B2(new_n704), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n502), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n440), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n760), .B1(new_n335), .B2(new_n541), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1033), .A2(new_n1029), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n233), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n758), .B1(new_n1036), .B2(new_n760), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1030), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n833), .B1(new_n1038), .B2(new_n768), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G303), .A2(new_n790), .B1(new_n786), .B2(G317), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n777), .A2(G322), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n850), .C2(new_n795), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n781), .A2(G283), .B1(new_n852), .B2(G294), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT49), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n639), .A2(new_n787), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n757), .B(new_n1049), .C1(G326), .C2(new_n791), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n798), .A2(new_n589), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G50), .A2(new_n786), .B1(new_n790), .B2(G68), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n852), .A2(new_n464), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n388), .C2(new_n795), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n788), .A2(G97), .B1(new_n791), .B2(G150), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1055), .B(new_n757), .C1(new_n802), .C2(new_n838), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1048), .A2(new_n1050), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1039), .B1(new_n1058), .B2(new_n814), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n697), .B2(new_n766), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n995), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n1000), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n740), .A2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n742), .B1(new_n739), .B2(new_n995), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(G393));
  AND2_X1   g0865(.A1(new_n998), .A2(new_n742), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n993), .A2(new_n997), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1066), .B1(new_n996), .B2(new_n1067), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n968), .A2(new_n817), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n768), .B1(new_n422), .B2(new_n207), .C1(new_n759), .C2(new_n243), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT114), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1072), .A2(new_n749), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(G283), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1008), .A2(new_n1023), .B1(new_n1075), .B2(new_n772), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G322), .B2(new_n791), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n269), .B(new_n807), .C1(G303), .C2(new_n782), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n639), .C2(new_n780), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n786), .A2(G311), .B1(new_n777), .B2(G317), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT52), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n798), .A2(G77), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n791), .A2(G143), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n375), .B2(new_n787), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G68), .B2(new_n852), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1031), .A2(new_n790), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1017), .B1(G50), .B2(new_n782), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1082), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n786), .A2(G159), .B1(new_n777), .B2(G150), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT51), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1079), .A2(new_n1081), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1074), .B1(new_n767), .B2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1067), .A2(new_n1000), .B1(new_n1069), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1068), .A2(new_n1093), .ZN(G390));
  AND2_X1   g0894(.A1(new_n737), .A2(G330), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n930), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n824), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n924), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n829), .A2(new_n934), .A3(new_n931), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n934), .B1(new_n829), .B2(new_n931), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n923), .A2(new_n928), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n897), .A2(new_n1098), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n823), .A2(new_n511), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n701), .B(new_n1104), .C1(new_n722), .C2(new_n723), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n931), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1103), .B1(new_n1106), .B2(new_n1096), .ZN(new_n1107));
  OAI211_X1 g0907(.A(KEYINPUT115), .B(new_n1097), .C1(new_n1102), .C2(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n927), .B1(new_n925), .B2(new_n926), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1109), .A2(new_n1110), .B1(new_n936), .B2(new_n924), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1106), .A2(new_n1096), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1103), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1097), .A2(KEYINPUT115), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1097), .A2(KEYINPUT115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1111), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1108), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n764), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n786), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1120), .A2(new_n276), .B1(new_n1023), .B2(new_n801), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n845), .B(new_n1121), .C1(G97), .C2(new_n790), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n777), .A2(G283), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n269), .B(new_n808), .C1(new_n273), .C2(new_n782), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1122), .A2(new_n1082), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n777), .A2(G128), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n269), .C1(new_n1127), .C2(new_n801), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G137), .B2(new_n782), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1008), .A2(new_n1130), .B1(new_n440), .B2(new_n787), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G132), .B2(new_n786), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n798), .A2(G159), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n772), .A2(new_n839), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n814), .B1(new_n1125), .B2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n833), .B(new_n1137), .C1(new_n388), .C2(new_n834), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1118), .A2(new_n1000), .B1(new_n1119), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1095), .A2(new_n525), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n668), .B(new_n1140), .C1(new_n725), .C2(new_n524), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT116), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n949), .A2(KEYINPUT116), .A3(new_n668), .A4(new_n1140), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1096), .B1(new_n1095), .B2(new_n824), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n738), .A2(new_n825), .A3(new_n930), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1145), .A2(new_n1146), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n930), .B1(new_n738), .B2(new_n825), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1097), .A2(new_n931), .A3(new_n1148), .A4(new_n1105), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1143), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1151), .A2(new_n1108), .A3(new_n1117), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1143), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n707), .B1(new_n1118), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT117), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AOI211_X1 g0956(.A(KEYINPUT117), .B(new_n707), .C1(new_n1118), .C2(new_n1153), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1139), .B1(new_n1156), .B2(new_n1157), .ZN(G378));
  INV_X1    g0958(.A(G41), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1017), .A2(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1120), .A2(new_n253), .B1(new_n341), .B2(new_n787), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(G283), .C2(new_n791), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1053), .B1(new_n838), .B2(new_n276), .C1(new_n504), .C2(new_n1008), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G97), .B2(new_n782), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1164), .A3(new_n1011), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT58), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G50), .B1(new_n266), .B2(new_n1159), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1165), .A2(new_n1166), .B1(new_n1160), .B2(new_n1167), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1008), .A2(new_n837), .B1(new_n772), .B2(new_n1130), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G128), .B2(new_n786), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n1127), .B2(new_n838), .C1(new_n843), .C2(new_n795), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G150), .B2(new_n798), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G33), .B(G41), .C1(new_n791), .C2(G124), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n802), .B2(new_n787), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1168), .B1(new_n1166), .B2(new_n1165), .C1(new_n1174), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n767), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n834), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1178), .B(new_n749), .C1(G50), .C2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1181));
  INV_X1    g0981(.A(KEYINPUT119), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n663), .B2(new_n521), .ZN(new_n1183));
  AOI211_X1 g0983(.A(KEYINPUT119), .B(new_n522), .C1(new_n661), .C2(new_n662), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1181), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n517), .A2(new_n688), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n662), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT89), .B1(new_n487), .B2(new_n491), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n521), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT119), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n663), .A2(new_n1182), .A3(new_n521), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1181), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1185), .A2(new_n1186), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1186), .B1(new_n1185), .B2(new_n1193), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1180), .B1(new_n1197), .B2(new_n764), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT120), .Z(new_n1199));
  NAND4_X1  g0999(.A1(new_n889), .A2(G330), .A3(new_n1196), .A4(new_n898), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n883), .A2(new_n887), .A3(new_n884), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n887), .B1(new_n883), .B2(new_n884), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n898), .B(G330), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1197), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n939), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT121), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1200), .B(new_n1204), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1204), .A2(new_n1200), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1206), .B1(new_n929), .B2(new_n938), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1199), .B1(new_n1211), .B2(new_n1000), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1118), .A2(new_n1153), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1204), .A2(new_n1200), .A3(new_n939), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n939), .B1(new_n1204), .B2(new_n1200), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT57), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT122), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1216), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1208), .A2(new_n1205), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1204), .A2(new_n1200), .A3(new_n939), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(KEYINPUT57), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1214), .B1(new_n1118), .B2(new_n1150), .ZN(new_n1226));
  OAI21_X1  g1026(.A(KEYINPUT122), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1222), .A2(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1213), .A2(new_n1215), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n742), .B1(new_n1229), .B2(KEYINPUT57), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1212), .B1(new_n1228), .B2(new_n1230), .ZN(G375));
  NAND3_X1  g1031(.A1(new_n1214), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n981), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1151), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n338), .B1(new_n801), .B2(new_n773), .C1(new_n795), .C2(new_n639), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n852), .A2(G97), .B1(new_n788), .B2(G77), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n1120), .B2(new_n1075), .C1(new_n496), .C2(new_n1008), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1235), .B(new_n1237), .C1(G294), .C2(new_n777), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n798), .A2(G50), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n757), .B1(new_n341), .B2(new_n787), .C1(new_n1008), .C2(new_n839), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n852), .A2(G159), .B1(G128), .B2(new_n791), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1120), .B2(new_n837), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n843), .A2(new_n838), .B1(new_n795), .B2(new_n1130), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1240), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1238), .A2(new_n1051), .B1(new_n1239), .B2(new_n1244), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n749), .B1(G68), .B2(new_n1179), .C1(new_n1245), .C2(new_n814), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n930), .B2(new_n764), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1150), .B2(new_n1000), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1234), .A2(new_n1248), .ZN(G381));
  OR4_X1    g1049(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1250), .A2(G387), .A3(G381), .ZN(new_n1251));
  INV_X1    g1051(.A(G378), .ZN(new_n1252));
  INV_X1    g1052(.A(G375), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(G407));
  NAND2_X1  g1054(.A1(new_n689), .A2(G213), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1252), .A3(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(G407), .A2(G213), .A3(new_n1257), .ZN(G409));
  XNOR2_X1  g1058(.A(new_n820), .B(G393), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G387), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT124), .B1(new_n1001), .B2(new_n1027), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G390), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1262), .B(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G378), .B(new_n1212), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1199), .B1(new_n1267), .B2(new_n1000), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1216), .A2(new_n1233), .A3(new_n1211), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1157), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1152), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1273), .A3(new_n1139), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1256), .B1(new_n1266), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1151), .A2(KEYINPUT60), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n742), .B1(new_n1276), .B2(new_n1232), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1276), .A2(new_n1232), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1248), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n832), .A3(new_n857), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G384), .B(new_n1248), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1275), .A2(KEYINPUT62), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT62), .B1(new_n1275), .B2(new_n1283), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1275), .A2(new_n1283), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1286), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1266), .A2(new_n1274), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1255), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1256), .A2(G2897), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1280), .A2(new_n1281), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1290), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1265), .B1(new_n1287), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1296), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1294), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1264), .B(new_n1301), .C1(new_n1303), .C2(new_n1275), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1275), .A2(KEYINPUT63), .A3(new_n1283), .ZN(new_n1306));
  AOI211_X1 g1106(.A(KEYINPUT123), .B(KEYINPUT63), .C1(new_n1275), .C2(new_n1283), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT123), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1288), .B2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1305), .B(new_n1306), .C1(new_n1307), .C2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1300), .A2(new_n1311), .ZN(G405));
  OAI21_X1  g1112(.A(new_n1282), .B1(new_n1253), .B2(G378), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1283), .A2(new_n1252), .A3(G375), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(KEYINPUT126), .A3(new_n1266), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1266), .A2(KEYINPUT126), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1313), .A2(new_n1317), .A3(new_n1314), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1316), .A2(new_n1318), .A3(new_n1265), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1265), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(G402));
endmodule


