//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT91), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G15gat), .ZN(new_n207));
  INV_X1    g006(.A(G15gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT90), .ZN(new_n213));
  INV_X1    g012(.A(G1gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n212), .A2(new_n213), .B1(KEYINPUT16), .B2(new_n214), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT90), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT90), .B1(new_n207), .B2(new_n209), .ZN(new_n217));
  NOR3_X1   g016(.A1(new_n216), .A2(new_n217), .A3(G1gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n204), .B(new_n205), .C1(new_n215), .C2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G43gat), .B(G50gat), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT14), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT14), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G29gat), .A2(G36gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT15), .B(new_n220), .C1(new_n226), .C2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n226), .B(KEYINPUT88), .ZN(new_n230));
  XOR2_X1   g029(.A(G43gat), .B(G50gat), .Z(new_n231));
  INV_X1    g030(.A(KEYINPUT15), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n227), .B(KEYINPUT89), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n229), .B1(new_n230), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n214), .A2(KEYINPUT16), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n216), .B2(new_n217), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n212), .A2(new_n214), .A3(new_n213), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n204), .A2(new_n205), .ZN(new_n241));
  NAND2_X1  g040(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n239), .A2(new_n240), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n219), .A2(new_n237), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n237), .B1(new_n219), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n203), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT92), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(KEYINPUT92), .B(new_n203), .C1(new_n244), .C2(new_n245), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n237), .A2(KEYINPUT17), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT17), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n229), .B(new_n252), .C1(new_n230), .C2(new_n236), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n219), .A2(new_n243), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n244), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n257), .A3(new_n202), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT18), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT18), .A4(new_n202), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n250), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G113gat), .B(G141gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(G197gat), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT11), .B(G169gat), .Z(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT12), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n250), .A2(new_n260), .A3(new_n267), .A4(new_n261), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT83), .ZN(new_n273));
  INV_X1    g072(.A(G127gat), .ZN(new_n274));
  INV_X1    g073(.A(G134gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G127gat), .A2(G134gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G113gat), .B(G120gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(KEYINPUT68), .A3(new_n277), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT69), .B(KEYINPUT1), .Z(new_n284));
  NAND4_X1  g083(.A1(new_n280), .A2(new_n282), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n276), .B(new_n277), .C1(new_n281), .C2(KEYINPUT1), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT70), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n289));
  NAND2_X1  g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT2), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT77), .ZN(new_n292));
  INV_X1    g091(.A(G155gat), .ZN(new_n293));
  INV_X1    g092(.A(G162gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n290), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G141gat), .B(G148gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n299), .B1(G155gat), .B2(G162gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n292), .B(new_n296), .C1(new_n298), .C2(new_n300), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n305), .A3(new_n286), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n288), .A2(new_n289), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n286), .A3(new_n285), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT79), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT4), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n308), .B2(KEYINPUT4), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n304), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n302), .A2(KEYINPUT3), .A3(new_n303), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n287), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n273), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AOI211_X1 g119(.A(KEYINPUT83), .B(new_n318), .C1(new_n312), .C2(new_n316), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n304), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n287), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n308), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n322), .B(KEYINPUT39), .C1(new_n319), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n316), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n308), .A2(KEYINPUT4), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT79), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT4), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n327), .B1(new_n331), .B2(new_n307), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT83), .B1(new_n332), .B2(new_n318), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n273), .A3(new_n319), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT39), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(G1gat), .B(G29gat), .Z(new_n336));
  XNOR2_X1  g135(.A(G57gat), .B(G85gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT82), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n335), .A2(KEYINPUT84), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT84), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT39), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n320), .B2(new_n321), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(new_n346), .B2(new_n341), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n326), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(KEYINPUT40), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G226gat), .ZN(new_n352));
  INV_X1    g151(.A(G233gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(KEYINPUT26), .ZN(new_n358));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n359), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G183gat), .ZN(new_n362));
  INV_X1    g161(.A(G190gat), .ZN(new_n363));
  OAI22_X1  g162(.A1(new_n358), .A2(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(KEYINPUT27), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT27), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G183gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT67), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT67), .ZN(new_n370));
  AOI21_X1  g169(.A(G190gat), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT28), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n368), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(KEYINPUT28), .A3(new_n363), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n364), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n356), .A2(KEYINPUT23), .ZN(new_n378));
  NAND3_X1  g177(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT64), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n359), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT65), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT66), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT24), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(G183gat), .A3(G190gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(G183gat), .B(G190gat), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n384), .B(new_n386), .C1(new_n387), .C2(new_n385), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n385), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT66), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT25), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n357), .B2(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n383), .A2(new_n388), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n357), .A2(new_n392), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n359), .A3(new_n378), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n396), .B2(new_n389), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n377), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n355), .B1(new_n398), .B2(KEYINPUT29), .ZN(new_n399));
  XNOR2_X1  g198(.A(G211gat), .B(G218gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT22), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT72), .B(G211gat), .ZN(new_n403));
  INV_X1    g202(.A(G218gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT73), .ZN(new_n406));
  XNOR2_X1  g205(.A(G197gat), .B(G204gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n406), .B1(new_n405), .B2(new_n407), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n401), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n410), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(new_n408), .A3(new_n400), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n390), .A2(new_n388), .A3(new_n393), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT65), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n382), .B(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n397), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n374), .A2(new_n376), .ZN(new_n420));
  INV_X1    g219(.A(new_n364), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT74), .B1(new_n423), .B2(new_n354), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT74), .ZN(new_n425));
  AOI211_X1 g224(.A(new_n425), .B(new_n355), .C1(new_n419), .C2(new_n422), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n399), .B(new_n415), .C1(new_n424), .C2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n354), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n398), .A2(new_n355), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n414), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n431), .A3(KEYINPUT75), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n425), .B1(new_n398), .B2(new_n355), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n423), .A2(KEYINPUT74), .A3(new_n354), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT75), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n415), .ZN(new_n437));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT76), .ZN(new_n439));
  XNOR2_X1  g238(.A(G64gat), .B(G92gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  AND3_X1   g240(.A1(new_n432), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n432), .B2(new_n437), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(KEYINPUT30), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n432), .A2(new_n437), .ZN(new_n445));
  INV_X1    g244(.A(new_n441), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT5), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n316), .A2(new_n450), .A3(new_n318), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n312), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n450), .B1(new_n325), .B2(new_n319), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n288), .A2(KEYINPUT4), .A3(new_n304), .A4(new_n306), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n308), .A2(new_n289), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n455), .A2(new_n316), .A3(new_n456), .A4(new_n318), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n444), .A2(new_n449), .B1(new_n459), .B2(new_n342), .ZN(new_n460));
  OAI221_X1 g259(.A(new_n326), .B1(new_n349), .B2(KEYINPUT40), .C1(new_n343), .C2(new_n347), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n351), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G78gat), .B(G106gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(G22gat), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n411), .A2(new_n413), .A3(new_n428), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT3), .B1(new_n466), .B2(KEYINPUT80), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n411), .A2(new_n413), .A3(new_n468), .A4(new_n428), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n304), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n314), .A2(new_n428), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n414), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(G228gat), .B(G233gat), .C1(new_n470), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G228gat), .A2(G233gat), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n466), .A2(new_n313), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n475), .B(new_n472), .C1(new_n476), .C2(new_n304), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT31), .B(G50gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n479), .B1(new_n474), .B2(new_n477), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n465), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n474), .A2(new_n477), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n478), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n464), .A3(new_n480), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n340), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n459), .A2(KEYINPUT6), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT86), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n312), .A2(new_n452), .B1(new_n454), .B2(new_n457), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT6), .B1(new_n492), .B2(new_n340), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n459), .A2(new_n342), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n492), .A2(new_n340), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT6), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n447), .A2(new_n491), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT37), .B1(new_n432), .B2(new_n437), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n399), .B(new_n414), .C1(new_n424), .C2(new_n426), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n415), .B1(new_n429), .B2(new_n430), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT37), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT38), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n500), .A2(new_n505), .A3(new_n446), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT87), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n445), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n509), .A2(new_n504), .A3(new_n441), .A4(new_n503), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n495), .A2(new_n498), .A3(new_n491), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT87), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .A4(new_n447), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n509), .A2(new_n441), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n445), .A2(new_n508), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT38), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n507), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n462), .A2(new_n488), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n442), .ZN(new_n519));
  INV_X1    g318(.A(new_n493), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n490), .B1(new_n520), .B2(new_n496), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n443), .A2(KEYINPUT30), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n449), .A2(new_n519), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n487), .A2(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(G15gat), .B(G43gat), .Z(new_n525));
  XNOR2_X1  g324(.A(G71gat), .B(G99gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G227gat), .A2(G233gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n288), .A2(new_n306), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n423), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n419), .A2(new_n422), .A3(new_n288), .A4(new_n306), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n527), .B1(new_n532), .B2(KEYINPUT33), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT32), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n531), .ZN(new_n537));
  INV_X1    g336(.A(new_n528), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT71), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT34), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n533), .A2(new_n535), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT34), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT71), .B(new_n542), .C1(new_n537), .C2(new_n538), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n536), .A2(new_n540), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n543), .ZN(new_n545));
  AOI211_X1 g344(.A(new_n534), .B(new_n532), .C1(KEYINPUT33), .C2(new_n527), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n533), .A2(new_n535), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n544), .A2(new_n548), .A3(KEYINPUT36), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT36), .B1(new_n544), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n524), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT81), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT81), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n524), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n518), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n444), .A2(new_n449), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n544), .A2(new_n548), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n488), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n483), .A2(new_n559), .A3(new_n486), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT35), .B1(new_n562), .B2(new_n523), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n272), .B1(new_n556), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(G57gat), .A2(G64gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(G57gat), .A2(G64gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT93), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G71gat), .ZN(new_n575));
  INV_X1    g374(.A(G78gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT93), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n578), .A3(new_n566), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n571), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n568), .A2(KEYINPUT94), .ZN(new_n582));
  AND2_X1   g381(.A1(G57gat), .A2(G64gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(G57gat), .A2(G64gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT94), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n566), .A2(new_n587), .A3(new_n567), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n582), .A2(new_n585), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n581), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(new_n274), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n572), .A2(new_n573), .ZN(new_n600));
  XNOR2_X1  g399(.A(G57gat), .B(G64gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n602), .A2(KEYINPUT95), .A3(new_n582), .A4(new_n588), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n589), .A2(new_n590), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n599), .B1(new_n605), .B2(new_n581), .ZN(new_n606));
  AOI211_X1 g405(.A(KEYINPUT96), .B(new_n580), .C1(new_n603), .C2(new_n604), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n255), .B1(new_n609), .B2(new_n594), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n598), .B(new_n610), .Z(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n293), .ZN(new_n613));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n598), .B(new_n610), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622));
  XOR2_X1   g421(.A(G99gat), .B(G106gat), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n626), .A2(new_n627), .A3(G85gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT8), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT98), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n633));
  INV_X1    g432(.A(G85gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n625), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n636), .A3(new_n630), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G85gat), .A2(G92gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT7), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n624), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  AOI211_X1 g441(.A(new_n623), .B(new_n642), .C1(new_n632), .C2(new_n637), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n622), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n635), .A2(new_n636), .A3(new_n630), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n636), .B1(new_n635), .B2(new_n630), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n623), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n638), .A2(new_n624), .A3(new_n640), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT99), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n254), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n644), .A2(new_n237), .A3(new_n650), .ZN(new_n653));
  XNOR2_X1  g452(.A(G190gat), .B(G218gat), .ZN(new_n654));
  AND2_X1   g453(.A1(G232gat), .A2(G233gat), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n654), .A2(KEYINPUT100), .B1(KEYINPUT41), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n654), .A2(KEYINPUT100), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n652), .A2(new_n660), .A3(new_n653), .A4(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n655), .A2(KEYINPUT41), .ZN(new_n663));
  XNOR2_X1  g462(.A(G134gat), .B(G162gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n659), .A2(new_n665), .A3(new_n661), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n593), .B1(new_n641), .B2(new_n643), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n580), .B1(new_n603), .B2(new_n604), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n648), .A2(new_n649), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n593), .A2(KEYINPUT96), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n599), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(KEYINPUT10), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n675), .B1(new_n651), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(G230gat), .A2(G233gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT101), .ZN(new_n682));
  INV_X1    g481(.A(new_n680), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n650), .A4(new_n644), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(new_n675), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(G120gat), .B(G148gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(G176gat), .B(G204gat), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n671), .A2(new_n674), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n692), .B2(new_n683), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n682), .A2(new_n687), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n683), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n690), .B1(new_n681), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n621), .A2(new_n670), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n565), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n521), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n214), .ZN(G1324gat));
  NAND2_X1  g501(.A1(new_n556), .A2(new_n564), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n699), .A2(new_n557), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n271), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n565), .A2(KEYINPUT102), .A3(new_n704), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(G8gat), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT105), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n707), .A2(new_n711), .A3(G8gat), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT16), .B(G8gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT103), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n705), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(KEYINPUT104), .ZN(new_n718));
  INV_X1    g517(.A(new_n708), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT102), .B1(new_n565), .B2(new_n704), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n717), .B1(new_n721), .B2(new_n714), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n713), .A2(new_n722), .ZN(G1325gat));
  OAI21_X1  g522(.A(G15gat), .B1(new_n700), .B2(new_n551), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n559), .A2(new_n208), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n700), .B2(new_n725), .ZN(G1326gat));
  NOR2_X1   g525(.A1(new_n700), .A2(new_n488), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT43), .B(G22gat), .Z(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  AOI211_X1 g528(.A(KEYINPUT101), .B(new_n683), .C1(new_n684), .C2(new_n675), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n686), .B1(new_n679), .B2(new_n680), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n696), .B1(new_n732), .B2(new_n693), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n621), .A2(new_n670), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n565), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n521), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(new_n221), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n669), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n703), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n552), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n518), .A2(new_n744), .B1(new_n563), .B2(new_n561), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n745), .B2(new_n669), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n620), .A2(new_n272), .A3(new_n698), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G29gat), .B1(new_n749), .B2(new_n521), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n738), .A2(new_n739), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n740), .A2(new_n750), .A3(new_n751), .ZN(G1328gat));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n222), .A3(new_n557), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n754));
  OAI21_X1  g553(.A(G36gat), .B1(new_n749), .B2(new_n558), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(G1329gat));
  INV_X1    g556(.A(new_n551), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n746), .A3(new_n758), .A4(new_n748), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G43gat), .ZN(new_n760));
  INV_X1    g559(.A(G43gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n736), .A2(new_n761), .A3(new_n559), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n760), .A2(new_n762), .A3(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1330gat));
  NAND4_X1  g566(.A1(new_n743), .A2(new_n746), .A3(new_n487), .A4(new_n748), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G50gat), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n488), .A2(G50gat), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT106), .Z(new_n771));
  AND3_X1   g570(.A1(new_n565), .A2(new_n735), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n775));
  NOR2_X1   g574(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT108), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n777), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n772), .B1(new_n768), .B2(G50gat), .ZN(new_n780));
  INV_X1    g579(.A(new_n775), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(G1331gat));
  NAND4_X1  g582(.A1(new_n620), .A2(new_n272), .A3(new_n669), .A4(new_n698), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n745), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n737), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g586(.A1(new_n518), .A2(new_n744), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n564), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n790));
  INV_X1    g589(.A(new_n784), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT109), .B1(new_n745), .B2(new_n784), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n558), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT110), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n792), .A2(new_n793), .A3(new_n797), .A4(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n800));
  NOR2_X1   g599(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n796), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1333gat));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n785), .B2(new_n559), .ZN(new_n805));
  AND4_X1   g604(.A1(new_n804), .A2(new_n789), .A3(new_n559), .A4(new_n791), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n575), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n793), .ZN(new_n808));
  OAI21_X1  g607(.A(G71gat), .B1(new_n808), .B2(new_n551), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n807), .B2(new_n809), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(G1334gat));
  NOR2_X1   g612(.A1(new_n808), .A2(new_n488), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(new_n576), .ZN(G1335gat));
  NOR2_X1   g614(.A1(new_n620), .A2(new_n271), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n733), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n747), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G85gat), .B1(new_n819), .B2(new_n521), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n669), .B1(new_n788), .B2(new_n564), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT51), .B1(new_n821), .B2(new_n816), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n823));
  NOR4_X1   g622(.A1(new_n745), .A2(new_n823), .A3(new_n669), .A4(new_n817), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n521), .A2(new_n733), .A3(G85gat), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT112), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n820), .B1(new_n826), .B2(new_n828), .ZN(G1336gat));
  NAND4_X1  g628(.A1(new_n743), .A2(new_n746), .A3(new_n557), .A4(new_n818), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n633), .A2(new_n625), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n558), .A2(G92gat), .A3(new_n733), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n822), .B2(new_n824), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT114), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n832), .A2(new_n833), .A3(new_n835), .A4(new_n838), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1337gat));
  XNOR2_X1  g641(.A(KEYINPUT115), .B(G99gat), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n825), .A2(new_n559), .A3(new_n698), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n819), .A2(new_n551), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n843), .ZN(G1338gat));
  NAND4_X1  g645(.A1(new_n743), .A2(new_n746), .A3(new_n487), .A4(new_n818), .ZN(new_n847));
  XOR2_X1   g646(.A(KEYINPUT116), .B(G106gat), .Z(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n488), .A2(G106gat), .A3(new_n733), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n822), .B2(new_n824), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n851), .B(KEYINPUT117), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n825), .A2(new_n854), .B1(new_n847), .B2(new_n848), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n855), .B2(new_n850), .ZN(G1339gat));
  NAND4_X1  g655(.A1(new_n620), .A2(new_n272), .A3(new_n669), .A4(new_n733), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n675), .B(new_n683), .C1(new_n651), .C2(new_n678), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(KEYINPUT54), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n682), .A2(new_n859), .A3(new_n687), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n690), .B1(new_n685), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(KEYINPUT55), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n694), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n202), .B1(new_n256), .B2(new_n257), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n244), .A2(new_n245), .A3(new_n203), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n266), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n270), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n668), .A3(new_n667), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT55), .B1(new_n860), .B2(new_n862), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n864), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n270), .A2(new_n867), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n733), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n698), .A2(new_n868), .A3(KEYINPUT118), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n691), .B1(new_n681), .B2(KEYINPUT54), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(new_n732), .B2(new_n859), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n271), .B1(new_n877), .B2(KEYINPUT55), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n874), .B(new_n875), .C1(new_n878), .C2(new_n864), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n871), .B1(new_n879), .B2(new_n669), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n857), .B1(new_n880), .B2(new_n620), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NOR4_X1   g681(.A1(new_n882), .A2(new_n521), .A3(new_n562), .A4(new_n557), .ZN(new_n883));
  AOI21_X1  g682(.A(G113gat), .B1(new_n883), .B2(new_n271), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n558), .A2(new_n737), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n882), .A2(new_n562), .A3(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n271), .A2(G113gat), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(G1340gat));
  AOI21_X1  g687(.A(G120gat), .B1(new_n883), .B2(new_n698), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n698), .A2(G120gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n886), .B2(new_n890), .ZN(G1341gat));
  NAND3_X1  g690(.A1(new_n886), .A2(G127gat), .A3(new_n620), .ZN(new_n892));
  XOR2_X1   g691(.A(new_n892), .B(KEYINPUT119), .Z(new_n893));
  AOI21_X1  g692(.A(G127gat), .B1(new_n883), .B2(new_n620), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(G1342gat));
  NAND3_X1  g694(.A1(new_n883), .A2(new_n275), .A3(new_n670), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n886), .A2(new_n670), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n897), .B(new_n898), .C1(new_n275), .C2(new_n899), .ZN(G1343gat));
  NOR2_X1   g699(.A1(new_n758), .A2(new_n885), .ZN(new_n901));
  INV_X1    g700(.A(new_n857), .ZN(new_n902));
  INV_X1    g701(.A(new_n871), .ZN(new_n903));
  INV_X1    g702(.A(new_n864), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n272), .A2(new_n870), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n904), .A2(new_n905), .B1(new_n698), .B2(new_n868), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(new_n670), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n902), .B1(new_n907), .B2(new_n621), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(new_n909), .A3(new_n488), .ZN(new_n910));
  XNOR2_X1  g709(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n881), .B2(new_n487), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n901), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G141gat), .B1(new_n914), .B2(new_n272), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n758), .A2(new_n488), .A3(new_n557), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n881), .A2(new_n737), .A3(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(G141gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n271), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT58), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT58), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n915), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1344gat));
  NAND4_X1  g723(.A1(new_n881), .A2(new_n737), .A3(new_n698), .A4(new_n916), .ZN(new_n925));
  AOI21_X1  g724(.A(G148gat), .B1(new_n925), .B2(KEYINPUT59), .ZN(new_n926));
  INV_X1    g725(.A(new_n901), .ZN(new_n927));
  INV_X1    g726(.A(new_n913), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n907), .A2(new_n621), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT57), .B(new_n487), .C1(new_n929), .C2(new_n902), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n927), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n733), .A2(KEYINPUT59), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n881), .A2(new_n487), .A3(new_n912), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT121), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n909), .B1(new_n908), .B2(new_n488), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n881), .A2(new_n937), .A3(new_n487), .A4(new_n912), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n927), .A2(new_n733), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g740(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n933), .B(KEYINPUT122), .C1(new_n941), .C2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945));
  INV_X1    g744(.A(new_n932), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n925), .A2(KEYINPUT59), .ZN(new_n947));
  OAI22_X1  g746(.A1(new_n914), .A2(new_n946), .B1(G148gat), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n943), .B1(new_n939), .B2(new_n940), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n944), .A2(new_n950), .ZN(G1345gat));
  NAND3_X1  g750(.A1(new_n917), .A2(new_n293), .A3(new_n620), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n931), .A2(new_n620), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n954), .B2(new_n293), .ZN(G1346gat));
  NAND3_X1  g754(.A1(new_n917), .A2(new_n294), .A3(new_n670), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n931), .A2(new_n670), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n958), .B2(new_n294), .ZN(G1347gat));
  NAND2_X1  g758(.A1(new_n557), .A2(new_n521), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n960), .A2(new_n562), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n878), .A2(new_n864), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n874), .A2(new_n875), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n669), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n620), .B1(new_n964), .B2(new_n903), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n961), .B1(new_n965), .B2(new_n902), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(G169gat), .B1(new_n967), .B2(new_n271), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n881), .A2(new_n969), .A3(new_n961), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n881), .B2(new_n961), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n271), .A2(G169gat), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(G1348gat));
  NAND3_X1  g773(.A1(new_n972), .A2(G176gat), .A3(new_n698), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n977));
  AOI21_X1  g776(.A(G176gat), .B1(new_n967), .B2(new_n698), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(G1349gat));
  NAND3_X1  g778(.A1(new_n967), .A2(new_n375), .A3(new_n620), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n970), .A2(new_n971), .A3(new_n621), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n981), .B2(new_n362), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n363), .A3(new_n670), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n966), .A2(KEYINPUT123), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n881), .A2(new_n969), .A3(new_n961), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n985), .A2(new_n670), .A3(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n987), .A2(new_n988), .A3(G190gat), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n988), .B1(new_n987), .B2(G190gat), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT61), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n970), .A2(new_n971), .A3(new_n669), .ZN(new_n993));
  OAI21_X1  g792(.A(KEYINPUT125), .B1(new_n993), .B2(new_n363), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n987), .A2(new_n988), .A3(G190gat), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n984), .B1(new_n991), .B2(new_n996), .ZN(G1351gat));
  NOR2_X1   g796(.A1(new_n758), .A2(new_n960), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n881), .A2(new_n487), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g798(.A(G197gat), .B1(new_n999), .B2(new_n271), .ZN(new_n1000));
  AND2_X1   g799(.A1(new_n939), .A2(new_n998), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n271), .A2(G197gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(G1352gat));
  NAND2_X1  g802(.A1(new_n1001), .A2(new_n698), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(G204gat), .ZN(new_n1005));
  INV_X1    g804(.A(G204gat), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n999), .A2(new_n1006), .A3(new_n698), .ZN(new_n1007));
  XOR2_X1   g806(.A(new_n1007), .B(KEYINPUT62), .Z(new_n1008));
  NAND2_X1  g807(.A1(new_n1005), .A2(new_n1008), .ZN(G1353gat));
  NAND3_X1  g808(.A1(new_n999), .A2(new_n403), .A3(new_n620), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n939), .A2(new_n620), .A3(new_n998), .ZN(new_n1011));
  AND3_X1   g810(.A1(new_n1011), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1012));
  AOI21_X1  g811(.A(KEYINPUT63), .B1(new_n1011), .B2(G211gat), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(G1354gat));
  AOI21_X1  g813(.A(G218gat), .B1(new_n999), .B2(new_n670), .ZN(new_n1015));
  XNOR2_X1  g814(.A(new_n1015), .B(KEYINPUT126), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n670), .A2(G218gat), .ZN(new_n1017));
  XNOR2_X1  g816(.A(new_n1017), .B(KEYINPUT127), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n1016), .B1(new_n1001), .B2(new_n1018), .ZN(G1355gat));
endmodule


