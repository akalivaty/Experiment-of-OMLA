//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  NOR2_X1   g001(.A1(G29gat), .A2(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT14), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G29gat), .A2(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT89), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT88), .B1(new_n211), .B2(KEYINPUT15), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n211), .A2(KEYINPUT88), .A3(KEYINPUT15), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n205), .A2(new_n206), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT15), .A3(new_n211), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(G1gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G1gat), .B2(new_n219), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(G8gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n218), .B(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n226), .B2(new_n223), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n202), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n218), .B(new_n223), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n228), .B(KEYINPUT13), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n218), .B(KEYINPUT17), .ZN(new_n234));
  INV_X1    g033(.A(new_n223), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n224), .A4(new_n228), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n230), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT11), .B(G169gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G197gat), .ZN(new_n240));
  XOR2_X1   g039(.A(G113gat), .B(G141gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT12), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n230), .A2(new_n243), .A3(new_n233), .A4(new_n237), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G22gat), .B(G50gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G228gat), .ZN(new_n253));
  INV_X1    g052(.A(G233gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G155gat), .A2(G162gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT2), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT76), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G141gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G148gat), .ZN(new_n262));
  INV_X1    g061(.A(G148gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G141gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n257), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n260), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n257), .ZN(new_n268));
  NOR2_X1   g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT77), .B1(new_n263), .B2(G141gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT77), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(new_n261), .A3(G148gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n274), .A3(new_n264), .ZN(new_n275));
  INV_X1    g074(.A(new_n269), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(KEYINPUT78), .A3(new_n257), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT78), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n268), .B2(new_n269), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n275), .A2(new_n277), .A3(new_n279), .A4(new_n258), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n271), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT22), .B1(new_n284), .B2(G218gat), .ZN(new_n285));
  AND2_X1   g084(.A1(G211gat), .A2(G218gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(G211gat), .A2(G218gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g087(.A1(G197gat), .A2(G204gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(G197gat), .A2(G204gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n285), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n288), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT22), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT73), .B(G211gat), .ZN(new_n295));
  INV_X1    g094(.A(G218gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n291), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n293), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT74), .B1(new_n292), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n288), .B1(new_n285), .B2(new_n291), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT29), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n281), .B1(new_n304), .B2(KEYINPUT3), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n297), .A2(new_n293), .A3(new_n298), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n299), .A2(KEYINPUT74), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT75), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n300), .A2(new_n310), .A3(new_n303), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(new_n281), .B2(KEYINPUT3), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n256), .B1(new_n305), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT3), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n292), .A2(new_n299), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(KEYINPUT29), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n281), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n313), .A2(new_n300), .A3(new_n303), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n256), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n252), .B1(new_n315), .B2(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n271), .A2(new_n280), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n312), .B1(new_n307), .B2(new_n308), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(new_n316), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n255), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n321), .A3(new_n251), .ZN(new_n329));
  XOR2_X1   g128(.A(G78gat), .B(G106gat), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n323), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n331), .B1(new_n323), .B2(new_n329), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n250), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n323), .A2(new_n329), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n330), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n323), .A2(new_n329), .A3(new_n331), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n249), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n325), .A2(new_n316), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n341));
  INV_X1    g140(.A(G134gat), .ZN(new_n342));
  INV_X1    g141(.A(G120gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G113gat), .ZN(new_n344));
  INV_X1    g143(.A(G113gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G120gat), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT1), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G127gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G113gat), .B(G120gat), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n350), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n342), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n348), .ZN(new_n353));
  OAI21_X1  g152(.A(G127gat), .B1(new_n350), .B2(KEYINPUT1), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n354), .A3(G134gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT79), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(KEYINPUT80), .B(KEYINPUT4), .C1(new_n356), .C2(new_n281), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT4), .B1(new_n356), .B2(new_n281), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n325), .A2(new_n365), .A3(new_n355), .A4(new_n352), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n361), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n356), .B(new_n281), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n370), .B2(new_n359), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n373), .B(KEYINPUT4), .C1(new_n356), .C2(new_n281), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n363), .A2(KEYINPUT81), .A3(new_n366), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n361), .A2(new_n369), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT0), .B(G57gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(G85gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n372), .A2(new_n381), .A3(new_n376), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n377), .A2(KEYINPUT6), .A3(new_n382), .ZN(new_n387));
  INV_X1    g186(.A(G226gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(new_n254), .ZN(new_n389));
  NAND2_X1  g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT24), .ZN(new_n393));
  INV_X1    g192(.A(G183gat), .ZN(new_n394));
  INV_X1    g193(.A(G190gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT24), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n390), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n393), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(G169gat), .ZN(new_n400));
  INV_X1    g199(.A(G176gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT23), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n403), .A2(G169gat), .A3(G176gat), .ZN(new_n405));
  AND2_X1   g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT66), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT66), .ZN(new_n408));
  NAND2_X1  g207(.A1(G169gat), .A2(G176gat), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n408), .B(new_n409), .C1(new_n402), .C2(new_n403), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n399), .A2(new_n404), .A3(new_n407), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT25), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT26), .ZN(new_n413));
  NOR2_X1   g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n406), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n402), .A2(KEYINPUT26), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n415), .A2(new_n416), .B1(G183gat), .B2(G190gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n394), .A2(KEYINPUT27), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT68), .ZN(new_n419));
  AOI21_X1  g218(.A(G190gat), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT27), .B1(new_n394), .B2(KEYINPUT68), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT28), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT27), .B(G183gat), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n423), .A2(KEYINPUT28), .A3(new_n395), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n417), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n401), .A2(KEYINPUT23), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n400), .A2(KEYINPUT64), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT64), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G169gat), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n426), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n409), .B1(new_n414), .B2(KEYINPUT23), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT65), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n403), .A2(G176gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n428), .A2(G169gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n400), .A2(KEYINPUT64), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT65), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n406), .B1(new_n402), .B2(new_n403), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n390), .ZN(new_n441));
  NAND3_X1  g240(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT25), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n432), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n412), .A2(new_n425), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n389), .B1(new_n445), .B2(new_n312), .ZN(new_n446));
  INV_X1    g245(.A(new_n389), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n425), .A2(new_n444), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n448), .B2(new_n412), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n309), .B(new_n311), .C1(new_n446), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n312), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n447), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n300), .A2(new_n303), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n445), .A2(new_n389), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457));
  INV_X1    g256(.A(G64gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G92gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  OR3_X1    g260(.A1(new_n456), .A2(KEYINPUT30), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n456), .A2(new_n461), .ZN(new_n463));
  INV_X1    g262(.A(new_n461), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n450), .A2(new_n455), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(KEYINPUT30), .A3(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n386), .A2(new_n387), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n339), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT69), .B1(new_n445), .B2(new_n356), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n352), .A2(new_n355), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT69), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n448), .A2(new_n470), .A3(new_n471), .A4(new_n412), .ZN(new_n472));
  NAND2_X1  g271(.A1(G227gat), .A2(G233gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n445), .A2(new_n356), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n469), .A2(new_n472), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT34), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT32), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n478));
  INV_X1    g277(.A(new_n473), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT33), .B1(new_n478), .B2(new_n479), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G43gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(G71gat), .B(G99gat), .ZN(new_n483));
  XOR2_X1   g282(.A(new_n482), .B(new_n483), .Z(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n480), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  AOI221_X4 g285(.A(new_n477), .B1(KEYINPUT33), .B2(new_n484), .C1(new_n478), .C2(new_n479), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n476), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n478), .A2(new_n479), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT33), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n480), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n475), .B(KEYINPUT34), .Z(new_n494));
  INV_X1    g293(.A(new_n487), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT72), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n488), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(KEYINPUT72), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT36), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n486), .A2(KEYINPUT70), .A3(new_n487), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT70), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n493), .B2(new_n495), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n476), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT71), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT71), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n506), .B(new_n476), .C1(new_n501), .C2(new_n503), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n496), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n500), .B1(new_n508), .B2(KEYINPUT36), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n511));
  NAND3_X1  g310(.A1(new_n450), .A2(new_n455), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n450), .A2(new_n455), .A3(KEYINPUT86), .A4(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n452), .A2(new_n454), .A3(new_n309), .A4(new_n311), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n453), .B1(new_n446), .B2(new_n449), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(KEYINPUT37), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n461), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT38), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n465), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n464), .B1(new_n514), .B2(new_n515), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n456), .B2(KEYINPUT37), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n385), .A2(new_n384), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n381), .B1(new_n372), .B2(new_n376), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n387), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n526), .A2(new_n531), .B1(new_n338), .B2(new_n334), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT84), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n375), .A2(new_n357), .A3(new_n374), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n359), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n370), .A2(new_n359), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n535), .A2(KEYINPUT39), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT39), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n538), .A3(new_n359), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n381), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT83), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT83), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n542), .A3(new_n381), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n537), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n533), .B1(new_n544), .B2(KEYINPUT40), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n466), .A2(new_n462), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(new_n528), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(KEYINPUT40), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n535), .A2(KEYINPUT39), .A3(new_n536), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n539), .A2(new_n542), .A3(new_n381), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n542), .B1(new_n539), .B2(new_n381), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT40), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(KEYINPUT84), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n545), .A2(new_n547), .A3(new_n548), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n510), .B1(new_n532), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n465), .ZN(new_n557));
  AOI211_X1 g356(.A(KEYINPUT38), .B(new_n557), .C1(new_n523), .C2(new_n519), .ZN(new_n558));
  INV_X1    g357(.A(new_n525), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n531), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND4_X1   g359(.A1(new_n510), .A2(new_n560), .A3(new_n339), .A4(new_n555), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n468), .B(new_n509), .C1(new_n556), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n498), .A2(new_n499), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n339), .A3(new_n467), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n505), .A2(new_n496), .A3(new_n339), .A4(new_n507), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n467), .A2(KEYINPUT35), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n248), .B1(new_n562), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  INV_X1    g375(.A(G85gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(KEYINPUT8), .A2(new_n576), .B1(new_n577), .B2(new_n460), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT7), .ZN(new_n579));
  OAI22_X1  g378(.A1(new_n577), .A2(new_n460), .B1(new_n579), .B2(KEYINPUT92), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n581), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G99gat), .B(G106gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n218), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n575), .B(new_n586), .C1(new_n226), .C2(new_n585), .ZN(new_n587));
  XOR2_X1   g386(.A(G190gat), .B(G218gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT93), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n574), .B1(new_n590), .B2(KEYINPUT94), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n587), .B(new_n589), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G57gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n458), .ZN(new_n598));
  NAND2_X1  g397(.A1(G57gat), .A2(G64gat), .ZN(new_n599));
  AND2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(KEYINPUT9), .ZN(new_n601));
  NOR2_X1   g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n602), .A2(KEYINPUT90), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n600), .A2(new_n602), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n223), .B1(KEYINPUT21), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(new_n394), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT91), .Z(new_n612));
  OR2_X1    g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n612), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G211gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n615), .B(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n618), .B1(new_n613), .B2(new_n614), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n596), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n585), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(KEYINPUT95), .A3(KEYINPUT10), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n606), .A2(new_n585), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT10), .B1(new_n624), .B2(KEYINPUT95), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n627), .A2(KEYINPUT96), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT96), .B1(new_n627), .B2(new_n628), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n623), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n622), .B1(new_n626), .B2(new_n624), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G204gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT97), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n401), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n631), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n627), .A2(new_n628), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n622), .ZN(new_n640));
  INV_X1    g439(.A(new_n632), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n621), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n571), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n531), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g447(.A1(new_n645), .A2(new_n546), .ZN(new_n649));
  NAND2_X1  g448(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n650));
  INV_X1    g449(.A(G8gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n220), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n655), .B(new_n656), .C1(new_n651), .C2(new_n649), .ZN(G1325gat));
  AOI21_X1  g456(.A(G15gat), .B1(new_n646), .B2(new_n563), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT98), .ZN(new_n659));
  INV_X1    g458(.A(new_n509), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n660), .A2(G15gat), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n659), .B1(new_n646), .B2(new_n661), .ZN(G1326gat));
  NOR2_X1   g461(.A1(new_n645), .A2(new_n339), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT43), .B(G22gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  NOR2_X1   g464(.A1(new_n619), .A2(new_n620), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n638), .A2(new_n642), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n595), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n571), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n386), .A2(new_n387), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n673), .A2(G29gat), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT45), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n666), .B(KEYINPUT100), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n667), .B(KEYINPUT101), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n677), .A2(new_n248), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n596), .A2(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n569), .A2(KEYINPUT102), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n566), .B(new_n683), .C1(new_n567), .C2(new_n568), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n685), .A2(new_n686), .A3(new_n562), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n685), .B2(new_n562), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n681), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n562), .A2(new_n570), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n595), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT44), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n680), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n531), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G29gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n676), .A2(new_n695), .ZN(G1328gat));
  NOR3_X1   g495(.A1(new_n673), .A2(G36gat), .A3(new_n546), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT46), .ZN(new_n698));
  INV_X1    g497(.A(new_n546), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G36gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(G1329gat));
  INV_X1    g501(.A(new_n563), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n673), .A2(G43gat), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n693), .A2(new_n660), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(G43gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g506(.A(new_n339), .ZN(new_n708));
  INV_X1    g507(.A(new_n681), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n505), .A2(new_n507), .ZN(new_n710));
  INV_X1    g509(.A(new_n568), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n710), .A2(new_n496), .A3(new_n711), .A4(new_n339), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n683), .B1(new_n712), .B2(new_n566), .ZN(new_n713));
  INV_X1    g512(.A(new_n684), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n562), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT103), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n685), .A2(new_n686), .A3(new_n562), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n709), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n691), .A2(KEYINPUT44), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n708), .B(new_n679), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G50gat), .ZN(new_n721));
  INV_X1    g520(.A(G50gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n708), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT104), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n571), .A2(new_n670), .A3(new_n671), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT48), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(KEYINPUT105), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT48), .B1(new_n725), .B2(KEYINPUT105), .ZN(new_n729));
  AOI211_X1 g528(.A(new_n728), .B(new_n729), .C1(new_n720), .C2(G50gat), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT106), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n722), .B1(new_n693), .B2(new_n708), .ZN(new_n733));
  INV_X1    g532(.A(new_n725), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n736));
  INV_X1    g535(.A(new_n729), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n727), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n731), .A2(new_n739), .ZN(G1331gat));
  NOR2_X1   g539(.A1(new_n621), .A2(new_n247), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n678), .B(new_n741), .C1(new_n687), .C2(new_n688), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n674), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n597), .ZN(G1332gat));
  NOR2_X1   g543(.A1(new_n742), .A2(new_n546), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT49), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n458), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT107), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n745), .A2(new_n751), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n750), .A2(new_n746), .A3(new_n752), .A4(new_n458), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n742), .B2(new_n509), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n742), .A2(new_n703), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n758), .B2(G71gat), .ZN(new_n759));
  XOR2_X1   g558(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1334gat));
  NOR2_X1   g560(.A1(new_n742), .A2(new_n339), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT109), .B(G78gat), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1335gat));
  NAND2_X1  g563(.A1(new_n666), .A2(new_n248), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT110), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n715), .A2(new_n595), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(new_n643), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n577), .A3(new_n531), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n643), .B(new_n766), .C1(new_n718), .C2(new_n719), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n674), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1336gat));
  OAI21_X1  g573(.A(G92gat), .B1(new_n772), .B2(new_n546), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n769), .A2(new_n460), .A3(new_n699), .A4(new_n678), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g577(.A(G99gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n770), .A2(new_n779), .A3(new_n563), .ZN(new_n780));
  OAI21_X1  g579(.A(G99gat), .B1(new_n772), .B2(new_n509), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1338gat));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  INV_X1    g582(.A(G106gat), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n784), .A3(new_n708), .A4(new_n678), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G106gat), .B1(new_n772), .B2(new_n339), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n788), .B(new_n785), .C1(new_n786), .C2(new_n783), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1339gat));
  NOR3_X1   g591(.A1(new_n621), .A2(new_n247), .A3(new_n643), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n228), .B1(new_n236), .B2(new_n224), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n231), .A2(new_n232), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n242), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n246), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n667), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT54), .B1(new_n639), .B2(new_n622), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n631), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n803));
  NAND3_X1  g602(.A1(new_n639), .A2(new_n622), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n802), .A2(KEYINPUT55), .A3(new_n637), .A4(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n638), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n637), .B(new_n804), .C1(new_n631), .C2(new_n801), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n805), .A2(new_n247), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n800), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n596), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n805), .A2(new_n809), .ZN(new_n814));
  INV_X1    g613(.A(new_n798), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n814), .A2(new_n595), .A3(new_n806), .A4(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n794), .B1(new_n817), .B2(new_n677), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n674), .A2(new_n699), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n567), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n345), .A3(new_n247), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(new_n563), .A3(new_n339), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n248), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1340gat));
  INV_X1    g625(.A(new_n678), .ZN(new_n827));
  OAI21_X1  g626(.A(G120gat), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n643), .A2(new_n343), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n822), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n831), .ZN(G1341gat));
  INV_X1    g631(.A(new_n666), .ZN(new_n833));
  AOI21_X1  g632(.A(G127gat), .B1(new_n822), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n677), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n824), .A2(new_n348), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(G1342gat));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n342), .A3(new_n595), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT56), .Z(new_n839));
  OAI21_X1  g638(.A(G134gat), .B1(new_n824), .B2(new_n596), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1343gat));
  NAND2_X1  g640(.A1(new_n818), .A2(new_n708), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n509), .A2(new_n819), .ZN(new_n843));
  NOR4_X1   g642(.A1(new_n842), .A2(G141gat), .A3(new_n248), .A4(new_n843), .ZN(new_n844));
  XOR2_X1   g643(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n643), .A2(new_n848), .A3(new_n815), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT116), .B1(new_n667), .B2(new_n798), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n810), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n596), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n833), .B1(new_n852), .B2(new_n816), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n708), .B1(new_n853), .B2(new_n793), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n843), .B1(new_n847), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n247), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n844), .B1(new_n858), .B2(G141gat), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT58), .Z(G1344gat));
  NAND2_X1  g659(.A1(new_n854), .A2(new_n855), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT118), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n818), .A2(new_n708), .A3(new_n845), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n854), .A2(new_n864), .A3(new_n855), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n843), .B(KEYINPUT117), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n643), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n842), .A2(new_n843), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n263), .A3(new_n643), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n263), .B1(new_n857), .B2(new_n643), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n869), .B(new_n871), .C1(new_n872), .C2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g672(.A(G155gat), .B1(new_n870), .B2(new_n833), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n677), .A2(G155gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n857), .B2(new_n875), .ZN(G1346gat));
  AOI21_X1  g675(.A(G162gat), .B1(new_n870), .B2(new_n595), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n857), .A2(new_n595), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(G162gat), .ZN(G1347gat));
  AND2_X1   g678(.A1(new_n818), .A2(new_n674), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n880), .A2(new_n699), .A3(new_n821), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n881), .B(new_n247), .C1(new_n434), .C2(new_n435), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n674), .A2(new_n699), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT119), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n703), .A3(new_n708), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n818), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G169gat), .B1(new_n886), .B2(new_n248), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n882), .A2(new_n887), .ZN(G1348gat));
  NOR3_X1   g687(.A1(new_n886), .A2(new_n401), .A3(new_n827), .ZN(new_n889));
  AOI21_X1  g688(.A(G176gat), .B1(new_n881), .B2(new_n643), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n890), .A2(KEYINPUT120), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(KEYINPUT120), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(G1349gat));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(KEYINPUT60), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n894), .A2(KEYINPUT60), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n886), .A2(new_n835), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(G183gat), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n423), .A3(new_n833), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n895), .B(new_n896), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  AND4_X1   g701(.A1(new_n894), .A2(new_n900), .A3(new_n901), .A4(KEYINPUT60), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n886), .B2(new_n596), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT61), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n881), .A2(new_n395), .A3(new_n595), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1351gat));
  NOR2_X1   g707(.A1(new_n660), .A2(new_n884), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n909), .B(KEYINPUT124), .Z(new_n910));
  NAND3_X1  g709(.A1(new_n866), .A2(new_n247), .A3(new_n910), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT125), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(KEYINPUT125), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(G197gat), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n509), .A2(new_n699), .A3(new_n708), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT123), .Z(new_n916));
  AND2_X1   g715(.A1(new_n880), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(G197gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n247), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n914), .A2(new_n919), .ZN(G1352gat));
  XOR2_X1   g719(.A(KEYINPUT126), .B(G204gat), .Z(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n643), .A3(new_n922), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT62), .Z(new_n924));
  NAND2_X1  g723(.A1(new_n866), .A2(new_n910), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n925), .B2(new_n827), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1353gat));
  NAND3_X1  g726(.A1(new_n866), .A2(new_n833), .A3(new_n910), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT127), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n866), .A2(new_n930), .A3(new_n833), .A4(new_n910), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n929), .A2(G211gat), .A3(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n929), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n917), .A2(new_n295), .A3(new_n833), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1354gat));
  OAI21_X1  g737(.A(G218gat), .B1(new_n925), .B2(new_n596), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n917), .A2(new_n296), .A3(new_n595), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1355gat));
endmodule


