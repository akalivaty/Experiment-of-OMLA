//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT91), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(G8gat), .ZN(new_n211));
  INV_X1    g010(.A(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G43gat), .ZN(new_n213));
  INV_X1    g012(.A(G43gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G50gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT88), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(KEYINPUT88), .A3(G50gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n217), .A2(KEYINPUT89), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OR3_X1    g019(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n221), .A2(new_n222), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT15), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n219), .A2(new_n218), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT89), .B1(new_n227), .B2(new_n217), .ZN(new_n228));
  INV_X1    g027(.A(new_n225), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n223), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n226), .A2(new_n230), .A3(KEYINPUT92), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n221), .A2(new_n222), .ZN(new_n232));
  NAND2_X1  g031(.A1(G29gat), .A2(G36gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT89), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n218), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n234), .B1(new_n238), .B2(new_n225), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n229), .B1(new_n220), .B2(new_n223), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n239), .A2(KEYINPUT90), .A3(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(KEYINPUT17), .B(new_n231), .C1(new_n241), .C2(KEYINPUT92), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT92), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n230), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n243), .B(new_n244), .C1(new_n245), .C2(KEYINPUT90), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n211), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n238), .A2(new_n225), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n250), .A2(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n211), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n247), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT18), .ZN(new_n255));
  INV_X1    g054(.A(G8gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n210), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT90), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT92), .B1(new_n251), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n231), .A2(KEYINPUT17), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n246), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(new_n248), .A3(new_n252), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT18), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT93), .B1(new_n211), .B2(new_n251), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n257), .A2(new_n268), .A3(new_n245), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n252), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n248), .B(KEYINPUT13), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G113gat), .B(G141gat), .ZN(new_n274));
  INV_X1    g073(.A(G197gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT11), .B(G169gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT12), .ZN(new_n279));
  AND4_X1   g078(.A1(new_n255), .A2(new_n266), .A3(new_n273), .A4(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n270), .A2(new_n272), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n281), .B1(new_n264), .B2(new_n265), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n279), .B1(new_n282), .B2(new_n255), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n202), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n279), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n273), .B1(new_n254), .B2(KEYINPUT18), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n264), .A2(new_n265), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n282), .A2(new_n255), .A3(new_n279), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(KEYINPUT94), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293));
  XNOR2_X1  g092(.A(G127gat), .B(G134gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G134gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(KEYINPUT71), .A3(G127gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(KEYINPUT1), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT72), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G113gat), .B(G120gat), .Z(new_n302));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n294), .A2(new_n295), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .A4(new_n298), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n294), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(G141gat), .B(G148gat), .Z(new_n312));
  INV_X1    g111(.A(G155gat), .ZN(new_n313));
  INV_X1    g112(.A(G162gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR3_X1   g114(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT79), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n312), .B(KEYINPUT79), .C1(new_n315), .C2(new_n316), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(G155gat), .B(G162gat), .Z(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n293), .B1(new_n311), .B2(new_n325), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n301), .A2(new_n307), .B1(new_n294), .B2(new_n309), .ZN(new_n327));
  INV_X1    g126(.A(new_n325), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT4), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n319), .A2(new_n332), .A3(new_n324), .A4(new_n320), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT80), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n317), .A2(new_n318), .B1(new_n322), .B2(new_n323), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n332), .A4(new_n320), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT81), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n308), .A2(new_n310), .B1(new_n325), .B2(KEYINPUT3), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n330), .B(new_n331), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n327), .B(new_n325), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n344), .A2(new_n331), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n292), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n326), .A2(new_n329), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n338), .A2(new_n340), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT81), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n338), .A2(new_n340), .A3(new_n339), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT5), .B1(new_n351), .B2(new_n331), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT6), .ZN(new_n353));
  XOR2_X1   g152(.A(G57gat), .B(G85gat), .Z(new_n354));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR4_X1   g158(.A1(new_n346), .A2(new_n352), .A3(new_n353), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n292), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n343), .A2(new_n345), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n361), .B(new_n358), .C1(new_n362), .C2(new_n292), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n359), .B1(new_n346), .B2(new_n352), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n364), .A3(new_n353), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n360), .B1(new_n365), .B2(KEYINPUT87), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT87), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n363), .A2(new_n364), .A3(new_n367), .A4(new_n353), .ZN(new_n368));
  AND2_X1   g167(.A1(G211gat), .A2(G218gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(G197gat), .A2(G204gat), .ZN(new_n370));
  AND2_X1   g169(.A1(G197gat), .A2(G204gat), .ZN(new_n371));
  OAI22_X1  g170(.A1(new_n369), .A2(KEYINPUT22), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n372), .A2(KEYINPUT74), .ZN(new_n373));
  XOR2_X1   g172(.A(G211gat), .B(G218gat), .Z(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n377));
  INV_X1    g176(.A(G183gat), .ZN(new_n378));
  INV_X1    g177(.A(G190gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT64), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT24), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n385), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT64), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n382), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(KEYINPUT23), .ZN(new_n392));
  NAND2_X1  g191(.A1(G169gat), .A2(G176gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n392), .B(new_n393), .C1(new_n394), .C2(new_n390), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n377), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT66), .ZN(new_n397));
  INV_X1    g196(.A(new_n381), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n387), .B1(new_n398), .B2(KEYINPUT67), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(new_n380), .C1(KEYINPUT67), .C2(new_n387), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n395), .A2(new_n377), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n396), .A2(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n395), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n386), .A3(new_n388), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT25), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT66), .ZN(new_n406));
  INV_X1    g205(.A(new_n393), .ZN(new_n407));
  INV_X1    g206(.A(new_n390), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(KEYINPUT26), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(KEYINPUT26), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n383), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT27), .B(G183gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(KEYINPUT68), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT68), .B1(new_n378), .B2(KEYINPUT27), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n379), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(KEYINPUT28), .A3(new_n379), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT70), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n411), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(KEYINPUT70), .A3(new_n418), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n402), .A2(new_n406), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n376), .B1(new_n423), .B2(KEYINPUT29), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n420), .ZN(new_n425));
  INV_X1    g224(.A(new_n411), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n406), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n401), .A2(new_n400), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n405), .B2(KEYINPUT66), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n427), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n376), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n431), .A2(KEYINPUT76), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT76), .B1(new_n431), .B2(new_n432), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n375), .B(new_n424), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n375), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT75), .B(KEYINPUT29), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n432), .B1(new_n431), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n376), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT37), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n435), .A2(new_n444), .A3(new_n441), .ZN(new_n446));
  XNOR2_X1  g245(.A(G8gat), .B(G36gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(G92gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT77), .B(G64gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT38), .B1(new_n445), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n450), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n453), .A2(KEYINPUT38), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n439), .A2(new_n440), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n444), .B1(new_n455), .B2(new_n375), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n436), .B(new_n424), .C1(new_n433), .C2(new_n434), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n458), .A2(new_n446), .B1(new_n443), .B2(new_n453), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n366), .A2(new_n368), .A3(new_n452), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G228gat), .A2(G233gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT3), .B1(new_n375), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n437), .B1(new_n334), .B2(new_n337), .ZN(new_n465));
  OAI221_X1 g264(.A(new_n462), .B1(new_n464), .B2(new_n328), .C1(new_n465), .C2(new_n375), .ZN(new_n466));
  INV_X1    g265(.A(new_n374), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n372), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n438), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n467), .A2(new_n372), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n332), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n325), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n465), .B2(new_n375), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT83), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n473), .A2(new_n474), .A3(new_n461), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n473), .B2(new_n461), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(G22gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT85), .ZN(new_n479));
  INV_X1    g278(.A(G22gat), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n480), .B(new_n466), .C1(new_n475), .C2(new_n476), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G78gat), .B(G106gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT31), .B(G50gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n477), .B2(G22gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n481), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n478), .A2(new_n490), .A3(new_n481), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n477), .A2(KEYINPUT84), .A3(G22gat), .ZN(new_n492));
  INV_X1    g291(.A(new_n485), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI22_X1  g293(.A1(new_n482), .A2(new_n489), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n442), .A2(new_n450), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n435), .A2(new_n441), .A3(new_n453), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(KEYINPUT30), .A3(new_n497), .ZN(new_n498));
  OR3_X1    g297(.A1(new_n442), .A2(KEYINPUT30), .A3(new_n450), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n351), .B2(new_n331), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n330), .B1(new_n341), .B2(new_n342), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n503), .A2(KEYINPUT86), .A3(G225gat), .A4(G233gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT39), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n506), .B1(new_n344), .B2(new_n331), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n502), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n359), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT40), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n507), .A2(KEYINPUT40), .A3(new_n359), .A4(new_n509), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n500), .A2(new_n512), .A3(new_n363), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n460), .A2(new_n495), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT34), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n431), .A2(new_n311), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n423), .A2(new_n327), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G227gat), .A2(G233gat), .ZN(new_n523));
  OAI211_X1 g322(.A(KEYINPUT32), .B(new_n519), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G43gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G71gat), .B(G99gat), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  AOI21_X1  g327(.A(new_n523), .B1(new_n520), .B2(new_n521), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n525), .B(new_n528), .C1(new_n529), .C2(KEYINPUT33), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT33), .ZN(new_n531));
  INV_X1    g330(.A(new_n528), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n522), .B(new_n523), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT32), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT34), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n524), .A2(new_n530), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n533), .A2(new_n530), .B1(new_n524), .B2(new_n535), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n517), .B(new_n518), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n530), .A2(new_n533), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n535), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n542), .A2(KEYINPUT73), .A3(new_n516), .A4(new_n536), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n489), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n487), .A2(new_n488), .ZN(new_n546));
  INV_X1    g345(.A(new_n494), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n478), .A2(new_n490), .A3(new_n481), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n346), .A2(new_n352), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT6), .A3(new_n358), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n365), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n498), .A2(new_n499), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n544), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n515), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n365), .A2(new_n551), .B1(new_n498), .B2(new_n499), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n537), .A2(new_n538), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n495), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT35), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n366), .A2(new_n368), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT35), .B1(new_n498), .B2(new_n499), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n561), .A2(new_n558), .A3(new_n495), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n291), .B1(new_n556), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567));
  OAI211_X1 g366(.A(G85gat), .B(G92gat), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT96), .B1(KEYINPUT95), .B2(KEYINPUT7), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G99gat), .B(G106gat), .Z(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G99gat), .ZN(new_n573));
  INV_X1    g372(.A(G106gat), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT8), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(G85gat), .A2(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n570), .A2(new_n572), .A3(new_n575), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n575), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n568), .A2(new_n569), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n571), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT41), .ZN(new_n585));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586));
  OAI22_X1  g385(.A1(new_n245), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n242), .A2(new_n246), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(new_n584), .ZN(new_n589));
  XOR2_X1   g388(.A(G134gat), .B(G162gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G190gat), .B(G218gat), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n586), .A2(new_n585), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n591), .A2(new_n594), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G71gat), .B(G78gat), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT9), .ZN(new_n601));
  INV_X1    g400(.A(G71gat), .ZN(new_n602));
  INV_X1    g401(.A(G78gat), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G57gat), .B(G64gat), .Z(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n599), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT21), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n257), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n257), .B2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(new_n378), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G211gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n615), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G127gat), .B(G155gat), .Z(new_n620));
  XOR2_X1   g419(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n598), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n580), .A2(new_n583), .A3(new_n608), .A4(new_n606), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT97), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(KEYINPUT97), .A3(KEYINPUT10), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n584), .A2(new_n609), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n627), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(G230gat), .A3(G233gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT98), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n636), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n626), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n565), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n552), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(new_n205), .ZN(G1324gat));
  INV_X1    g448(.A(new_n647), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n500), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT16), .B(G8gat), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT99), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n653), .A2(KEYINPUT42), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(G8gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(KEYINPUT42), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(G1325gat));
  INV_X1    g456(.A(G15gat), .ZN(new_n658));
  INV_X1    g457(.A(new_n544), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n647), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n650), .A2(new_n558), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n658), .B2(new_n661), .ZN(G1326gat));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n495), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT43), .B(G22gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  INV_X1    g464(.A(new_n625), .ZN(new_n666));
  INV_X1    g465(.A(new_n645), .ZN(new_n667));
  AND4_X1   g466(.A1(new_n565), .A2(new_n666), .A3(new_n597), .A4(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n552), .A2(G29gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT100), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(new_n672), .A3(new_n669), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n671), .A2(KEYINPUT45), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT45), .B1(new_n671), .B2(new_n673), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n598), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n556), .B2(new_n564), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n549), .A2(new_n554), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT102), .B1(new_n495), .B2(new_n557), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n684), .A3(new_n659), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n460), .A2(new_n495), .A3(new_n514), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n564), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n597), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n681), .B1(new_n688), .B2(new_n678), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n280), .B2(new_n283), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n288), .A2(KEYINPUT101), .A3(new_n289), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n666), .A2(new_n667), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n689), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n677), .B1(new_n697), .B2(new_n552), .ZN(new_n698));
  INV_X1    g497(.A(new_n552), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n689), .A2(KEYINPUT103), .A3(new_n699), .A4(new_n696), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(G29gat), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n676), .A2(new_n701), .ZN(G1328gat));
  INV_X1    g501(.A(G36gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n668), .A2(new_n703), .A3(new_n500), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT46), .Z(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n697), .B2(new_n553), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1329gat));
  OAI21_X1  g506(.A(G43gat), .B1(new_n697), .B2(new_n659), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n668), .A2(new_n214), .A3(new_n558), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n708), .B2(new_n710), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(G1330gat));
  OAI21_X1  g512(.A(G50gat), .B1(new_n697), .B2(new_n495), .ZN(new_n714));
  NAND2_X1  g513(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n549), .A2(new_n212), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT104), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n668), .B2(new_n718), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n714), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n715), .B1(new_n714), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(G1331gat));
  NOR3_X1   g521(.A1(new_n626), .A2(new_n693), .A3(new_n667), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n687), .A2(new_n723), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n724), .A2(KEYINPUT106), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(KEYINPUT106), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n552), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT107), .B(G57gat), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1332gat));
  XOR2_X1   g529(.A(KEYINPUT108), .B(KEYINPUT109), .Z(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n725), .A2(new_n726), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n500), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT49), .B(G64gat), .Z(new_n735));
  NOR3_X1   g534(.A1(new_n727), .A2(new_n553), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n731), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n735), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n733), .A2(new_n500), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n731), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n727), .A2(new_n553), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n732), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n737), .A2(new_n742), .ZN(G1333gat));
  XNOR2_X1  g542(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n602), .B1(new_n733), .B2(new_n544), .ZN(new_n746));
  INV_X1    g545(.A(new_n558), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n727), .A2(G71gat), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n602), .A3(new_n558), .ZN(new_n750));
  OAI21_X1  g549(.A(G71gat), .B1(new_n727), .B2(new_n659), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(new_n751), .A3(new_n744), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1334gat));
  NOR2_X1   g552(.A1(new_n727), .A2(new_n495), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n603), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n693), .A2(new_n625), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n687), .A2(new_n597), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n515), .A2(new_n659), .A3(new_n683), .A4(new_n684), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n598), .B1(new_n760), .B2(new_n564), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n761), .B2(new_n756), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT112), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n757), .A2(new_n758), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n761), .A2(KEYINPUT51), .A3(new_n756), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n552), .A2(G85gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n763), .A2(new_n645), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n693), .A2(new_n625), .A3(new_n667), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n689), .A2(KEYINPUT111), .A3(new_n699), .A4(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n515), .A2(new_n555), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n495), .A2(new_n558), .A3(new_n562), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n774), .A2(new_n561), .B1(new_n559), .B2(KEYINPUT35), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n679), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n776), .B(new_n770), .C1(new_n761), .C2(KEYINPUT44), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n772), .B1(new_n777), .B2(new_n552), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n771), .A2(new_n778), .A3(G85gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n769), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n769), .A2(new_n779), .A3(KEYINPUT113), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1336gat));
  NAND3_X1  g583(.A1(new_n689), .A2(new_n500), .A3(new_n770), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n759), .A2(new_n762), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n553), .A2(G92gat), .A3(new_n667), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n788), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n789), .B(KEYINPUT114), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n792), .A2(new_n793), .B1(G92gat), .B2(new_n785), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n791), .B1(new_n794), .B2(new_n787), .ZN(G1337gat));
  OAI21_X1  g594(.A(G99gat), .B1(new_n777), .B2(new_n659), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n763), .A2(new_n645), .A3(new_n767), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n558), .A2(new_n573), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(G1338gat));
  OAI21_X1  g598(.A(G106gat), .B1(new_n777), .B2(new_n495), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n549), .A2(new_n574), .A3(new_n645), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n788), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n802), .B(new_n803), .Z(G1339gat));
  AOI22_X1  g603(.A1(new_n628), .A2(new_n629), .B1(new_n609), .B2(new_n584), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n805), .A2(new_n806), .A3(new_n631), .A4(new_n632), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n634), .A2(KEYINPUT54), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n631), .B1(new_n805), .B2(new_n632), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n642), .B(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n644), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  OAI211_X1 g614(.A(KEYINPUT116), .B(new_n644), .C1(new_n810), .C2(new_n811), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n691), .B2(new_n692), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n248), .B1(new_n263), .B2(new_n252), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n270), .A2(new_n272), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n278), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n289), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n667), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT117), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n817), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n288), .A2(KEYINPUT101), .A3(new_n289), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT101), .B1(new_n288), .B2(new_n289), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829));
  INV_X1    g628(.A(new_n823), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n824), .A2(new_n831), .A3(new_n598), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n598), .A2(new_n817), .A3(new_n822), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n625), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n646), .A2(new_n694), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n495), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n840), .B(new_n495), .C1(new_n835), .C2(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n500), .A2(new_n552), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n747), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n291), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n828), .A2(new_n830), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n597), .B1(new_n848), .B2(KEYINPUT117), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n833), .B1(new_n849), .B2(new_n831), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n836), .B1(new_n850), .B2(new_n625), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n495), .A3(new_n845), .ZN(new_n852));
  OR3_X1    g651(.A1(new_n852), .A2(G113gat), .A3(new_n694), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n847), .A2(new_n853), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n846), .B2(new_n667), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n852), .A2(G120gat), .A3(new_n667), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1341gat));
  INV_X1    g656(.A(new_n852), .ZN(new_n858));
  AOI21_X1  g657(.A(G127gat), .B1(new_n858), .B2(new_n625), .ZN(new_n859));
  INV_X1    g658(.A(new_n846), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n625), .A2(G127gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(G1342gat));
  OAI21_X1  g661(.A(G134gat), .B1(new_n846), .B2(new_n598), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n597), .A2(new_n297), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT56), .B1(new_n852), .B2(new_n864), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n852), .A2(KEYINPUT56), .A3(new_n864), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  INV_X1    g666(.A(G141gat), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n284), .A2(new_n290), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(KEYINPUT119), .A3(new_n830), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n598), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT119), .B1(new_n871), .B2(new_n830), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n871), .A2(new_n830), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n878), .A2(KEYINPUT120), .A3(new_n598), .A4(new_n872), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n875), .A2(new_n834), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n837), .B1(new_n880), .B2(new_n666), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT57), .B1(new_n881), .B2(new_n495), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n883), .B(new_n549), .C1(new_n835), .C2(new_n837), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n844), .A2(new_n544), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n291), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n868), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n835), .A2(new_n837), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n495), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n885), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n888), .A2(new_n868), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n882), .A2(new_n886), .A3(new_n693), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(G141gat), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n889), .A2(new_n895), .B1(new_n898), .B2(new_n890), .ZN(G1344gat));
  OR3_X1    g698(.A1(new_n893), .A2(G148gat), .A3(new_n667), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G148gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n887), .B2(new_n645), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n878), .A2(new_n598), .A3(new_n872), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n834), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n666), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n646), .A2(new_n291), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n625), .B1(new_n904), .B2(new_n834), .ZN(new_n910));
  INV_X1    g709(.A(new_n908), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT121), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n909), .A2(new_n912), .A3(new_n883), .A4(new_n549), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT57), .B1(new_n891), .B2(new_n495), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n913), .A2(new_n914), .A3(new_n645), .A4(new_n885), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n901), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n900), .B1(new_n903), .B2(new_n916), .ZN(G1345gat));
  INV_X1    g716(.A(new_n893), .ZN(new_n918));
  AOI21_X1  g717(.A(G155gat), .B1(new_n918), .B2(new_n625), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n666), .A2(new_n313), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n887), .B2(new_n920), .ZN(G1346gat));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n314), .A3(new_n597), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n887), .A2(new_n597), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n314), .ZN(G1347gat));
  NOR3_X1   g723(.A1(new_n699), .A2(new_n747), .A3(new_n553), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n495), .B(new_n925), .C1(new_n835), .C2(new_n837), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(G169gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n928), .A3(new_n693), .ZN(new_n929));
  INV_X1    g728(.A(new_n925), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n930), .B1(new_n839), .B2(new_n841), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(new_n888), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n932), .B2(new_n928), .ZN(G1348gat));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n842), .A2(new_n645), .A3(new_n925), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G176gat), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n926), .A2(G176gat), .A3(new_n667), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n934), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  AOI211_X1 g738(.A(KEYINPUT122), .B(new_n937), .C1(new_n935), .C2(G176gat), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(G1349gat));
  AOI21_X1  g740(.A(new_n840), .B1(new_n851), .B2(new_n495), .ZN(new_n942));
  INV_X1    g741(.A(new_n841), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n625), .B(new_n925), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(G183gat), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n625), .A2(new_n413), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n927), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT123), .B1(new_n926), .B2(new_n951), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n945), .A2(new_n948), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n948), .B1(new_n945), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(G1350gat));
  NOR3_X1   g757(.A1(new_n926), .A2(G190gat), .A3(new_n598), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT125), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n379), .B1(new_n931), .B2(new_n597), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(G1351gat));
  AND2_X1   g764(.A1(new_n913), .A2(new_n914), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n659), .A2(new_n552), .A3(new_n500), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n966), .A2(new_n888), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n659), .A2(new_n500), .A3(new_n549), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n972), .A2(new_n699), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n851), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n693), .A2(new_n275), .ZN(new_n975));
  OAI22_X1  g774(.A1(new_n969), .A2(new_n275), .B1(new_n974), .B2(new_n975), .ZN(G1352gat));
  OR3_X1    g775(.A1(new_n974), .A2(G204gat), .A3(new_n667), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n966), .A2(new_n645), .A3(new_n968), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G204gat), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(G1353gat));
  OR3_X1    g781(.A1(new_n974), .A2(G211gat), .A3(new_n666), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n913), .A2(new_n914), .A3(new_n625), .A4(new_n968), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(G1354gat));
  INV_X1    g786(.A(G218gat), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n598), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n913), .A2(new_n914), .A3(new_n968), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n988), .B1(new_n974), .B2(new_n598), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n992), .B(new_n993), .ZN(G1355gat));
endmodule


