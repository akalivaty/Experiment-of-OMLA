

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594;

  XNOR2_X1 U327 ( .A(n342), .B(n341), .ZN(n346) );
  XNOR2_X1 U328 ( .A(n367), .B(n366), .ZN(n368) );
  AND2_X1 U329 ( .A1(G230GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U330 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n356) );
  XNOR2_X1 U331 ( .A(n357), .B(n356), .ZN(n373) );
  XNOR2_X1 U332 ( .A(n340), .B(n339), .ZN(n341) );
  NOR2_X1 U333 ( .A1(n532), .A2(n504), .ZN(n418) );
  XNOR2_X1 U334 ( .A(n358), .B(n295), .ZN(n360) );
  XNOR2_X1 U335 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U336 ( .A(KEYINPUT36), .B(KEYINPUT78), .ZN(n355) );
  XNOR2_X1 U337 ( .A(n360), .B(n446), .ZN(n362) );
  XNOR2_X1 U338 ( .A(n350), .B(n349), .ZN(n354) );
  XNOR2_X1 U339 ( .A(n395), .B(n355), .ZN(n495) );
  XNOR2_X1 U340 ( .A(n369), .B(n368), .ZN(n372) );
  XNOR2_X1 U341 ( .A(n465), .B(G176GAT), .ZN(n466) );
  XNOR2_X1 U342 ( .A(n467), .B(n466), .ZN(G1349GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n297) );
  XNOR2_X1 U344 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U346 ( .A(KEYINPUT18), .B(n298), .Z(n415) );
  XOR2_X1 U347 ( .A(G190GAT), .B(G99GAT), .Z(n300) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U350 ( .A(KEYINPUT83), .B(KEYINPUT87), .Z(n302) );
  XNOR2_X1 U351 ( .A(G169GAT), .B(G15GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U353 ( .A(n304), .B(n303), .Z(n314) );
  XOR2_X1 U354 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n306) );
  XNOR2_X1 U355 ( .A(G176GAT), .B(KEYINPUT85), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n312) );
  XOR2_X1 U357 ( .A(G120GAT), .B(G71GAT), .Z(n358) );
  XOR2_X1 U358 ( .A(G127GAT), .B(KEYINPUT0), .Z(n308) );
  XNOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n440) );
  XOR2_X1 U361 ( .A(n358), .B(n440), .Z(n310) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n415), .B(n315), .ZN(n507) );
  XOR2_X1 U367 ( .A(KEYINPUT80), .B(G64GAT), .Z(n317) );
  XNOR2_X1 U368 ( .A(G8GAT), .B(G71GAT), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U370 ( .A(KEYINPUT79), .B(KEYINPUT81), .Z(n319) );
  XNOR2_X1 U371 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n332) );
  XOR2_X1 U374 ( .A(G57GAT), .B(KEYINPUT13), .Z(n370) );
  XOR2_X1 U375 ( .A(G22GAT), .B(G155GAT), .Z(n449) );
  XOR2_X1 U376 ( .A(n370), .B(n449), .Z(n323) );
  XNOR2_X1 U377 ( .A(G78GAT), .B(G211GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n328) );
  XNOR2_X1 U379 ( .A(G15GAT), .B(G1GAT), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n324), .B(KEYINPUT71), .ZN(n375) );
  XOR2_X1 U381 ( .A(KEYINPUT15), .B(n375), .Z(n326) );
  NAND2_X1 U382 ( .A1(G231GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U384 ( .A(n328), .B(n327), .Z(n330) );
  XNOR2_X1 U385 ( .A(G183GAT), .B(G127GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n589) );
  XNOR2_X1 U388 ( .A(G99GAT), .B(G106GAT), .ZN(n338) );
  INV_X1 U389 ( .A(G85GAT), .ZN(n333) );
  NAND2_X1 U390 ( .A1(KEYINPUT73), .A2(n333), .ZN(n336) );
  INV_X1 U391 ( .A(KEYINPUT73), .ZN(n334) );
  NAND2_X1 U392 ( .A1(n334), .A2(G85GAT), .ZN(n335) );
  NAND2_X1 U393 ( .A1(n336), .A2(n335), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n363) );
  XOR2_X1 U395 ( .A(G50GAT), .B(G162GAT), .Z(n450) );
  XNOR2_X1 U396 ( .A(n363), .B(n450), .ZN(n342) );
  AND2_X1 U397 ( .A1(G232GAT), .A2(G233GAT), .ZN(n340) );
  INV_X1 U398 ( .A(KEYINPUT10), .ZN(n339) );
  XOR2_X1 U399 ( .A(G29GAT), .B(G43GAT), .Z(n344) );
  XNOR2_X1 U400 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n378) );
  XNOR2_X1 U402 ( .A(n378), .B(KEYINPUT9), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U404 ( .A(G134GAT), .B(KEYINPUT76), .Z(n432) );
  XNOR2_X1 U405 ( .A(n432), .B(KEYINPUT11), .ZN(n348) );
  INV_X1 U406 ( .A(KEYINPUT75), .ZN(n347) );
  XOR2_X1 U407 ( .A(KEYINPUT77), .B(G92GAT), .Z(n352) );
  XNOR2_X1 U408 ( .A(G190GAT), .B(G218GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(n353), .ZN(n416) );
  XNOR2_X1 U411 ( .A(n354), .B(n416), .ZN(n395) );
  NOR2_X1 U412 ( .A1(n589), .A2(n495), .ZN(n357) );
  XNOR2_X1 U413 ( .A(G78GAT), .B(G204GAT), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n359), .B(G148GAT), .ZN(n446) );
  INV_X1 U415 ( .A(KEYINPUT31), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n369) );
  XNOR2_X1 U417 ( .A(n363), .B(KEYINPUT74), .ZN(n367) );
  XOR2_X1 U418 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n365) );
  XNOR2_X1 U419 ( .A(G92GAT), .B(KEYINPUT32), .ZN(n364) );
  XOR2_X1 U420 ( .A(n365), .B(n364), .Z(n366) );
  XOR2_X1 U421 ( .A(G176GAT), .B(G64GAT), .Z(n410) );
  XNOR2_X1 U422 ( .A(n370), .B(n410), .ZN(n371) );
  XNOR2_X1 U423 ( .A(n372), .B(n371), .ZN(n583) );
  NAND2_X1 U424 ( .A1(n373), .A2(n583), .ZN(n374) );
  XNOR2_X1 U425 ( .A(n374), .B(KEYINPUT111), .ZN(n391) );
  XOR2_X1 U426 ( .A(G169GAT), .B(G8GAT), .Z(n411) );
  XOR2_X1 U427 ( .A(n375), .B(n411), .Z(n377) );
  XNOR2_X1 U428 ( .A(G50GAT), .B(G36GAT), .ZN(n376) );
  XNOR2_X1 U429 ( .A(n377), .B(n376), .ZN(n382) );
  XOR2_X1 U430 ( .A(n378), .B(KEYINPUT30), .Z(n380) );
  NAND2_X1 U431 ( .A1(G229GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U433 ( .A(n382), .B(n381), .Z(n390) );
  XOR2_X1 U434 ( .A(G113GAT), .B(G22GAT), .Z(n384) );
  XNOR2_X1 U435 ( .A(G197GAT), .B(G141GAT), .ZN(n383) );
  XNOR2_X1 U436 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U437 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n386) );
  XNOR2_X1 U438 ( .A(KEYINPUT29), .B(KEYINPUT69), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U441 ( .A(n390), .B(n389), .ZN(n563) );
  INV_X1 U442 ( .A(n563), .ZN(n578) );
  NAND2_X1 U443 ( .A1(n391), .A2(n578), .ZN(n400) );
  XOR2_X1 U444 ( .A(KEYINPUT110), .B(KEYINPUT47), .Z(n398) );
  INV_X1 U445 ( .A(n589), .ZN(n566) );
  XNOR2_X1 U446 ( .A(n583), .B(KEYINPUT64), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n392), .B(KEYINPUT41), .ZN(n553) );
  NAND2_X1 U448 ( .A1(n563), .A2(n553), .ZN(n393) );
  XOR2_X1 U449 ( .A(KEYINPUT46), .B(n393), .Z(n394) );
  NOR2_X1 U450 ( .A1(n566), .A2(n394), .ZN(n396) );
  NAND2_X1 U451 ( .A1(n396), .A2(n395), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n399) );
  NAND2_X1 U453 ( .A1(n400), .A2(n399), .ZN(n402) );
  XOR2_X1 U454 ( .A(KEYINPUT112), .B(KEYINPUT48), .Z(n401) );
  XNOR2_X1 U455 ( .A(n402), .B(n401), .ZN(n532) );
  XOR2_X1 U456 ( .A(KEYINPUT97), .B(KEYINPUT99), .Z(n404) );
  XNOR2_X1 U457 ( .A(G204GAT), .B(KEYINPUT98), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n409) );
  XNOR2_X1 U459 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n405), .B(G211GAT), .ZN(n458) );
  XOR2_X1 U461 ( .A(n458), .B(KEYINPUT100), .Z(n407) );
  NAND2_X1 U462 ( .A1(G226GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U464 ( .A(n409), .B(n408), .Z(n413) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U466 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n415), .B(n414), .ZN(n417) );
  XNOR2_X1 U468 ( .A(n417), .B(n416), .ZN(n504) );
  XNOR2_X1 U469 ( .A(n418), .B(KEYINPUT54), .ZN(n443) );
  XOR2_X1 U470 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n420) );
  XNOR2_X1 U471 ( .A(G1GAT), .B(G57GAT), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U473 ( .A(KEYINPUT96), .B(KEYINPUT6), .Z(n422) );
  XNOR2_X1 U474 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U476 ( .A(n424), .B(n423), .Z(n429) );
  XOR2_X1 U477 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n426) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U480 ( .A(KEYINPUT5), .B(n427), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n437) );
  XOR2_X1 U482 ( .A(G85GAT), .B(G155GAT), .Z(n431) );
  XNOR2_X1 U483 ( .A(G120GAT), .B(G148GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U485 ( .A(n433), .B(n432), .Z(n435) );
  XNOR2_X1 U486 ( .A(G29GAT), .B(G162GAT), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U488 ( .A(n437), .B(n436), .Z(n442) );
  XOR2_X1 U489 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n439) );
  XNOR2_X1 U490 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n445) );
  XNOR2_X1 U492 ( .A(n440), .B(n445), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n501) );
  NAND2_X1 U494 ( .A1(n443), .A2(n501), .ZN(n444) );
  XNOR2_X1 U495 ( .A(n444), .B(KEYINPUT65), .ZN(n576) );
  XNOR2_X1 U496 ( .A(n446), .B(n445), .ZN(n462) );
  XOR2_X1 U497 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n448) );
  XNOR2_X1 U498 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n454) );
  XOR2_X1 U500 ( .A(G106GAT), .B(G218GAT), .Z(n452) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U503 ( .A(n454), .B(n453), .Z(n456) );
  NAND2_X1 U504 ( .A1(G228GAT), .A2(G233GAT), .ZN(n455) );
  XNOR2_X1 U505 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U506 ( .A(n457), .B(KEYINPUT91), .Z(n460) );
  XNOR2_X1 U507 ( .A(n458), .B(KEYINPUT90), .ZN(n459) );
  XNOR2_X1 U508 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U509 ( .A(n462), .B(n461), .ZN(n473) );
  AND2_X1 U510 ( .A1(n576), .A2(n473), .ZN(n463) );
  XNOR2_X1 U511 ( .A(n463), .B(KEYINPUT55), .ZN(n464) );
  NOR2_X2 U512 ( .A1(n507), .A2(n464), .ZN(n569) );
  NAND2_X1 U513 ( .A1(n569), .A2(n553), .ZN(n467) );
  XOR2_X1 U514 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n465) );
  XNOR2_X1 U515 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n487) );
  NAND2_X1 U516 ( .A1(n563), .A2(n583), .ZN(n498) );
  XNOR2_X1 U517 ( .A(n473), .B(KEYINPUT67), .ZN(n468) );
  XNOR2_X1 U518 ( .A(n468), .B(KEYINPUT28), .ZN(n528) );
  NOR2_X1 U519 ( .A1(n501), .A2(n528), .ZN(n469) );
  XOR2_X1 U520 ( .A(KEYINPUT27), .B(n504), .Z(n477) );
  NAND2_X1 U521 ( .A1(n469), .A2(n477), .ZN(n533) );
  XNOR2_X1 U522 ( .A(n533), .B(KEYINPUT101), .ZN(n470) );
  NAND2_X1 U523 ( .A1(n470), .A2(n507), .ZN(n482) );
  INV_X1 U524 ( .A(n507), .ZN(n535) );
  INV_X1 U525 ( .A(n504), .ZN(n525) );
  NAND2_X1 U526 ( .A1(n535), .A2(n525), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n473), .A2(n471), .ZN(n472) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(n472), .Z(n478) );
  XNOR2_X1 U529 ( .A(KEYINPUT103), .B(KEYINPUT26), .ZN(n475) );
  NOR2_X1 U530 ( .A1(n535), .A2(n473), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT102), .B(n476), .Z(n577) );
  NAND2_X1 U533 ( .A1(n577), .A2(n477), .ZN(n547) );
  NAND2_X1 U534 ( .A1(n478), .A2(n547), .ZN(n479) );
  XNOR2_X1 U535 ( .A(KEYINPUT104), .B(n479), .ZN(n480) );
  NAND2_X1 U536 ( .A1(n480), .A2(n501), .ZN(n481) );
  NAND2_X1 U537 ( .A1(n482), .A2(n481), .ZN(n494) );
  XNOR2_X1 U538 ( .A(KEYINPUT78), .B(n395), .ZN(n571) );
  NAND2_X1 U539 ( .A1(n571), .A2(n566), .ZN(n483) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n483), .Z(n484) );
  NAND2_X1 U541 ( .A1(n494), .A2(n484), .ZN(n485) );
  XOR2_X1 U542 ( .A(KEYINPUT105), .B(n485), .Z(n513) );
  NOR2_X1 U543 ( .A1(n498), .A2(n513), .ZN(n491) );
  INV_X1 U544 ( .A(n501), .ZN(n549) );
  NAND2_X1 U545 ( .A1(n491), .A2(n549), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U547 ( .A1(n491), .A2(n525), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U550 ( .A1(n491), .A2(n535), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U552 ( .A1(n491), .A2(n528), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT106), .ZN(n493) );
  XNOR2_X1 U554 ( .A(G22GAT), .B(n493), .ZN(G1327GAT) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n503) );
  NAND2_X1 U556 ( .A1(n589), .A2(n494), .ZN(n496) );
  NOR2_X1 U557 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n497), .B(KEYINPUT37), .ZN(n523) );
  NOR2_X1 U559 ( .A1(n523), .A2(n498), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT107), .B(KEYINPUT38), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n511) );
  NOR2_X1 U562 ( .A1(n501), .A2(n511), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n511), .A2(n504), .ZN(n505) );
  XOR2_X1 U565 ( .A(KEYINPUT108), .B(n505), .Z(n506) );
  XNOR2_X1 U566 ( .A(G36GAT), .B(n506), .ZN(G1329GAT) );
  NOR2_X1 U567 ( .A1(n511), .A2(n507), .ZN(n508) );
  XOR2_X1 U568 ( .A(KEYINPUT40), .B(n508), .Z(n509) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n509), .ZN(G1330GAT) );
  INV_X1 U570 ( .A(n528), .ZN(n510) );
  NOR2_X1 U571 ( .A1(n511), .A2(n510), .ZN(n512) );
  XOR2_X1 U572 ( .A(G50GAT), .B(n512), .Z(G1331GAT) );
  NAND2_X1 U573 ( .A1(n553), .A2(n578), .ZN(n522) );
  NOR2_X1 U574 ( .A1(n522), .A2(n513), .ZN(n514) );
  XOR2_X1 U575 ( .A(KEYINPUT109), .B(n514), .Z(n519) );
  NAND2_X1 U576 ( .A1(n549), .A2(n519), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n515), .B(KEYINPUT42), .ZN(n516) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n516), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n519), .A2(n525), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n517), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n519), .A2(n535), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U584 ( .A1(n519), .A2(n528), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NOR2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n529), .A2(n549), .ZN(n524) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n529), .A2(n525), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n529), .A2(n535), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n532), .A2(n533), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n544) );
  NOR2_X1 U598 ( .A1(n578), .A2(n544), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  INV_X1 U601 ( .A(n553), .ZN(n538) );
  NOR2_X1 U602 ( .A1(n538), .A2(n544), .ZN(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  NOR2_X1 U606 ( .A1(n589), .A2(n544), .ZN(n542) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(n542), .Z(n543) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  NOR2_X1 U609 ( .A1(n571), .A2(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n532), .A2(n547), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n550), .B(KEYINPUT115), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n559), .A2(n563), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n551), .B(KEYINPUT116), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n555) );
  NAND2_X1 U619 ( .A1(n559), .A2(n553), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .Z(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n566), .A2(n559), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U625 ( .A(n559), .ZN(n560) );
  NOR2_X1 U626 ( .A1(n395), .A2(n560), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT118), .B(n561), .Z(n562) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(n562), .ZN(G1347GAT) );
  XOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT119), .Z(n565) );
  NAND2_X1 U630 ( .A1(n569), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n569), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT120), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U635 ( .A(n569), .ZN(n570) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n575) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT121), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT122), .B(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1351GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n577), .ZN(n591) );
  NOR2_X1 U642 ( .A1(n591), .A2(n578), .ZN(n582) );
  XOR2_X1 U643 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n591), .ZN(n588) );
  XOR2_X1 U648 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n585) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(KEYINPUT124), .B(n586), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n591), .ZN(n590) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n590), .Z(G1354GAT) );
  NOR2_X1 U655 ( .A1(n495), .A2(n591), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

