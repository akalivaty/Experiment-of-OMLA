//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT68), .ZN(new_n203));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208));
  NAND2_X1  g007(.A1(G113gat), .A2(G120gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(KEYINPUT69), .B(KEYINPUT1), .Z(new_n211));
  NAND4_X1  g010(.A1(new_n203), .A2(new_n204), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n204), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(KEYINPUT1), .B2(new_n202), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(G183gat), .A3(G190gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(G183gat), .B(G190gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(new_n217), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n222), .B(new_n218), .C1(new_n219), .C2(new_n217), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G169gat), .ZN(new_n228));
  INV_X1    g027(.A(G176gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n230), .B1(KEYINPUT23), .B2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n221), .A2(new_n223), .A3(new_n227), .A4(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n233), .A2(KEYINPUT25), .ZN(new_n234));
  INV_X1    g033(.A(new_n231), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n230), .B1(KEYINPUT26), .B2(new_n235), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n235), .A2(KEYINPUT26), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n236), .A2(new_n237), .B1(G183gat), .B2(G190gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G183gat), .ZN(new_n240));
  INV_X1    g039(.A(G183gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT27), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(G190gat), .B1(new_n240), .B2(KEYINPUT67), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT28), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT28), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n243), .A2(new_n248), .A3(G190gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n238), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n228), .A2(KEYINPUT64), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G169gat), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT23), .A4(new_n229), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n230), .A2(KEYINPUT25), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(new_n220), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n227), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n216), .B1(new_n234), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G227gat), .ZN(new_n261));
  INV_X1    g060(.A(G233gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT27), .B(G183gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT67), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n266));
  INV_X1    g065(.A(G190gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n248), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n249), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n271), .A2(new_n238), .B1(new_n227), .B2(new_n257), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n233), .A2(KEYINPUT25), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n215), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n260), .A2(new_n263), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n260), .A2(KEYINPUT70), .A3(new_n263), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT32), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT33), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G15gat), .B(G43gat), .Z(new_n283));
  XNOR2_X1  g082(.A(G71gat), .B(G99gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n277), .B2(new_n278), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT33), .B1(new_n277), .B2(new_n278), .ZN(new_n289));
  INV_X1    g088(.A(new_n285), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n260), .A2(new_n274), .ZN(new_n292));
  INV_X1    g091(.A(new_n263), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT34), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT34), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(new_n296), .A3(new_n293), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n286), .A2(new_n291), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G228gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(new_n262), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G155gat), .B(G162gat), .ZN(new_n303));
  OR2_X1    g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT76), .B(G162gat), .ZN(new_n307));
  INV_X1    g106(.A(G155gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT2), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311));
  INV_X1    g110(.A(new_n303), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT2), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n304), .A2(new_n313), .A3(new_n305), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n310), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G211gat), .B(G218gat), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(KEYINPUT73), .A2(G197gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(KEYINPUT73), .A2(G197gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G204gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(G204gat), .A3(new_n322), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n320), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AOI211_X1 g129(.A(new_n328), .B(new_n319), .C1(new_n325), .C2(new_n326), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n302), .B1(new_n318), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n317), .B1(new_n330), .B2(new_n331), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT82), .ZN(new_n336));
  INV_X1    g135(.A(new_n326), .ZN(new_n337));
  AOI21_X1  g136(.A(G204gat), .B1(new_n321), .B2(new_n322), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n329), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n319), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n327), .A2(new_n320), .A3(new_n329), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT82), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(new_n317), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n336), .A2(new_n344), .A3(new_n311), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT76), .B(G162gat), .Z(new_n346));
  AOI21_X1  g145(.A(new_n313), .B1(new_n346), .B2(G155gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n315), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n334), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n318), .A2(new_n332), .B1(KEYINPUT3), .B2(new_n349), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n317), .A3(new_n349), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n301), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(G22gat), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n352), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n302), .ZN(new_n356));
  INV_X1    g155(.A(G22gat), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n306), .A2(new_n309), .B1(new_n314), .B2(new_n312), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT3), .B1(new_n335), .B2(KEYINPUT82), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n344), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n356), .B(new_n357), .C1(new_n360), .C2(new_n334), .ZN(new_n361));
  XNOR2_X1  g160(.A(G78gat), .B(G106gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT31), .B(G50gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  NAND4_X1  g163(.A1(new_n354), .A2(new_n361), .A3(KEYINPUT83), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n354), .A2(new_n361), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n349), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n353), .B1(new_n367), .B2(new_n333), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT83), .B1(new_n368), .B2(new_n357), .ZN(new_n369));
  INV_X1    g168(.A(new_n364), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n299), .A2(new_n365), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT71), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n374));
  AOI221_X4 g173(.A(new_n287), .B1(KEYINPUT33), .B2(new_n285), .C1(new_n277), .C2(new_n278), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n298), .B(KEYINPUT72), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n286), .A2(KEYINPUT71), .A3(new_n291), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(new_n316), .A3(new_n215), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n310), .A2(new_n212), .A3(new_n315), .A4(new_n214), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n358), .A2(KEYINPUT4), .A3(new_n214), .A4(new_n212), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n382), .A2(new_n383), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n349), .A2(new_n215), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n384), .ZN(new_n390));
  INV_X1    g189(.A(new_n383), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT77), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n393));
  AOI211_X1 g192(.A(new_n393), .B(new_n383), .C1(new_n389), .C2(new_n384), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT5), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n380), .B(new_n388), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n349), .A2(new_n215), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n310), .A2(new_n315), .B1(new_n212), .B2(new_n214), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n391), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n393), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n390), .A2(KEYINPUT77), .A3(new_n391), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n388), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n380), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(KEYINPUT5), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G57gat), .B(G85gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT80), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n405), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n397), .B2(new_n405), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n414), .B(new_n413), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  AOI211_X1 g217(.A(KEYINPUT81), .B(new_n412), .C1(new_n397), .C2(new_n405), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n317), .B1(new_n234), .B2(new_n259), .ZN(new_n425));
  NAND2_X1  g224(.A1(G226gat), .A2(G233gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n273), .A2(new_n250), .A3(new_n258), .ZN(new_n428));
  INV_X1    g227(.A(new_n426), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT75), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  AOI211_X1 g230(.A(new_n431), .B(new_n426), .C1(new_n272), .C2(new_n273), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n427), .B(new_n342), .C1(new_n430), .C2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT74), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n429), .B1(new_n428), .B2(new_n317), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n426), .B1(new_n272), .B2(new_n273), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n434), .B(new_n332), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n429), .B1(new_n234), .B2(new_n259), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT29), .B1(new_n272), .B2(new_n273), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(new_n429), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n434), .B1(new_n441), .B2(new_n332), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n424), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n436), .B1(new_n425), .B2(new_n426), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT74), .B1(new_n444), .B2(new_n342), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n445), .A2(new_n433), .A3(new_n437), .A4(new_n423), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(KEYINPUT30), .A3(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n433), .A2(new_n437), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n445), .A4(new_n423), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n372), .A2(new_n379), .A3(new_n420), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n420), .A2(new_n451), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(KEYINPUT35), .ZN(new_n455));
  INV_X1    g254(.A(new_n298), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n374), .B2(new_n375), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n299), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n371), .A2(new_n365), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  INV_X1    g262(.A(new_n316), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n215), .B1(new_n358), .B2(new_n311), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n386), .B(new_n387), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n391), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n389), .A2(new_n383), .A3(new_n384), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n389), .A2(new_n470), .A3(new_n384), .A4(new_n383), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n467), .A2(new_n472), .A3(KEYINPUT39), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n466), .A2(new_n474), .A3(new_n391), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n411), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n463), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n467), .A2(new_n472), .A3(KEYINPUT39), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n478), .A2(KEYINPUT40), .A3(new_n411), .A4(new_n475), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n413), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n447), .A2(new_n450), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n371), .A2(new_n365), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n397), .A2(new_n405), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n411), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n416), .A2(new_n417), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(new_n414), .A3(new_n487), .A4(new_n413), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n445), .A2(new_n433), .A3(new_n437), .A4(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT37), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n441), .B2(new_n342), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n427), .B(new_n332), .C1(new_n430), .C2(new_n432), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT38), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n494), .A3(new_n424), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n495), .A2(new_n446), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n491), .B1(new_n448), .B2(new_n445), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n490), .A2(new_n424), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT38), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n488), .A2(new_n496), .A3(new_n499), .A4(new_n415), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n483), .A2(new_n500), .B1(new_n454), .B2(new_n459), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n299), .A2(KEYINPUT36), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n379), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n458), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n462), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(G197gat), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT11), .B(G169gat), .Z(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT12), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n357), .A2(G15gat), .ZN(new_n514));
  INV_X1    g313(.A(G15gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G22gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G1gat), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT89), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G8gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT16), .B1(new_n521), .B2(G1gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n518), .A2(KEYINPUT88), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n514), .B(new_n516), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n519), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n520), .B1(new_n519), .B2(new_n524), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528));
  INV_X1    g327(.A(G29gat), .ZN(new_n529));
  INV_X1    g328(.A(G36gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT14), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n531), .B(new_n533), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  NOR2_X1   g334(.A1(G43gat), .A2(G50gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G43gat), .A2(G50gat), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(KEYINPUT87), .A2(G29gat), .A3(G36gat), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT87), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G43gat), .A2(G50gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT15), .B1(new_n544), .B2(new_n536), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n543), .A2(new_n545), .A3(new_n533), .A4(new_n531), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n538), .A2(new_n535), .ZN(new_n547));
  AND2_X1   g346(.A1(KEYINPUT86), .A2(G50gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(KEYINPUT86), .A2(G50gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G43gat), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n528), .B(new_n540), .C1(new_n546), .C2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n555));
  INV_X1    g354(.A(G50gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(KEYINPUT86), .A2(G50gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n551), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n547), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n531), .A2(new_n533), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n561), .A2(new_n562), .A3(new_n545), .A4(new_n543), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n528), .B1(new_n563), .B2(new_n540), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n527), .B1(new_n554), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n540), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(new_n526), .B2(new_n525), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT90), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n513), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n565), .A2(KEYINPUT18), .A3(new_n566), .A4(new_n568), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n566), .B(KEYINPUT13), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n567), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n527), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n578), .B2(new_n568), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n571), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n579), .B1(new_n569), .B2(new_n570), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT90), .B1(new_n569), .B2(new_n570), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n583), .B(new_n574), .C1(new_n584), .C2(new_n513), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT9), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n589), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n591), .B(new_n590), .C1(new_n588), .C2(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n527), .B1(new_n587), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(G231gat), .A3(G233gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n597), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT92), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G183gat), .B(G211gat), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n603), .A2(new_n608), .A3(new_n605), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n612), .B1(new_n610), .B2(new_n613), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n600), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  INV_X1    g417(.A(new_n600), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n619), .A3(new_n614), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT8), .ZN(new_n623));
  NAND2_X1  g422(.A1(G85gat), .A2(G92gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT7), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G85gat), .ZN(new_n627));
  INV_X1    g426(.A(G92gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n623), .A2(new_n626), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT93), .ZN(new_n632));
  XNOR2_X1  g431(.A(G99gat), .B(G106gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n634), .ZN(new_n636));
  AOI22_X1  g435(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n627), .B2(new_n628), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n637), .A2(new_n633), .A3(new_n626), .A4(new_n630), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(KEYINPUT93), .A3(new_n638), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n635), .B(new_n639), .C1(new_n554), .C2(new_n564), .ZN(new_n640));
  XOR2_X1   g439(.A(G190gat), .B(G218gat), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n635), .ZN(new_n643));
  AND2_X1   g442(.A1(G232gat), .A2(G233gat), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n643), .A2(new_n567), .B1(KEYINPUT41), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n640), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n642), .B1(new_n640), .B2(new_n645), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n644), .A2(KEYINPUT41), .ZN(new_n648));
  XNOR2_X1  g447(.A(G134gat), .B(G162gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OR3_X1    g450(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n646), .B2(new_n647), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n639), .A2(new_n597), .A3(new_n635), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n595), .A2(new_n636), .A3(new_n596), .A4(new_n638), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT94), .B(KEYINPUT10), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT95), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT95), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n662), .A2(new_n667), .A3(new_n663), .A4(new_n664), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT10), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n643), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n661), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n662), .A2(new_n663), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n661), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT96), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n659), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n674), .B(new_n677), .ZN(new_n678));
  AOI22_X1  g477(.A1(new_n666), .A2(new_n668), .B1(new_n643), .B2(new_n670), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n678), .B(new_n658), .C1(new_n679), .C2(new_n661), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n621), .A2(new_n655), .A3(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT97), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT97), .ZN(new_n684));
  AND4_X1   g483(.A1(new_n508), .A2(new_n586), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n420), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  INV_X1    g487(.A(new_n451), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  AND3_X1   g489(.A1(new_n685), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n520), .B1(new_n685), .B2(new_n689), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT42), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(KEYINPUT42), .B2(new_n691), .ZN(G1325gat));
  INV_X1    g493(.A(new_n458), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n685), .A2(new_n515), .A3(new_n695), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n379), .A2(new_n502), .B1(new_n458), .B2(new_n504), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n685), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(new_n515), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n685), .A2(new_n459), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  INV_X1    g501(.A(new_n621), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n681), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n655), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT98), .Z(new_n706));
  NAND2_X1  g505(.A1(new_n481), .A2(new_n482), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n495), .A2(new_n446), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n420), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(new_n499), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n482), .B1(new_n420), .B2(new_n451), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(new_n697), .A3(new_n711), .ZN(new_n712));
  AOI22_X1  g511(.A1(KEYINPUT35), .A2(new_n452), .B1(new_n455), .B2(new_n460), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n586), .B(new_n706), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(G29gat), .A3(new_n420), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT99), .B(KEYINPUT45), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n453), .A2(new_n461), .B1(new_n501), .B2(new_n506), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(new_n654), .ZN(new_n720));
  OAI211_X1 g519(.A(KEYINPUT44), .B(new_n655), .C1(new_n712), .C2(new_n713), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT100), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n586), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n582), .A2(new_n585), .A3(KEYINPUT100), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n704), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT101), .Z(new_n728));
  AND4_X1   g527(.A1(new_n686), .A2(new_n720), .A3(new_n721), .A4(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n717), .B1(new_n529), .B2(new_n729), .ZN(G1328gat));
  NAND4_X1  g529(.A1(new_n720), .A2(new_n689), .A3(new_n721), .A4(new_n728), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G36gat), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n451), .A2(G36gat), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n508), .A2(new_n586), .A3(new_n706), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n732), .A2(KEYINPUT102), .A3(new_n735), .A4(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(G1329gat));
  OAI21_X1  g540(.A(new_n551), .B1(new_n714), .B2(new_n458), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n720), .A2(new_n721), .A3(new_n728), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n697), .A2(G43gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g545(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n459), .A2(new_n550), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n714), .B2(KEYINPUT103), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n508), .A2(new_n750), .A3(new_n586), .A4(new_n706), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n747), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n720), .A2(new_n459), .A3(new_n721), .A4(new_n728), .ZN(new_n753));
  INV_X1    g552(.A(new_n550), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT105), .Z(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n752), .A2(new_n755), .A3(new_n758), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1331gat));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n763));
  INV_X1    g562(.A(new_n681), .ZN(new_n764));
  NOR4_X1   g563(.A1(new_n726), .A2(new_n621), .A3(new_n655), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n508), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n765), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT106), .B1(new_n719), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n686), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g570(.A(new_n451), .B(KEYINPUT107), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  OR2_X1    g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1333gat));
  NOR2_X1   g575(.A1(new_n458), .A2(G71gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n769), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n766), .A2(new_n768), .ZN(new_n779));
  OAI21_X1  g578(.A(G71gat), .B1(new_n779), .B2(new_n506), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(new_n780), .A3(KEYINPUT50), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1334gat));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n459), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT108), .B(G78gat), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n786), .B(new_n787), .ZN(G1335gat));
  NAND3_X1  g587(.A1(new_n686), .A2(new_n627), .A3(new_n681), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n726), .A2(new_n703), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n655), .B(new_n791), .C1(new_n712), .C2(new_n713), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n654), .B1(new_n462), .B2(new_n507), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT51), .B1(new_n795), .B2(new_n791), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n791), .A2(new_n681), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n720), .A2(new_n686), .A3(new_n721), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G85gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT109), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n797), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(G1336gat));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n792), .A2(new_n807), .A3(KEYINPUT51), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n792), .B2(new_n807), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n772), .A2(G92gat), .A3(new_n764), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n720), .A2(new_n689), .A3(new_n721), .A4(new_n799), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(G92gat), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT52), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n720), .A2(new_n721), .A3(new_n799), .ZN(new_n816));
  OAI21_X1  g615(.A(G92gat), .B1(new_n816), .B2(new_n772), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n794), .A2(new_n796), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n811), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n815), .A2(new_n820), .ZN(G1337gat));
  NAND4_X1  g620(.A1(new_n720), .A2(new_n697), .A3(new_n721), .A4(new_n799), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G99gat), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n822), .A2(new_n823), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n458), .A2(G99gat), .A3(new_n764), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n825), .A2(new_n826), .B1(new_n819), .B2(new_n827), .ZN(G1338gat));
  NOR3_X1   g627(.A1(new_n482), .A2(G106gat), .A3(new_n764), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n808), .A2(new_n809), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n720), .A2(new_n459), .A3(new_n721), .A4(new_n799), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(G106gat), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT53), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(G106gat), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n835), .B(new_n836), .C1(new_n819), .C2(new_n830), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(G1339gat));
  INV_X1    g637(.A(new_n680), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n658), .B1(new_n672), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  INV_X1    g641(.A(new_n672), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n660), .B1(new_n643), .B2(new_n670), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n840), .B1(new_n669), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n842), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n839), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n669), .A2(new_n844), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n848), .B(KEYINPUT54), .C1(new_n679), .C2(new_n661), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n841), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n842), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n847), .A2(new_n724), .A3(new_n723), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n566), .B1(new_n565), .B2(new_n568), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n578), .A2(new_n568), .A3(new_n576), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n512), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n583), .A2(new_n513), .A3(new_n574), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n681), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n655), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT55), .B1(new_n859), .B2(new_n672), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n669), .A2(new_n671), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n840), .A3(new_n660), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n659), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n680), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT55), .B1(new_n841), .B2(new_n849), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n652), .A2(new_n856), .A3(new_n653), .A4(new_n855), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n621), .B1(new_n858), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n682), .A2(KEYINPUT112), .A3(new_n725), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT112), .B1(new_n682), .B2(new_n725), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n460), .ZN(new_n873));
  INV_X1    g672(.A(new_n772), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n420), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n205), .B1(new_n876), .B2(new_n586), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT113), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n420), .B1(new_n868), .B2(new_n871), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n372), .A2(new_n379), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n879), .A2(new_n880), .A3(new_n772), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n205), .A3(new_n726), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n882), .ZN(G1340gat));
  AOI21_X1  g682(.A(G120gat), .B1(new_n881), .B2(new_n681), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n764), .A2(new_n206), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n876), .B2(new_n885), .ZN(G1341gat));
  INV_X1    g685(.A(new_n876), .ZN(new_n887));
  OAI21_X1  g686(.A(G127gat), .B1(new_n887), .B2(new_n621), .ZN(new_n888));
  INV_X1    g687(.A(G127gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n881), .A2(new_n889), .A3(new_n703), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1342gat));
  INV_X1    g690(.A(G134gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n689), .A2(new_n654), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n879), .A2(new_n892), .A3(new_n880), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT114), .ZN(new_n896));
  OAI21_X1  g695(.A(G134gat), .B1(new_n887), .B2(new_n654), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n896), .B(new_n897), .C1(KEYINPUT56), .C2(new_n894), .ZN(G1343gat));
  NOR3_X1   g697(.A1(new_n874), .A2(new_n697), .A3(new_n420), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n872), .B2(new_n459), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n459), .A2(KEYINPUT57), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n849), .A2(KEYINPUT55), .A3(new_n659), .A4(new_n862), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n851), .A2(new_n586), .A3(new_n680), .A4(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n655), .B1(new_n903), .B2(new_n857), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n621), .B1(new_n904), .B2(new_n867), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n905), .B2(new_n871), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n899), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n586), .ZN(new_n908));
  OAI21_X1  g707(.A(G141gat), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  OR3_X1    g709(.A1(new_n697), .A2(KEYINPUT115), .A3(new_n482), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT115), .B1(new_n697), .B2(new_n482), .ZN(new_n912));
  AND4_X1   g711(.A1(new_n772), .A2(new_n911), .A3(new_n879), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n908), .A2(G141gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n909), .A2(new_n910), .A3(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n726), .B(new_n899), .C1(new_n900), .C2(new_n906), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G141gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n915), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT116), .B1(new_n919), .B2(KEYINPUT58), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n921));
  AOI211_X1 g720(.A(new_n921), .B(new_n910), .C1(new_n918), .C2(new_n915), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n916), .B1(new_n920), .B2(new_n922), .ZN(G1344gat));
  INV_X1    g722(.A(G148gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n913), .A2(new_n924), .A3(new_n681), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n872), .A2(KEYINPUT57), .A3(new_n459), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n683), .A2(new_n908), .A3(new_n684), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n902), .A2(new_n586), .A3(new_n680), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n857), .B1(new_n929), .B2(new_n865), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n867), .B1(new_n930), .B2(new_n654), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n621), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n904), .A2(KEYINPUT117), .A3(new_n867), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT57), .B1(new_n935), .B2(new_n459), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n927), .B1(new_n936), .B2(KEYINPUT118), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n938));
  AOI211_X1 g737(.A(new_n938), .B(KEYINPUT57), .C1(new_n935), .C2(new_n459), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n681), .B(new_n899), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n926), .B1(new_n940), .B2(G148gat), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n926), .A2(G148gat), .ZN(new_n942));
  INV_X1    g741(.A(new_n907), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n681), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n925), .B1(new_n941), .B2(new_n944), .ZN(G1345gat));
  AOI21_X1  g744(.A(G155gat), .B1(new_n913), .B2(new_n703), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n703), .A2(G155gat), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT119), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n943), .B2(new_n948), .ZN(G1346gat));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n943), .A2(new_n950), .A3(new_n655), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n346), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n943), .B2(new_n655), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n911), .A2(new_n879), .A3(new_n912), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n893), .A2(new_n307), .ZN(new_n955));
  OAI22_X1  g754(.A1(new_n952), .A2(new_n953), .B1(new_n954), .B2(new_n955), .ZN(G1347gat));
  NAND2_X1  g755(.A1(new_n872), .A2(new_n420), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT121), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n874), .A2(new_n880), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT122), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n251), .A2(new_n253), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NOR4_X1   g762(.A1(new_n961), .A2(KEYINPUT123), .A3(new_n963), .A4(new_n725), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT123), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n958), .A2(new_n960), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n725), .A2(new_n963), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n686), .A2(new_n451), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n873), .A2(new_n586), .A3(new_n969), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT124), .B1(new_n970), .B2(G169gat), .ZN(new_n972));
  OAI22_X1  g771(.A1(new_n964), .A2(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1348gat));
  NAND2_X1  g772(.A1(new_n873), .A2(new_n969), .ZN(new_n974));
  OAI21_X1  g773(.A(G176gat), .B1(new_n974), .B2(new_n764), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n681), .A2(new_n229), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n961), .B2(new_n976), .ZN(G1349gat));
  OAI21_X1  g776(.A(G183gat), .B1(new_n974), .B2(new_n621), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n703), .A2(new_n264), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n961), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT60), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT60), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n982), .B(new_n978), .C1(new_n961), .C2(new_n979), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1350gat));
  OAI21_X1  g783(.A(G190gat), .B1(new_n974), .B2(new_n654), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT125), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n987), .A2(KEYINPUT61), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n966), .A2(new_n267), .A3(new_n655), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n985), .A2(new_n986), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n987), .A2(KEYINPUT61), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n988), .B(new_n989), .C1(new_n990), .C2(new_n991), .ZN(G1351gat));
  NOR3_X1   g791(.A1(new_n697), .A2(new_n772), .A3(new_n482), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n958), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(G197gat), .B1(new_n994), .B2(new_n726), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n937), .A2(new_n939), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n697), .A2(new_n686), .A3(new_n451), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n586), .A2(G197gat), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(G1352gat));
  NAND3_X1  g799(.A1(new_n996), .A2(new_n681), .A3(new_n997), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(G204gat), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n1003));
  AOI211_X1 g802(.A(G204gat), .B(new_n764), .C1(new_n1003), .C2(KEYINPUT62), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n957), .A2(KEYINPUT121), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n957), .A2(KEYINPUT121), .ZN(new_n1006));
  OAI211_X1 g805(.A(new_n993), .B(new_n1004), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1002), .A2(new_n1009), .ZN(G1353gat));
  INV_X1    g809(.A(G211gat), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n994), .A2(new_n1011), .A3(new_n703), .ZN(new_n1012));
  OAI211_X1 g811(.A(new_n703), .B(new_n997), .C1(new_n937), .C2(new_n939), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n1013), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1014));
  AOI21_X1  g813(.A(KEYINPUT63), .B1(new_n1013), .B2(G211gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(G1354gat));
  NAND3_X1  g815(.A1(new_n996), .A2(new_n655), .A3(new_n997), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(G218gat), .ZN(new_n1018));
  INV_X1    g817(.A(G218gat), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n994), .A2(new_n1019), .A3(new_n655), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1018), .A2(new_n1020), .ZN(G1355gat));
endmodule


