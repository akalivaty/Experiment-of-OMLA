//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT66), .B(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n464), .A2(KEYINPUT67), .A3(G137), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n461), .A2(KEYINPUT66), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(new_n462), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n470), .A2(G137), .A3(new_n465), .A4(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n466), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT68), .B1(new_n463), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n468), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n461), .A2(KEYINPUT66), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n477), .B(new_n465), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(KEYINPUT69), .B1(new_n481), .B2(G101), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  INV_X1    g058(.A(G101), .ZN(new_n484));
  AOI211_X1 g059(.A(new_n483), .B(new_n484), .C1(new_n476), .C2(new_n480), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n475), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT70), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(new_n475), .C1(new_n482), .C2(new_n485), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n491), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n492), .A2(new_n465), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G160));
  INV_X1    g070(.A(new_n464), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G136), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n496), .A2(new_n465), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G124), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n465), .A2(G112), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n498), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n503), .B(KEYINPUT71), .ZN(G162));
  AND2_X1   g079(.A1(new_n465), .A2(G138), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n470), .A2(new_n471), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT73), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n505), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n506), .A2(KEYINPUT4), .B1(new_n511), .B2(new_n491), .ZN(new_n512));
  AND2_X1   g087(.A1(G126), .A2(G2105), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n470), .A2(new_n471), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  INV_X1    g092(.A(G114), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(G2105), .ZN(new_n519));
  NOR3_X1   g094(.A1(new_n465), .A2(KEYINPUT72), .A3(G114), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n512), .A2(new_n522), .ZN(G164));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G166));
  AND2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n525), .A2(KEYINPUT74), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n541), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  INV_X1    g119(.A(G51), .ZN(new_n545));
  INV_X1    g120(.A(G89), .ZN(new_n546));
  OAI221_X1 g121(.A(new_n544), .B1(new_n528), .B2(new_n545), .C1(new_n546), .C2(new_n526), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n542), .A2(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(new_n541), .A2(G64), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n532), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  INV_X1    g127(.A(G52), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n526), .A2(new_n552), .B1(new_n528), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(G171));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT75), .B(G43), .Z(new_n557));
  OAI22_X1  g132(.A1(new_n526), .A2(new_n556), .B1(new_n528), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n541), .A2(G56), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n558), .B1(new_n561), .B2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  INV_X1    g142(.A(new_n528), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G53), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT9), .Z(new_n570));
  AOI22_X1  g145(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n571), .A2(new_n532), .B1(new_n526), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  OAI21_X1  g153(.A(G651), .B1(new_n541), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OR3_X1    g157(.A1(new_n526), .A2(KEYINPUT76), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT76), .B1(new_n526), .B2(new_n582), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n583), .A2(new_n584), .B1(G49), .B2(new_n568), .ZN(new_n585));
  OAI211_X1 g160(.A(KEYINPUT77), .B(G651), .C1(new_n541), .C2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(G288));
  AOI22_X1  g162(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT78), .B1(new_n588), .B2(new_n532), .ZN(new_n589));
  OAI21_X1  g164(.A(G61), .B1(new_n535), .B2(new_n536), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n592), .A2(new_n593), .A3(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n526), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G86), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n568), .A2(G48), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(G85), .A2(new_n596), .B1(new_n568), .B2(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n541), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n532), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n596), .A2(G92), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT10), .Z(new_n605));
  NAND2_X1  g180(.A1(new_n568), .A2(KEYINPUT79), .ZN(new_n606));
  INV_X1    g181(.A(G54), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n528), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n537), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n606), .A2(new_n609), .B1(G651), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n603), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n603), .B1(new_n615), .B2(G868), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n574), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n618), .B1(new_n574), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n615), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n615), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n481), .A2(new_n491), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT13), .Z(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n497), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n499), .A2(G123), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n465), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND3_X1  g213(.A1(new_n631), .A2(new_n632), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT80), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n654), .A3(G14), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT81), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT82), .Z(new_n659));
  NOR2_X1   g234(.A1(G2072), .A2(G2078), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n444), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(KEYINPUT17), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n662), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n657), .B(new_n658), .C1(new_n444), .C2(new_n660), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n659), .A3(new_n657), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2096), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n672), .A2(new_n677), .A3(new_n675), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n677), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n680));
  AOI211_X1 g255(.A(new_n676), .B(new_n678), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT23), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n574), .B2(new_n689), .ZN(new_n692));
  INV_X1    g267(.A(G1956), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(G19), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n562), .B2(new_n689), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(G1341), .Z(new_n697));
  INV_X1    g272(.A(G1961), .ZN(new_n698));
  NOR2_X1   g273(.A1(G171), .A2(new_n689), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G5), .B2(new_n689), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n694), .B(new_n697), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  AOI22_X1  g276(.A1(G129), .A2(new_n499), .B1(new_n497), .B2(G141), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT95), .B(KEYINPUT26), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G105), .B2(new_n481), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G32), .B(new_n707), .S(G29), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT27), .B(G1996), .Z(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G27), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G164), .B2(new_n710), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n708), .A2(new_n709), .B1(new_n712), .B2(G2078), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n700), .A2(new_n698), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n713), .B(new_n714), .C1(new_n708), .C2(new_n709), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n701), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT31), .B(G11), .Z(new_n717));
  NOR2_X1   g292(.A1(new_n637), .A2(new_n710), .ZN(new_n718));
  INV_X1    g293(.A(G28), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(KEYINPUT30), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT96), .Z(new_n721));
  AOI21_X1  g296(.A(G29), .B1(new_n719), .B2(KEYINPUT30), .ZN(new_n722));
  AOI211_X1 g297(.A(new_n717), .B(new_n718), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G1966), .ZN(new_n724));
  NOR2_X1   g299(.A1(G168), .A2(new_n689), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n689), .B2(G21), .ZN(new_n726));
  OAI221_X1 g301(.A(new_n723), .B1(G2078), .B2(new_n712), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n710), .A2(G33), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT25), .Z(new_n730));
  AOI22_X1  g305(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n465), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G139), .B2(new_n497), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n728), .B1(new_n733), .B2(new_n710), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(new_n442), .ZN(new_n735));
  INV_X1    g310(.A(new_n726), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G1966), .ZN(new_n737));
  NOR2_X1   g312(.A1(G4), .A2(G16), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT93), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n614), .B2(new_n689), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G1348), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n710), .A2(G26), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n497), .A2(G140), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n499), .A2(G128), .ZN(new_n745));
  OR2_X1    g320(.A1(G104), .A2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n746), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n744), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n743), .B1(new_n750), .B2(new_n710), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2067), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n727), .A2(new_n737), .A3(new_n741), .A4(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G2090), .ZN(new_n754));
  NOR2_X1   g329(.A1(G29), .A2(G35), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G162), .B2(G29), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT29), .Z(new_n757));
  OAI211_X1 g332(.A(new_n716), .B(new_n753), .C1(new_n754), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n754), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT24), .ZN(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G160), .B2(new_n710), .ZN(new_n764));
  INV_X1    g339(.A(G2084), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n770));
  INV_X1    g345(.A(G6), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G305), .B2(G16), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(KEYINPUT86), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT86), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT32), .B(G1981), .ZN(new_n778));
  AND3_X1   g353(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n775), .B2(new_n777), .ZN(new_n780));
  OR3_X1    g355(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT87), .ZN(new_n781));
  NOR2_X1   g356(.A1(G166), .A2(new_n689), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n689), .A2(G22), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OR3_X1    g359(.A1(new_n782), .A2(KEYINPUT90), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(KEYINPUT90), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G1971), .ZN(new_n788));
  INV_X1    g363(.A(G1971), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n785), .A2(new_n789), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n581), .A2(new_n585), .A3(G16), .A4(new_n586), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G23), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT88), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(KEYINPUT89), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT89), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n792), .A2(new_n797), .A3(new_n794), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT33), .B(G1976), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n800), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n796), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  AND3_X1   g378(.A1(new_n791), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(KEYINPUT87), .B1(new_n779), .B2(new_n780), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n781), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT34), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT34), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n781), .A2(new_n804), .A3(new_n808), .A4(new_n805), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G24), .ZN(new_n810));
  XOR2_X1   g385(.A(G290), .B(KEYINPUT85), .Z(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G16), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G1986), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n497), .A2(G131), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n499), .A2(G119), .ZN(new_n815));
  OR2_X1    g390(.A1(G95), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT84), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n814), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  MUX2_X1   g394(.A(G25), .B(new_n819), .S(G29), .Z(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n807), .A2(new_n809), .A3(new_n813), .A4(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n770), .A2(KEYINPUT36), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n770), .B(KEYINPUT36), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n770), .A2(KEYINPUT36), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n769), .B1(new_n828), .B2(new_n832), .ZN(G311));
  NAND2_X1  g408(.A1(new_n828), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(new_n768), .ZN(G150));
  AOI22_X1  g410(.A1(new_n541), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(new_n532), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n526), .A2(new_n838), .B1(new_n528), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT37), .ZN(new_n844));
  INV_X1    g419(.A(new_n841), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n562), .B1(new_n845), .B2(KEYINPUT98), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n841), .A2(new_n847), .A3(new_n562), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n615), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n842), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n844), .B1(new_n856), .B2(new_n857), .ZN(G145));
  NAND2_X1  g433(.A1(new_n497), .A2(G142), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n499), .A2(G130), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n465), .A2(G118), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT103), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n628), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n819), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n750), .B(new_n707), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n511), .A2(new_n491), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n514), .A2(KEYINPUT99), .A3(new_n521), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT99), .B1(new_n514), .B2(new_n521), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT100), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n870), .B(new_n875), .C1(new_n871), .C2(new_n872), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n877), .A2(KEYINPUT101), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(KEYINPUT101), .ZN(new_n879));
  OR3_X1    g454(.A1(new_n867), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n733), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT102), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n867), .B1(new_n878), .B2(new_n879), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n881), .A2(KEYINPUT102), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n880), .A2(new_n887), .A3(new_n882), .A4(new_n883), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n866), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n866), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n494), .B(new_n637), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n889), .B2(new_n890), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g472(.A1(new_n574), .A2(new_n614), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n574), .A2(new_n614), .A3(KEYINPUT104), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n574), .A2(new_n614), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(KEYINPUT105), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(KEYINPUT105), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n851), .B(new_n623), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n902), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n903), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n900), .A2(KEYINPUT106), .A3(new_n901), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  INV_X1    g490(.A(new_n902), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n903), .A2(new_n915), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n914), .A2(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n909), .B1(new_n908), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n920));
  XNOR2_X1  g495(.A(G288), .B(G290), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  XNOR2_X1  g499(.A(G166), .B(KEYINPUT107), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(G305), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n924), .A2(new_n926), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n909), .B(new_n931), .C1(new_n908), .C2(new_n918), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n920), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n930), .B1(new_n920), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(G868), .B2(new_n841), .ZN(G295));
  OAI21_X1  g511(.A(new_n935), .B1(G868), .B2(new_n841), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  XNOR2_X1  g513(.A(G171), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(G286), .ZN(new_n940));
  XNOR2_X1  g515(.A(G171), .B(KEYINPUT110), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(G168), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n943), .A2(new_n851), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n940), .A2(new_n942), .B1(new_n849), .B2(new_n850), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n916), .A2(new_n912), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n943), .A2(new_n851), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(new_n945), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n918), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n930), .B1(new_n951), .B2(KEYINPUT111), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n948), .B(new_n953), .C1(new_n918), .C2(new_n950), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n948), .B(new_n930), .C1(new_n918), .C2(new_n950), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n950), .A2(new_n905), .A3(new_n906), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n911), .A2(new_n913), .A3(new_n917), .ZN(new_n961));
  OAI221_X1 g536(.A(new_n961), .B1(new_n904), .B2(KEYINPUT41), .C1(new_n949), .C2(new_n945), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n962), .A3(new_n929), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(new_n894), .A3(new_n957), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n959), .B1(new_n964), .B2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(new_n965), .ZN(new_n966));
  AND4_X1   g541(.A1(new_n956), .A2(new_n963), .A3(new_n894), .A4(new_n957), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n951), .A2(KEYINPUT111), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n929), .A3(new_n954), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(new_n894), .A3(new_n957), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n967), .B1(new_n970), .B2(KEYINPUT43), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(G397));
  INV_X1    g548(.A(G1976), .ZN(new_n974));
  OR2_X1    g549(.A1(G288), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT99), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n522), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n514), .A2(KEYINPUT99), .A3(new_n521), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n512), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT113), .B1(new_n979), .B2(G1384), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n873), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n493), .A2(G40), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n487), .A2(new_n489), .A3(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(G8), .B(new_n975), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT52), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n980), .A2(new_n983), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n989), .A2(new_n487), .A3(new_n489), .A4(new_n985), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT52), .B1(G288), .B2(new_n974), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(G8), .A3(new_n975), .A4(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT114), .B(G86), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n526), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n595), .A2(new_n598), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G1981), .ZN(new_n996));
  INV_X1    g571(.A(G1981), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n595), .A2(new_n997), .A3(new_n597), .A4(new_n598), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT49), .B1(new_n996), .B2(new_n998), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(new_n990), .A3(G8), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n988), .A2(new_n992), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G303), .A2(G8), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT55), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n980), .A2(new_n1007), .A3(new_n983), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n870), .A2(new_n514), .A3(new_n521), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1009), .A2(KEYINPUT50), .A3(new_n982), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n487), .A2(new_n754), .A3(new_n489), .A4(new_n985), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n874), .A2(KEYINPUT45), .A3(new_n982), .A4(new_n876), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(G164), .B2(G1384), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n487), .A2(new_n489), .A3(new_n985), .A4(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n789), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g595(.A(new_n1004), .B(new_n1006), .C1(new_n1014), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1003), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n990), .A2(G8), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT115), .Z(new_n1024));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n1025));
  INV_X1    g600(.A(new_n998), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G288), .A2(G1976), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n1002), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1024), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1028), .A2(new_n1025), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1022), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1006), .ZN(new_n1032));
  INV_X1    g607(.A(new_n986), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n980), .A2(KEYINPUT50), .A3(new_n983), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1007), .B(new_n982), .C1(new_n512), .C2(new_n522), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1033), .A2(new_n754), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1020), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1032), .B1(new_n1039), .B2(G8), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n988), .A2(new_n992), .A3(new_n1002), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1040), .A2(new_n1021), .A3(new_n1041), .ZN(new_n1042));
  AND4_X1   g617(.A1(new_n487), .A2(new_n489), .A3(new_n985), .A4(new_n1018), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n443), .A3(new_n1015), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1011), .A2(new_n1033), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n698), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1009), .A2(KEYINPUT45), .A3(new_n982), .ZN(new_n1049));
  AND4_X1   g624(.A1(new_n487), .A2(new_n489), .A3(new_n1049), .A4(new_n985), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n980), .A2(new_n1017), .A3(new_n983), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1045), .A2(G2078), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1046), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT125), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1054), .A2(new_n1055), .A3(G171), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n1054), .B2(G171), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1042), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G168), .A2(new_n1004), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT51), .B1(new_n1060), .B2(KEYINPUT124), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1051), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n487), .A2(new_n1049), .A3(new_n489), .A4(new_n985), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n724), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n487), .A2(new_n765), .A3(new_n489), .A4(new_n985), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1011), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(G8), .B(new_n1062), .C1(new_n1069), .C2(G286), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1966), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1066), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1072));
  OAI21_X1  g647(.A(G8), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1060), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(new_n1074), .A3(new_n1061), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1069), .A2(new_n1060), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1059), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1058), .A2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1070), .A2(new_n1075), .B1(new_n1069), .B2(new_n1060), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1059), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1031), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1069), .A2(G8), .A3(G168), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT63), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1083), .A2(new_n1021), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1971), .B1(new_n1043), .B2(new_n1015), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1012), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1087));
  OAI21_X1  g662(.A(G8), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1006), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1003), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n1003), .B2(new_n1089), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1085), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(KEYINPUT119), .B(new_n1085), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1096));
  OR3_X1    g671(.A1(new_n1040), .A2(new_n1021), .A3(new_n1041), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1084), .B1(new_n1097), .B2(new_n1083), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1037), .A2(new_n487), .A3(new_n489), .A4(new_n985), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1034), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n693), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT56), .B(G2072), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1043), .A2(new_n1015), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n574), .A2(KEYINPUT120), .A3(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1105), .A2(KEYINPUT120), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(KEYINPUT120), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1107), .B(new_n1108), .C1(new_n570), .C2(new_n573), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1102), .A2(new_n1104), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1035), .B(KEYINPUT117), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n986), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(G1956), .B1(new_n1115), .B2(new_n1034), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1043), .A2(new_n1015), .A3(new_n1103), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1110), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT121), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1111), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(G1348), .B1(new_n1011), .B2(new_n1033), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n990), .A2(G2067), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n615), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1113), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1119), .A2(new_n1122), .A3(KEYINPUT61), .A4(new_n1112), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n615), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1124), .A2(new_n1125), .A3(new_n1129), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1016), .A2(new_n1019), .A3(G1996), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT58), .B(G1341), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1033), .B2(new_n989), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n562), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT59), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1139), .B(new_n562), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1138), .A2(new_n1140), .B1(new_n1132), .B2(new_n614), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1128), .A2(new_n1133), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT61), .B1(new_n1120), .B2(KEYINPUT122), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1118), .A2(new_n1144), .A3(new_n1112), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1127), .B1(new_n1142), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n874), .A2(new_n982), .A3(new_n876), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1017), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1033), .A2(new_n1152), .A3(new_n1015), .A4(new_n1052), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1156));
  AOI21_X1  g731(.A(G301), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT54), .B1(new_n1054), .B2(G171), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1042), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1159), .A2(new_n1080), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1057), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1054), .A2(new_n1055), .A3(G171), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1155), .A2(new_n1156), .A3(G301), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1082), .B(new_n1099), .C1(new_n1150), .C2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1152), .A2(new_n986), .ZN(new_n1169));
  INV_X1    g744(.A(new_n821), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n819), .B(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT112), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n707), .B(G1996), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n749), .B(G2067), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(G290), .B(G1986), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1169), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1168), .A2(new_n1178), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1152), .A2(new_n986), .A3(G1996), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT46), .Z(new_n1181));
  OAI21_X1  g756(.A(new_n1169), .B1(new_n707), .B2(new_n1174), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT47), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n819), .A2(new_n1170), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1175), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(G2067), .B2(new_n749), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1169), .ZN(new_n1188));
  NOR2_X1   g763(.A1(G290), .A2(G1986), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1169), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT127), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT48), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1176), .A2(new_n1169), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1191), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1194), .B1(new_n1195), .B2(KEYINPUT48), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1184), .B(new_n1188), .C1(new_n1193), .C2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1179), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(G319), .ZN(new_n1201));
  NOR4_X1   g775(.A1(G229), .A2(G401), .A3(new_n1201), .A4(G227), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n896), .A2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g777(.A1(new_n971), .A2(new_n1203), .ZN(G308));
  AOI21_X1  g778(.A(new_n956), .B1(new_n955), .B2(new_n957), .ZN(new_n1205));
  OAI211_X1 g779(.A(new_n896), .B(new_n1202), .C1(new_n1205), .C2(new_n967), .ZN(G225));
endmodule


