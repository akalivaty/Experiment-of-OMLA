//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n212), .B1(new_n215), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT64), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n220), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n202), .A2(G68), .ZN(new_n242));
  INV_X1    g0042(.A(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n241), .B(new_n247), .Z(G351));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n207), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI22_X1  g0053(.A1(new_n249), .A2(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(G20), .B2(new_n203), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n213), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n257), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n206), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G50), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(new_n266), .B1(new_n202), .B2(new_n262), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT66), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n270), .A2(new_n274), .A3(new_n271), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G226), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n206), .A2(G274), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT65), .B(G45), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(G41), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G222), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G223), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n286), .C1(G77), .C2(new_n281), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n277), .A2(new_n280), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n268), .B(new_n290), .C1(G179), .C2(new_n288), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n260), .A2(KEYINPUT9), .A3(new_n267), .ZN(new_n293));
  INV_X1    g0093(.A(new_n288), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G190), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(G200), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  INV_X1    g0097(.A(new_n267), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(new_n259), .B2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n293), .A2(new_n295), .A3(new_n296), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n299), .A2(new_n296), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n302), .A2(new_n303), .A3(new_n293), .A4(new_n295), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n292), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n281), .A2(G238), .A3(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G107), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n281), .A2(new_n283), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n306), .B1(new_n307), .B2(new_n281), .C1(new_n308), .C2(new_n220), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n286), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n276), .A2(G244), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n280), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(G200), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT15), .B(G87), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n316), .A2(new_n250), .ZN(new_n317));
  INV_X1    g0117(.A(G77), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT68), .B1(new_n207), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT68), .ZN(new_n321));
  XOR2_X1   g0121(.A(new_n249), .B(KEYINPUT67), .Z(new_n322));
  OAI221_X1 g0122(.A(new_n320), .B1(new_n321), .B2(new_n317), .C1(new_n322), .C2(new_n253), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n257), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n318), .B1(new_n206), .B2(G20), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n263), .A2(new_n325), .B1(new_n318), .B2(new_n262), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n314), .A2(new_n315), .A3(new_n324), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n326), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n312), .A2(G179), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n312), .A2(new_n289), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n305), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G33), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n334), .A2(new_n336), .A3(G226), .A4(G1698), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT73), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n281), .A2(KEYINPUT73), .A3(G226), .A4(G1698), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n334), .A2(new_n336), .A3(G223), .A4(new_n283), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G87), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n270), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n280), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(G169), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n348), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n344), .B1(new_n339), .B2(new_n340), .ZN(new_n351));
  OAI211_X1 g0151(.A(G179), .B(new_n350), .C1(new_n351), .C2(new_n270), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n249), .B1(new_n206), .B2(G20), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n263), .B1(new_n262), .B2(new_n249), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n219), .A2(new_n243), .ZN(new_n357));
  OAI21_X1  g0157(.A(G20), .B1(new_n357), .B2(new_n201), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n252), .A2(G159), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n281), .B2(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n334), .A2(new_n336), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n360), .B1(new_n365), .B2(G68), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n258), .B1(new_n366), .B2(KEYINPUT16), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT72), .B1(new_n335), .B2(G33), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(new_n333), .A3(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n371), .A3(new_n336), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n361), .A2(G20), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n243), .B1(new_n374), .B2(new_n362), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n368), .B1(new_n375), .B2(new_n360), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n356), .B1(new_n367), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT18), .B1(new_n353), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT7), .B1(new_n363), .B2(new_n207), .ZN(new_n379));
  AOI211_X1 g0179(.A(new_n361), .B(G20), .C1(new_n334), .C2(new_n336), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n360), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n376), .A2(new_n257), .A3(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(G190), .B(new_n350), .C1(new_n351), .C2(new_n270), .ZN(new_n385));
  OAI21_X1  g0185(.A(G200), .B1(new_n346), .B2(new_n348), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n384), .A2(new_n355), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT17), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n386), .A2(new_n385), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(new_n377), .A3(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n383), .A2(new_n257), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n374), .A2(new_n362), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G68), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT16), .B1(new_n394), .B2(new_n382), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n355), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n349), .A2(new_n352), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n378), .A2(new_n389), .A3(new_n391), .A4(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n332), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n262), .A2(new_n243), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT12), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n243), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n318), .B2(new_n250), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n263), .A2(G68), .A3(new_n264), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT11), .B1(new_n405), .B2(new_n257), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT14), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT69), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n270), .A2(new_n274), .A3(new_n271), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n274), .B1(new_n270), .B2(new_n271), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n273), .A2(KEYINPUT69), .A3(new_n275), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(G238), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n280), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT70), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(KEYINPUT70), .A3(new_n280), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G97), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n220), .A2(G1698), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G226), .B2(G1698), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n425), .B1(new_n427), .B2(new_n363), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n286), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n413), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n419), .A2(KEYINPUT70), .A3(new_n280), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT70), .B1(new_n419), .B2(new_n280), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n413), .B(new_n429), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n412), .B(G169), .C1(new_n430), .C2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT13), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(G179), .A3(new_n433), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n433), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n412), .B1(new_n440), .B2(G169), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n411), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n430), .A2(new_n434), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n411), .B1(new_n443), .B2(G190), .ZN(new_n444));
  INV_X1    g0244(.A(G200), .ZN(new_n445));
  AOI211_X1 g0245(.A(KEYINPUT71), .B(new_n445), .C1(new_n437), .C2(new_n433), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT71), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n447), .B1(new_n440), .B2(G200), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n444), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n401), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1), .ZN(new_n452));
  NAND2_X1  g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n270), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT75), .B1(new_n457), .B2(new_n222), .ZN(new_n458));
  OR2_X1    g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n453), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(G274), .A3(new_n452), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT75), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n456), .A2(new_n462), .A3(G257), .A4(new_n270), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n334), .A2(new_n336), .A3(G244), .A4(new_n283), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n283), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n281), .A2(G250), .A3(G1698), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n467), .A2(new_n468), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n464), .A2(KEYINPUT76), .B1(new_n286), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT77), .ZN(new_n473));
  INV_X1    g0273(.A(G179), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT76), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n458), .A2(new_n475), .A3(new_n461), .A4(new_n463), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n286), .B1(new_n452), .B2(new_n460), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n462), .B1(new_n478), .B2(G257), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n463), .A2(new_n461), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT76), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n471), .A2(new_n286), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n481), .A2(new_n476), .A3(new_n474), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT77), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(new_n476), .A3(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n393), .A2(G107), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  AND2_X1   g0288(.A1(G97), .A2(G107), .ZN(new_n489));
  NOR2_X1   g0289(.A1(G97), .A2(G107), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n307), .A2(KEYINPUT6), .A3(G97), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n207), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n253), .A2(new_n318), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT74), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT74), .ZN(new_n496));
  INV_X1    g0296(.A(new_n494), .ZN(new_n497));
  INV_X1    g0297(.A(new_n492), .ZN(new_n498));
  XNOR2_X1  g0298(.A(G97), .B(G107), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n498), .B1(new_n488), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n496), .B(new_n497), .C1(new_n500), .C2(new_n207), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n487), .A2(new_n495), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n257), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n261), .A2(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n206), .A2(G33), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n261), .A2(new_n505), .A3(new_n213), .A4(new_n256), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n504), .B1(new_n507), .B2(G97), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n289), .A2(new_n486), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n481), .A2(new_n476), .A3(G190), .A4(new_n482), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n510), .A2(new_n503), .A3(new_n508), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n486), .A2(G200), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n485), .A2(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n456), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n478), .A2(G270), .B1(new_n515), .B2(G274), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n334), .A2(new_n336), .A3(G264), .A4(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n334), .A2(new_n336), .A3(G257), .A4(new_n283), .ZN(new_n518));
  INV_X1    g0318(.A(G303), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n517), .B(new_n518), .C1(new_n519), .C2(new_n281), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n286), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n507), .A2(G116), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n262), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n256), .A2(new_n213), .B1(G20), .B2(new_n524), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n469), .B(new_n207), .C1(G33), .C2(new_n221), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n526), .A2(KEYINPUT20), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT20), .B1(new_n526), .B2(new_n527), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n523), .B(new_n525), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n522), .A2(G169), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT80), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(KEYINPUT21), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n530), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n516), .A2(new_n521), .A3(G190), .ZN(new_n536));
  INV_X1    g0336(.A(G270), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n461), .B1(new_n457), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n286), .B2(new_n520), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n535), .B(new_n536), .C1(new_n539), .C2(new_n445), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(G179), .A3(new_n530), .ZN(new_n541));
  INV_X1    g0341(.A(new_n533), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n522), .A2(new_n530), .A3(G169), .A4(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n534), .A2(new_n540), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n334), .A2(new_n336), .A3(G244), .A4(G1698), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n334), .A2(new_n336), .A3(G238), .A4(new_n283), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n545), .B(new_n546), .C1(new_n333), .C2(new_n524), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n286), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n278), .A2(G45), .ZN(new_n549));
  OAI21_X1  g0349(.A(G250), .B1(new_n451), .B2(G1), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n286), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n207), .B1(new_n425), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n490), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n334), .A2(new_n336), .A3(new_n207), .A4(G68), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n555), .B1(new_n250), .B2(new_n221), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT78), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n258), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT78), .A4(new_n561), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n564), .A2(new_n565), .B1(new_n262), .B2(new_n316), .ZN(new_n566));
  OR3_X1    g0366(.A1(new_n506), .A2(KEYINPUT79), .A3(new_n557), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT79), .B1(new_n506), .B2(new_n557), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n551), .B1(new_n547), .B2(new_n286), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G190), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n554), .A2(new_n566), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n562), .A2(new_n563), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(new_n257), .A3(new_n565), .ZN(new_n574));
  INV_X1    g0374(.A(new_n316), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n507), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n316), .A2(new_n262), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n553), .A2(new_n289), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n570), .A2(new_n474), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n572), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n544), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n262), .A2(KEYINPUT25), .A3(new_n307), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT83), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT25), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n261), .B2(G107), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n585), .B(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n307), .B2(new_n506), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n334), .A2(new_n336), .A3(new_n207), .A4(G87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT22), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n281), .A2(new_n592), .A3(new_n207), .A4(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n307), .A2(G20), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(KEYINPUT23), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(KEYINPUT23), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT81), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n594), .A2(new_n595), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n595), .B1(new_n594), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n257), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT82), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(KEYINPUT82), .B(new_n257), .C1(new_n604), .C2(new_n605), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n589), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n456), .A2(G264), .A3(new_n270), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT84), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n478), .A2(KEYINPUT84), .A3(G264), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n281), .A2(G257), .A3(G1698), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n281), .A2(G250), .A3(new_n283), .ZN(new_n616));
  INV_X1    g0416(.A(G294), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n615), .B(new_n616), .C1(new_n333), .C2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n613), .A2(new_n614), .B1(new_n618), .B2(new_n286), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n619), .A2(new_n461), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n286), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(new_n461), .A3(new_n611), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n620), .A2(G200), .B1(G190), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n610), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n620), .A2(G179), .B1(G169), .B2(new_n622), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n583), .B(new_n624), .C1(new_n625), .C2(new_n610), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n450), .A2(new_n514), .A3(new_n626), .ZN(G372));
  AND3_X1   g0427(.A1(new_n396), .A2(new_n398), .A3(new_n397), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n398), .B1(new_n396), .B2(new_n397), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n331), .ZN(new_n631));
  OAI21_X1  g0431(.A(G169), .B1(new_n430), .B2(new_n434), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n438), .A3(new_n435), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n449), .A2(new_n631), .B1(new_n634), .B2(new_n411), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n389), .A2(new_n391), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n630), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n301), .A2(new_n304), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n292), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n566), .A2(new_n576), .B1(new_n474), .B2(new_n570), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n547), .A2(KEYINPUT85), .A3(new_n286), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT85), .B1(new_n547), .B2(new_n286), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n552), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n289), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n571), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n574), .A2(new_n577), .A3(new_n569), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(G200), .B2(new_n644), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT86), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT85), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n548), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n547), .A2(KEYINPUT85), .A3(new_n286), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n445), .B1(new_n656), .B2(new_n552), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT86), .B1(new_n657), .B2(new_n649), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n647), .B1(new_n652), .B2(new_n658), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n534), .A2(new_n541), .A3(new_n543), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n610), .B2(new_n625), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n659), .A2(new_n513), .A3(new_n624), .A4(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n485), .A2(new_n509), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT26), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n572), .A2(new_n581), .ZN(new_n666));
  AND4_X1   g0466(.A1(KEYINPUT26), .A2(new_n666), .A3(new_n485), .A4(new_n509), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n646), .B(new_n662), .C1(new_n665), .C2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n640), .B1(new_n450), .B2(new_n669), .ZN(G369));
  NAND3_X1  g0470(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G343), .ZN(new_n675));
  XOR2_X1   g0475(.A(new_n675), .B(KEYINPUT87), .Z(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n535), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n544), .B2(KEYINPUT88), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(KEYINPUT88), .B2(new_n544), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n660), .A2(new_n677), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT89), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(KEYINPUT89), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n610), .A2(new_n623), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n610), .A2(new_n625), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n610), .B2(new_n676), .ZN(new_n690));
  INV_X1    g0490(.A(new_n688), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n676), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n688), .A2(new_n676), .ZN(new_n694));
  INV_X1    g0494(.A(new_n676), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n660), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n689), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n693), .A2(new_n694), .A3(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n210), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n558), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n217), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n662), .A2(new_n646), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n644), .A2(G200), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n651), .A3(new_n566), .A4(new_n569), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n658), .A2(new_n709), .A3(new_n571), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n485), .A3(new_n509), .A4(new_n646), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT26), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n667), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n676), .B1(new_n707), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT93), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n668), .A2(KEYINPUT93), .A3(new_n676), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n662), .A2(new_n646), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n666), .A2(new_n485), .A3(new_n509), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n712), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT94), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n659), .A2(new_n664), .A3(KEYINPUT26), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT94), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(new_n725), .A3(new_n712), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n695), .B1(new_n720), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n719), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT92), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n614), .A2(new_n613), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n621), .A3(new_n570), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n733), .A2(new_n474), .A3(new_n522), .ZN(new_n734));
  INV_X1    g0534(.A(new_n486), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(KEYINPUT30), .ZN(new_n736));
  XOR2_X1   g0536(.A(KEYINPUT90), .B(KEYINPUT30), .Z(new_n737));
  NAND4_X1  g0537(.A1(new_n619), .A2(new_n539), .A3(G179), .A4(new_n570), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n737), .B1(new_n738), .B2(new_n486), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n539), .A2(G179), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n619), .A2(new_n461), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n486), .A2(new_n740), .A3(new_n741), .A4(new_n644), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n736), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n695), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT91), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n739), .B2(new_n742), .ZN(new_n748));
  INV_X1    g0548(.A(new_n736), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n739), .A2(new_n747), .A3(new_n742), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n676), .A2(new_n745), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n731), .B(new_n746), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n754), .B1(new_n750), .B2(new_n751), .ZN(new_n756));
  AOI21_X1  g0556(.A(KEYINPUT31), .B1(new_n743), .B2(new_n695), .ZN(new_n757));
  OAI21_X1  g0557(.A(KEYINPUT92), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n689), .A2(new_n513), .A3(new_n583), .A4(new_n676), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G330), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n730), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n706), .B1(new_n763), .B2(G1), .ZN(G364));
  AND2_X1   g0564(.A1(new_n207), .A2(G13), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n206), .B1(new_n765), .B2(G45), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n701), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n210), .A2(G355), .A3(new_n281), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n700), .A2(new_n281), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n217), .B2(new_n279), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n247), .A2(new_n451), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n770), .B1(G116), .B2(new_n210), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n213), .B1(G20), .B2(new_n289), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n769), .B1(new_n774), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n207), .A2(new_n474), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n782), .A2(G190), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n782), .A2(new_n445), .A3(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  OAI221_X1 g0588(.A(new_n363), .B1(new_n784), .B2(new_n785), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G179), .A2(G200), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n790), .A2(G20), .A3(new_n313), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT96), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n789), .B1(G329), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n781), .A2(G190), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n445), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G326), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n207), .A2(new_n445), .A3(G179), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G190), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n800), .A2(new_n801), .B1(new_n519), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n798), .A2(G200), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(G322), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n802), .A2(new_n313), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT97), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT97), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n207), .B1(new_n790), .B2(G190), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n811), .A2(G283), .B1(G294), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g0617(.A1(new_n797), .A2(new_n806), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G159), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n795), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT32), .Z(new_n821));
  AOI22_X1  g0621(.A1(G68), .A2(new_n786), .B1(new_n783), .B2(G77), .ZN(new_n822));
  INV_X1    g0622(.A(new_n805), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n823), .A2(KEYINPUT95), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(KEYINPUT95), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n822), .B1(new_n202), .B2(new_n800), .C1(new_n826), .C2(new_n219), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n821), .B(new_n827), .C1(G97), .C2(new_n816), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n811), .A2(G107), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(new_n281), .C1(new_n557), .C2(new_n803), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT98), .Z(new_n831));
  AOI21_X1  g0631(.A(new_n818), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n778), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n780), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n681), .B2(new_n777), .ZN(new_n835));
  INV_X1    g0635(.A(new_n686), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n768), .B1(new_n681), .B2(new_n682), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G396));
  NAND2_X1  g0639(.A1(new_n695), .A2(new_n328), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n327), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n331), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n631), .A2(new_n676), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n716), .A2(new_n718), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n845), .A2(KEYINPUT100), .ZN(new_n846));
  INV_X1    g0646(.A(new_n844), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n676), .B(new_n847), .C1(new_n707), .C2(new_n713), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n845), .B2(KEYINPUT100), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n761), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT101), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n768), .B1(new_n850), .B2(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT101), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n854), .B(new_n761), .C1(new_n846), .C2(new_n849), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n778), .A2(new_n775), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n769), .B1(new_n318), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G283), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n363), .B1(new_n784), .B2(new_n524), .C1(new_n859), .C2(new_n787), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n810), .A2(new_n557), .B1(new_n221), .B2(new_n815), .ZN(new_n861));
  INV_X1    g0661(.A(new_n803), .ZN(new_n862));
  AOI22_X1  g0662(.A1(G107), .A2(new_n862), .B1(new_n805), .B2(G294), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n519), .B2(new_n800), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n795), .A2(new_n785), .ZN(new_n865));
  NOR4_X1   g0665(.A1(new_n860), .A2(new_n861), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G150), .A2(new_n786), .B1(new_n783), .B2(G159), .ZN(new_n867));
  INV_X1    g0667(.A(G137), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(new_n800), .ZN(new_n869));
  INV_X1    g0669(.A(new_n826), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n870), .B2(G143), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n871), .A2(KEYINPUT34), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n811), .A2(G68), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n816), .A2(G58), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n796), .A2(G132), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n363), .B1(new_n862), .B2(G50), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n873), .A2(new_n874), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n871), .B2(KEYINPUT34), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n866), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n858), .B1(new_n833), .B2(new_n879), .C1(new_n847), .C2(new_n776), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n856), .A2(new_n880), .ZN(G384));
  INV_X1    g0681(.A(new_n500), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n524), .B(new_n215), .C1(new_n882), .C2(KEYINPUT35), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(KEYINPUT35), .B2(new_n882), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT36), .Z(new_n885));
  OR3_X1    g0685(.A1(new_n217), .A2(new_n318), .A3(new_n357), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n206), .B(G13), .C1(new_n886), .C2(new_n242), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n387), .B1(new_n353), .B2(new_n377), .ZN(new_n889));
  INV_X1    g0689(.A(new_n674), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n377), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n396), .A2(new_n397), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n396), .A2(new_n674), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n387), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n400), .A2(new_n891), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n243), .B1(new_n362), .B2(new_n364), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n368), .B1(new_n901), .B2(new_n360), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n383), .A2(new_n902), .A3(new_n257), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n355), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(KEYINPUT102), .A3(new_n355), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n674), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n400), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n896), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n349), .A2(new_n352), .A3(new_n890), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n895), .B1(new_n913), .B2(new_n387), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n910), .B(KEYINPUT38), .C1(new_n911), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n900), .A2(new_n915), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n744), .A2(new_n745), .B1(new_n743), .B2(new_n753), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n844), .B1(new_n759), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n695), .A2(new_n411), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n442), .A2(new_n449), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(new_n442), .B2(new_n449), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n916), .B(new_n918), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n626), .A2(new_n514), .A3(new_n695), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n743), .A2(new_n753), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n746), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n847), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n410), .B1(new_n440), .B2(new_n313), .ZN(new_n927));
  OAI21_X1  g0727(.A(G200), .B1(new_n430), .B2(new_n434), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT71), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n440), .A2(new_n447), .A3(G200), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n411), .B(new_n695), .C1(new_n931), .C2(new_n634), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n442), .A2(new_n449), .A3(new_n919), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n926), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT38), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n914), .A2(new_n911), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n908), .B1(new_n636), .B2(new_n630), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT40), .B1(new_n938), .B2(new_n915), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n922), .A2(KEYINPUT40), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT105), .ZN(new_n941));
  INV_X1    g0741(.A(new_n450), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n923), .B2(new_n925), .ZN(new_n943));
  OAI21_X1  g0743(.A(G330), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n941), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT103), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n938), .A2(KEYINPUT39), .A3(new_n915), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n634), .A2(new_n411), .A3(new_n676), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n913), .A2(new_n387), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT37), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n951), .A2(new_n896), .B1(new_n400), .B2(new_n909), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n899), .B1(KEYINPUT38), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n947), .B(new_n949), .C1(new_n953), .C2(KEYINPUT39), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n890), .B1(new_n628), .B2(new_n629), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n848), .A2(new_n843), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n932), .A2(new_n933), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n938), .A2(new_n915), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n946), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n960), .A2(new_n946), .A3(new_n955), .A4(new_n954), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT104), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n450), .B1(new_n728), .B2(KEYINPUT29), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n719), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n965), .B1(new_n719), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n640), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n964), .B(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n945), .A2(new_n971), .B1(new_n206), .B2(new_n765), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n945), .A2(new_n971), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n888), .B1(new_n972), .B2(new_n973), .ZN(G367));
  INV_X1    g0774(.A(new_n771), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n233), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n779), .B1(new_n210), .B2(new_n316), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n768), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n281), .B1(new_n786), .B2(G294), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n785), .B2(new_n800), .C1(new_n859), .C2(new_n784), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(new_n870), .B2(G303), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n811), .A2(G97), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(new_n307), .C2(new_n815), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n862), .A2(KEYINPUT46), .A3(G116), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT46), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n803), .B2(new_n524), .ZN(new_n986));
  INV_X1    g0786(.A(G317), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n984), .B(new_n986), .C1(new_n987), .C2(new_n795), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n281), .B1(new_n784), .B2(new_n202), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G159), .B2(new_n786), .ZN(new_n990));
  INV_X1    g0790(.A(G143), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n800), .A2(new_n991), .B1(new_n219), .B2(new_n803), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G150), .B2(new_n805), .ZN(new_n993));
  XNOR2_X1  g0793(.A(KEYINPUT112), .B(G137), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n990), .B(new_n993), .C1(new_n795), .C2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n816), .A2(G68), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n318), .B2(new_n810), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n983), .A2(new_n988), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT47), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n978), .B1(new_n999), .B2(new_n778), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT113), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n695), .A2(new_n649), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(new_n646), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT106), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n659), .A2(new_n1002), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1001), .B1(new_n777), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n698), .A2(new_n694), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n503), .A2(new_n508), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(new_n676), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n513), .A2(new_n1012), .B1(new_n664), .B2(new_n695), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT44), .Z(new_n1015));
  NOR2_X1   g0815(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT45), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(new_n693), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n693), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(KEYINPUT109), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1018), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n693), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(KEYINPUT109), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT110), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n692), .A2(new_n697), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n698), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1027), .B1(new_n1030), .B2(new_n686), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n836), .A2(KEYINPUT110), .A3(new_n1029), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(KEYINPUT111), .A3(new_n686), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT111), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n836), .B2(new_n1029), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1031), .A2(new_n1032), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n763), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1026), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n763), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n701), .B(KEYINPUT41), .Z(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n767), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(KEYINPUT42), .B1(new_n1013), .B2(new_n698), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n511), .A2(new_n512), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n664), .B1(new_n1045), .B2(new_n688), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n695), .B2(new_n1046), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1013), .A2(new_n698), .A3(KEYINPUT42), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT107), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1006), .B(KEYINPUT43), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n693), .A2(new_n1013), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT43), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1050), .A2(new_n1054), .A3(new_n1007), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT108), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n693), .B2(new_n1013), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1056), .A2(KEYINPUT108), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1009), .B1(new_n1043), .B2(new_n1061), .ZN(G387));
  OAI211_X1 g0862(.A(new_n690), .B(new_n777), .C1(new_n691), .C2(new_n676), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G303), .A2(new_n783), .B1(new_n786), .B2(G311), .ZN(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT115), .B(G322), .Z(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n800), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n870), .B2(G317), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT48), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(KEYINPUT48), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n816), .A2(G283), .B1(G294), .B2(new_n862), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT49), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n363), .B1(new_n795), .B2(new_n801), .C1(new_n810), .C2(new_n524), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n281), .B1(new_n784), .B2(new_n243), .C1(new_n249), .C2(new_n787), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G150), .B2(new_n796), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n803), .A2(new_n318), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n800), .A2(new_n819), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(G50), .C2(new_n805), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n816), .A2(new_n575), .ZN(new_n1082));
  AND4_X1   g0882(.A1(new_n982), .A2(new_n1078), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n778), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n779), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n210), .A2(new_n281), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1086), .A2(new_n703), .B1(G107), .B2(new_n210), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n322), .A2(G50), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n703), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n975), .B1(new_n237), .B2(new_n279), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1087), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1084), .B(new_n768), .C1(new_n1085), .C2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT116), .Z(new_n1096));
  AOI22_X1  g0896(.A1(new_n1036), .A2(new_n767), .B1(new_n1063), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1037), .A2(new_n701), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1036), .A2(new_n763), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(G393));
  AOI21_X1  g0900(.A(new_n702), .B1(new_n1026), .B2(new_n1038), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1019), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n1020), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1037), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G150), .A2(new_n799), .B1(new_n805), .B2(G159), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT51), .Z(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n318), .B2(new_n815), .C1(new_n557), .C2(new_n810), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n281), .B1(new_n787), .B2(new_n202), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G68), .B2(new_n862), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n991), .B2(new_n795), .C1(new_n322), .C2(new_n784), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n363), .B1(new_n784), .B2(new_n617), .C1(new_n519), .C2(new_n787), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G283), .B2(new_n862), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n795), .A2(new_n1065), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n816), .A2(G116), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1113), .A2(new_n829), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G311), .A2(new_n805), .B1(new_n799), .B2(G317), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT52), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1108), .A2(new_n1111), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n778), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n771), .A2(new_n241), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1085), .B1(G97), .B2(new_n700), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n769), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n1013), .B2(new_n777), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1103), .B2(new_n766), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1105), .A2(new_n1128), .ZN(G390));
  NAND2_X1  g0929(.A1(new_n934), .A2(G330), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n760), .A2(G330), .A3(new_n847), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n958), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n676), .B(new_n842), .C1(new_n1133), .C2(new_n707), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n843), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n682), .B1(new_n759), .B2(new_n917), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n844), .B1(new_n1136), .B2(KEYINPUT117), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(KEYINPUT117), .B2(new_n1136), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n958), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1135), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1131), .A2(new_n958), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n957), .A2(new_n1132), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n942), .A2(new_n1136), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n640), .B(new_n1144), .C1(new_n967), .C2(new_n968), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1130), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n938), .A2(KEYINPUT39), .A3(new_n915), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT39), .B1(new_n900), .B2(new_n915), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n957), .A2(new_n958), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1151), .B1(new_n1152), .B2(new_n948), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n916), .A2(new_n948), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n1135), .B2(new_n958), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1148), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1135), .A2(new_n958), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n953), .A2(new_n949), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n843), .A2(new_n848), .B1(new_n932), .B2(new_n933), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1160), .A2(new_n949), .B1(new_n1150), .B2(new_n1149), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1161), .A3(new_n1141), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1156), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1147), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1163), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n1146), .A3(new_n1143), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n701), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n767), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n363), .B1(new_n784), .B2(new_n221), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G107), .B2(new_n786), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n800), .A2(new_n859), .B1(new_n557), .B2(new_n803), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G116), .B2(new_n805), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(new_n617), .C2(new_n795), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n873), .B1(new_n318), .B2(new_n815), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n281), .B1(new_n787), .B2(new_n994), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G128), .B2(new_n799), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT54), .B(G143), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT118), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n796), .A2(G125), .B1(new_n783), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(G132), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1176), .B(new_n1179), .C1(new_n1180), .C2(new_n823), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n803), .A2(new_n251), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT53), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n202), .B2(new_n810), .C1(new_n819), .C2(new_n815), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1173), .A2(new_n1174), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n778), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n769), .B1(new_n249), .B2(new_n857), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n1151), .C2(new_n776), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1168), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT119), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT119), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1168), .A2(new_n1191), .A3(new_n1188), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1167), .A2(new_n1190), .A3(new_n1192), .ZN(G378));
  INV_X1    g0993(.A(new_n857), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n768), .B1(G50), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n281), .A2(G41), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n784), .B2(new_n316), .C1(new_n221), .C2(new_n787), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G283), .B2(new_n796), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n800), .A2(new_n524), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1079), .B(new_n1199), .C1(G107), .C2(new_n805), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n811), .A2(G58), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1198), .A2(new_n996), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT58), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1196), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1205), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n799), .A2(G125), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n787), .B2(new_n1180), .C1(new_n868), .C2(new_n784), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G150), .B2(new_n816), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1178), .A2(new_n862), .B1(G128), .B2(new_n805), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT120), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT121), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n811), .A2(G159), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G33), .B(G41), .C1(new_n796), .C2(G124), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1207), .B1(new_n1203), .B2(new_n1202), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1195), .B1(new_n1221), .B2(new_n778), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n268), .A2(new_n674), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n305), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n305), .A2(new_n1223), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OR3_X1    g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1228), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n775), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1222), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1232), .B1(new_n940), .B2(new_n682), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT40), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n934), .B2(new_n916), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n958), .A2(new_n918), .A3(new_n939), .ZN(new_n1239));
  OAI211_X1 g1039(.A(G330), .B(new_n1231), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1236), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n964), .A3(KEYINPUT122), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n954), .A2(new_n955), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT103), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(KEYINPUT122), .A3(new_n962), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n1236), .A3(new_n1240), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1242), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1235), .B1(new_n1248), .B2(new_n767), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT57), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1241), .B(new_n1246), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1146), .B1(new_n1163), .B2(new_n1142), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1250), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1241), .A2(new_n964), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1245), .A2(new_n962), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n1236), .A3(new_n1240), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1250), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n702), .B1(new_n1258), .B2(new_n1252), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT123), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1254), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  AOI211_X1 g1061(.A(KEYINPUT123), .B(new_n702), .C1(new_n1258), .C2(new_n1252), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1249), .B1(new_n1261), .B2(new_n1262), .ZN(G375));
  NAND2_X1  g1063(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1147), .A2(new_n1042), .A3(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n768), .B1(G68), .B2(new_n1194), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n281), .B1(new_n784), .B2(new_n251), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G159), .B2(new_n862), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n796), .A2(G128), .B1(new_n786), .B2(new_n1178), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(new_n1180), .C2(new_n800), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1201), .B1(new_n202), .B2(new_n815), .C1(new_n826), .C2(new_n994), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n823), .A2(new_n859), .B1(new_n800), .B2(new_n617), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G97), .B2(new_n862), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n363), .B1(new_n784), .B2(new_n307), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G116), .B2(new_n786), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1273), .B(new_n1275), .C1(new_n519), .C2(new_n795), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1082), .B1(new_n318), .B2(new_n810), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n1270), .A2(new_n1271), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1266), .B1(new_n1278), .B2(new_n778), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n958), .B2(new_n776), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1142), .B2(new_n766), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1265), .A2(new_n1282), .ZN(G381));
  NAND2_X1  g1083(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n766), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1061), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1008), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(G390), .A2(new_n1289), .A3(G384), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1189), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1167), .A2(new_n1292), .ZN(new_n1293));
  OR4_X1    g1093(.A1(G375), .A2(new_n1291), .A3(G381), .A4(new_n1293), .ZN(G407));
  INV_X1    g1094(.A(new_n1249), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT57), .B1(new_n1248), .B2(new_n1252), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1257), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1256), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1252), .B(KEYINPUT57), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n701), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1296), .B1(new_n1300), .B2(KEYINPUT123), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1295), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1293), .ZN(new_n1304));
  INV_X1    g1104(.A(G343), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(G213), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1303), .A2(new_n1304), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(G407), .A2(G213), .A3(new_n1308), .ZN(G409));
  AOI21_X1  g1109(.A(new_n1127), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G393), .A2(G396), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1310), .B1(new_n1312), .B2(new_n1288), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(G390), .A2(new_n1289), .A3(new_n1311), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1287), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1313), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(G387), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1317), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G378), .B(new_n1249), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1248), .A2(new_n1042), .A3(new_n1252), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1235), .B1(new_n1321), .B2(new_n767), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1304), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1319), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1142), .A2(KEYINPUT60), .A3(new_n1145), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1326), .A2(new_n701), .ZN(new_n1327));
  OAI21_X1  g1127(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1264), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1281), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT124), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n856), .A2(new_n1331), .A3(new_n880), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n856), .A2(new_n1331), .A3(new_n880), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1331), .B1(new_n856), .B2(new_n880), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1333), .B1(new_n1330), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1325), .A2(new_n1306), .A3(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(KEYINPUT62), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT126), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT61), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1307), .B1(new_n1319), .B2(new_n1324), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1307), .A2(G2897), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1337), .A2(new_n1345), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1333), .B(new_n1344), .C1(new_n1330), .C2(new_n1336), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  OAI211_X1 g1148(.A(new_n1341), .B(new_n1342), .C1(new_n1343), .C2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT62), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1343), .A2(new_n1350), .A3(new_n1338), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1340), .A2(new_n1349), .A3(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1347), .ZN(new_n1353));
  AND2_X1   g1153(.A1(new_n1327), .A2(new_n1329), .ZN(new_n1354));
  OAI22_X1  g1154(.A1(new_n1354), .A2(new_n1281), .B1(new_n1335), .B2(new_n1334), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1344), .B1(new_n1355), .B2(new_n1333), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1353), .A2(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1293), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1358), .B1(new_n1303), .B2(G378), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1357), .B1(new_n1359), .B2(new_n1307), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1341), .B1(new_n1360), .B2(new_n1342), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1318), .B1(new_n1352), .B2(new_n1361), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1318), .A2(KEYINPUT61), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT125), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1357), .A2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1348), .A2(KEYINPUT125), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n1365), .B(new_n1366), .C1(new_n1307), .C2(new_n1359), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1343), .A2(KEYINPUT63), .A3(new_n1338), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT63), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1339), .A2(new_n1369), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1363), .A2(new_n1367), .A3(new_n1368), .A4(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1362), .A2(new_n1371), .ZN(G405));
  NAND3_X1  g1172(.A1(new_n1315), .A2(new_n1317), .A3(KEYINPUT127), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(G375), .A2(new_n1304), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1374), .A2(new_n1319), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1375), .A2(new_n1338), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1374), .A2(new_n1319), .A3(new_n1337), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1373), .A2(new_n1376), .A3(new_n1377), .ZN(new_n1378));
  AOI21_X1  g1178(.A(KEYINPUT127), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1379));
  XNOR2_X1  g1179(.A(new_n1378), .B(new_n1379), .ZN(G402));
endmodule


