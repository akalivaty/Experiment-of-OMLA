//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT69), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n462), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n464), .A2(new_n466), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n462), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n464), .A2(new_n466), .A3(new_n462), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT70), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(new_n462), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT72), .Z(new_n489));
  NAND3_X1  g064(.A1(new_n478), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n481), .A2(new_n498), .A3(G138), .A4(new_n462), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n505), .B1(new_n502), .B2(G543), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(G543), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT74), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n502), .A2(G543), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n504), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT73), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n518));
  OAI211_X1 g093(.A(G62), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n512), .B1(new_n515), .B2(new_n523), .ZN(G166));
  NAND2_X1  g099(.A1(new_n503), .A2(new_n505), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(new_n516), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT75), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n506), .A2(new_n529), .A3(G63), .A4(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n511), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n507), .A2(KEYINPUT76), .A3(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n506), .A2(new_n507), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  AND4_X1   g115(.A1(new_n531), .A2(new_n536), .A3(new_n538), .A4(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(new_n535), .A2(G52), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n506), .A2(G90), .A3(new_n507), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n542), .A2(KEYINPUT78), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT78), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n533), .B2(new_n534), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n548), .B2(new_n543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n526), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n514), .B1(new_n553), .B2(KEYINPUT77), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n554), .B1(KEYINPUT77), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  AOI22_X1  g132(.A1(new_n535), .A2(G43), .B1(new_n537), .B2(G81), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n514), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(G860), .A3(new_n560), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n526), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n507), .A2(G53), .A3(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n537), .A2(G91), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(G299));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(new_n511), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n537), .A2(G88), .B1(G50), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n522), .B1(new_n521), .B2(G651), .ZN(new_n578));
  AOI211_X1 g153(.A(KEYINPUT74), .B(new_n514), .C1(new_n519), .C2(new_n520), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(G303));
  OAI21_X1  g155(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n506), .A2(G87), .A3(new_n507), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n507), .A2(G49), .A3(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT79), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n581), .A2(new_n582), .A3(new_n586), .A4(new_n583), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G288));
  NAND3_X1  g164(.A1(new_n525), .A2(G61), .A3(new_n516), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n514), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n525), .A2(G86), .A3(new_n516), .A4(new_n507), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n507), .A2(G48), .A3(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n535), .A2(G47), .B1(new_n537), .B2(G85), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n514), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n526), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(G54), .A2(new_n535), .B1(new_n604), .B2(G651), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n506), .A2(G92), .A3(new_n507), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT80), .B1(new_n610), .B2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  MUX2_X1   g187(.A(KEYINPUT80), .B(new_n611), .S(new_n612), .Z(G284));
  MUX2_X1   g188(.A(KEYINPUT80), .B(new_n611), .S(new_n612), .Z(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n610), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n610), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(KEYINPUT81), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(KEYINPUT81), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n558), .A2(new_n560), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n615), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g203(.A1(new_n479), .A2(new_n463), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2100), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n485), .A2(G135), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n462), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n475), .A2(G123), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT82), .B(G2096), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n632), .A2(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT84), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n645), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n662), .B(KEYINPUT17), .Z(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n659), .B2(new_n660), .ZN(new_n667));
  INV_X1    g242(.A(new_n659), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(new_n662), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n661), .B1(new_n669), .B2(new_n660), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n665), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT86), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  MUX2_X1   g261(.A(new_n686), .B(new_n685), .S(new_n678), .Z(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G20), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT23), .ZN(new_n697));
  INV_X1    g272(.A(G299), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n695), .ZN(new_n699));
  INV_X1    g274(.A(G1956), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G35), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G162), .B2(new_n702), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT29), .Z(new_n705));
  INV_X1    g280(.A(G2090), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n701), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT97), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n702), .A2(G33), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n480), .A2(new_n483), .A3(G139), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(G115), .A2(G2104), .ZN(new_n712));
  INV_X1    g287(.A(G127), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n474), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G2105), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT25), .Z(new_n717));
  NAND4_X1  g292(.A1(new_n711), .A2(KEYINPUT92), .A3(new_n715), .A4(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n715), .A2(new_n717), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n710), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n709), .B1(new_n723), .B2(new_n702), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G2072), .ZN(new_n725));
  NOR2_X1   g300(.A1(G4), .A2(G16), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n610), .B2(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n725), .B1(G1348), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G1348), .B2(new_n727), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n724), .A2(G2072), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n695), .A2(G5), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G171), .B2(new_n695), .ZN(new_n733));
  INV_X1    g308(.A(G1961), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n729), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n702), .A2(G32), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT26), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n481), .A2(G129), .A3(G2105), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n480), .A2(new_n483), .A3(G141), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n737), .B1(new_n745), .B2(new_n702), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT27), .B(G1996), .Z(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT94), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n746), .B(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT30), .B(G28), .ZN(new_n750));
  OR2_X1    g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  NAND2_X1  g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n750), .A2(new_n702), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n638), .B2(new_n702), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT95), .Z(new_n755));
  MUX2_X1   g330(.A(G19), .B(new_n625), .S(G16), .Z(new_n756));
  XOR2_X1   g331(.A(KEYINPUT91), .B(G1341), .Z(new_n757));
  AOI211_X1 g332(.A(new_n749), .B(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n705), .A2(new_n706), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n702), .A2(G26), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT28), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n480), .A2(new_n483), .A3(G140), .ZN(new_n762));
  OR2_X1    g337(.A1(G104), .A2(G2105), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n763), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n464), .A2(new_n466), .A3(G128), .A4(G2105), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n761), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2067), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n756), .B2(new_n757), .ZN(new_n770));
  NAND2_X1  g345(.A1(G164), .A2(G29), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G27), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT96), .B(G2078), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  AND2_X1   g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n702), .B1(KEYINPUT24), .B2(G34), .ZN(new_n777));
  OAI22_X1  g352(.A1(G160), .A2(new_n702), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2084), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n770), .A2(new_n774), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n695), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n695), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n758), .A2(new_n759), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n708), .A2(new_n736), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G6), .A2(G16), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n596), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT32), .ZN(new_n789));
  INV_X1    g364(.A(G1981), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G23), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT88), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n584), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT88), .A4(new_n583), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n792), .B1(new_n797), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT33), .B(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G16), .A2(G22), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G166), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1971), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n791), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT89), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n805), .A2(KEYINPUT89), .A3(KEYINPUT34), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G24), .ZN(new_n810));
  XNOR2_X1  g385(.A(G290), .B(KEYINPUT87), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1986), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n702), .A2(G25), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n485), .A2(G131), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n462), .A2(G107), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n475), .A2(G119), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n814), .B1(new_n821), .B2(new_n702), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XOR2_X1   g398(.A(new_n822), .B(new_n823), .Z(new_n824));
  NOR3_X1   g399(.A1(new_n809), .A2(new_n813), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(KEYINPUT90), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n807), .A2(new_n808), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n807), .A2(new_n808), .A3(new_n825), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT90), .B(KEYINPUT36), .Z(new_n830));
  OAI211_X1 g405(.A(new_n786), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(G150));
  INV_X1    g406(.A(G150), .ZN(G311));
  NAND2_X1  g407(.A1(new_n610), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n535), .A2(G55), .B1(new_n537), .B2(G93), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(new_n514), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n625), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n558), .A2(new_n835), .A3(new_n560), .A4(new_n837), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n834), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n842), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n838), .A2(G860), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT98), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT99), .ZN(G145));
  NAND2_X1  g425(.A1(new_n485), .A2(G142), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n462), .A2(G118), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n475), .A2(G130), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n497), .A2(new_n499), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n493), .A2(new_n494), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n859), .A2(new_n762), .A3(new_n766), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n767), .A2(G164), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n745), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n745), .B1(new_n860), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n720), .A2(new_n710), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n860), .A2(new_n861), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n743), .A2(new_n744), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n722), .B1(new_n869), .B2(new_n862), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n856), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n820), .B(new_n630), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n723), .B1(new_n863), .B2(new_n864), .ZN(new_n873));
  INV_X1    g448(.A(new_n865), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n874), .A3(new_n862), .ZN(new_n875));
  INV_X1    g450(.A(new_n856), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n871), .A2(new_n872), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT100), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n872), .B1(new_n871), .B2(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(G160), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n638), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n871), .A2(new_n877), .ZN(new_n883));
  INV_X1    g458(.A(new_n872), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G160), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n885), .A2(KEYINPUT100), .A3(new_n886), .A4(new_n878), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n881), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n882), .B1(new_n881), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(G162), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n881), .A2(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n638), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n881), .A2(new_n882), .A3(new_n887), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n490), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n890), .A2(new_n894), .A3(new_n895), .A4(new_n897), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(G395));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n609), .A2(new_n698), .ZN(new_n903));
  AOI21_X1  g478(.A(G299), .B1(new_n608), .B2(new_n605), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT102), .B1(new_n609), .B2(new_n698), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(KEYINPUT41), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT103), .A4(KEYINPUT41), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n903), .A2(new_n904), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n909), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n841), .B(new_n621), .Z(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n905), .A2(new_n906), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n796), .A2(G290), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n796), .A2(G290), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT104), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n925), .A3(new_n922), .ZN(new_n926));
  XNOR2_X1  g501(.A(G303), .B(new_n596), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  OR3_X1    g503(.A1(new_n923), .A2(new_n927), .A3(KEYINPUT104), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n916), .A2(new_n931), .A3(new_n918), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n920), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n930), .B1(new_n920), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n838), .A2(new_n615), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n936), .ZN(G331));
  INV_X1    g513(.A(new_n930), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n550), .A2(G168), .A3(new_n555), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G168), .B1(new_n550), .B2(new_n555), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n841), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G301), .A2(G286), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n944), .A2(new_n839), .A3(new_n840), .A4(new_n940), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n917), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n943), .A2(new_n945), .A3(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(KEYINPUT105), .B(new_n841), .C1(new_n941), .C2(new_n942), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n939), .B(new_n949), .C1(new_n914), .C2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n905), .A2(new_n912), .A3(new_n906), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n946), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n930), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n954), .A2(new_n960), .A3(new_n895), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n951), .A2(new_n952), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n909), .A2(new_n910), .A3(new_n913), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n948), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(G37), .B1(new_n968), .B2(new_n939), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n949), .B1(new_n914), .B2(new_n953), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n930), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n964), .A2(KEYINPUT44), .A3(new_n965), .A4(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n972), .B1(new_n969), .B2(new_n971), .ZN(new_n976));
  AND4_X1   g551(.A1(new_n972), .A2(new_n954), .A3(new_n960), .A4(new_n895), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n978), .ZN(G397));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n980));
  INV_X1    g555(.A(G8), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(G166), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n469), .A2(new_n472), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(G1384), .B1(new_n857), .B2(new_n858), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n988), .B2(KEYINPUT45), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT107), .B(G1384), .ZN(new_n991));
  NOR3_X1   g566(.A1(G164), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n803), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT115), .B1(new_n988), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n988), .A2(new_n995), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n988), .A2(KEYINPUT115), .A3(new_n995), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n987), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G2090), .B1(new_n1000), .B2(KEYINPUT116), .ZN(new_n1001));
  INV_X1    g576(.A(new_n472), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n467), .A2(new_n468), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G2105), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1004), .A3(G40), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n996), .B2(new_n997), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n999), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n994), .B1(new_n1001), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n985), .B1(new_n1009), .B2(new_n981), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n1011));
  NOR3_X1   g586(.A1(G166), .A2(new_n980), .A3(new_n981), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT108), .B1(new_n988), .B2(new_n995), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1005), .B1(new_n988), .B2(new_n995), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1017), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n706), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n981), .B1(new_n1019), .B2(new_n993), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n982), .A2(KEYINPUT109), .A3(new_n983), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1014), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1014), .A2(new_n1020), .A3(KEYINPUT110), .A4(new_n1021), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n794), .A2(G1976), .A3(new_n795), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n981), .B1(new_n988), .B2(new_n987), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n585), .A2(new_n1032), .A3(new_n587), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1033), .A2(new_n1027), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1030), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n590), .A2(new_n591), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G651), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n593), .A2(new_n594), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n790), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n592), .B2(new_n595), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT49), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n988), .A2(new_n987), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT111), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n790), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n592), .A2(new_n595), .A3(G1981), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AND4_X1   g625(.A1(KEYINPUT111), .A2(new_n1050), .A3(new_n1045), .A4(new_n1029), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1035), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n536), .A2(new_n540), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1054), .A2(G8), .A3(new_n531), .A4(new_n538), .ZN(new_n1055));
  INV_X1    g630(.A(G2084), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1015), .A2(new_n1016), .A3(new_n1056), .A4(new_n1018), .ZN(new_n1057));
  NOR3_X1   g632(.A1(G164), .A2(new_n990), .A3(G1384), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n783), .B1(new_n989), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1010), .A2(new_n1026), .A3(new_n1053), .A4(new_n1060), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1060), .B(KEYINPUT63), .C1(new_n1020), .C2(new_n984), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1064), .B(new_n1052), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1039), .B(KEYINPUT113), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1050), .A2(new_n1045), .A3(new_n1029), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT111), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1044), .A2(KEYINPUT111), .A3(new_n1045), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n588), .A2(new_n1032), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1069), .B(new_n1071), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT114), .B1(new_n1080), .B2(new_n1070), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1029), .B(KEYINPUT112), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1053), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1067), .A2(new_n1068), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1065), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT118), .B1(new_n1088), .B2(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1000), .A2(new_n700), .ZN(new_n1090));
  INV_X1    g665(.A(new_n989), .ZN(new_n1091));
  INV_X1    g666(.A(new_n991), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n859), .A2(KEYINPUT45), .A3(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(G299), .B(KEYINPUT57), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1090), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1956), .B1(new_n1006), .B2(new_n999), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1095), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1101), .A3(KEYINPUT61), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT121), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1098), .A2(new_n1101), .A3(new_n1104), .A4(KEYINPUT61), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n558), .A2(new_n560), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n990), .B1(G164), .B2(G1384), .ZN(new_n1109));
  INV_X1    g684(.A(G1996), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(new_n1093), .A3(new_n1110), .A4(new_n987), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(G1341), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1042), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1108), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1116), .B(new_n1108), .C1(new_n1111), .C2(new_n1114), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1121));
  INV_X1    g696(.A(G1348), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n1124));
  INV_X1    g699(.A(G2067), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n988), .A2(new_n1125), .A3(new_n987), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1123), .A2(new_n1124), .A3(new_n610), .A4(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n610), .A3(new_n1126), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT60), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n610), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1120), .B(new_n1127), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT61), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1106), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n609), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1098), .A2(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1136), .A2(new_n1101), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1121), .A2(new_n734), .ZN(new_n1139));
  INV_X1    g714(.A(G2078), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1058), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1091), .A2(KEYINPUT53), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1109), .A2(new_n1093), .A3(new_n1140), .A4(new_n987), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1139), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(G171), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT45), .B1(new_n859), .B2(new_n1092), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n472), .A2(KEYINPUT123), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n472), .A2(KEYINPUT123), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1140), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1152));
  NOR4_X1   g727(.A1(new_n1150), .A2(new_n1151), .A3(new_n469), .A4(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1149), .A2(new_n1093), .A3(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1139), .A2(G301), .A3(new_n1145), .A4(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1147), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT124), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n1159));
  AOI211_X1 g734(.A(new_n1159), .B(KEYINPUT54), .C1(new_n1147), .C2(new_n1155), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1139), .A2(new_n1145), .A3(new_n1154), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1157), .B1(new_n1162), .B2(G171), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(G171), .B2(new_n1146), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1010), .A2(new_n1026), .A3(new_n1164), .A4(new_n1053), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1057), .A2(new_n1059), .A3(G168), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(G8), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1168), .A2(KEYINPUT51), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n1170));
  AOI21_X1  g745(.A(G168), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT51), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1138), .A2(new_n1166), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1010), .A2(new_n1026), .A3(new_n1053), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1180), .A2(new_n1147), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1175), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1182), .A2(KEYINPUT62), .A3(new_n1173), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1179), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1087), .A2(new_n1089), .A3(new_n1177), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1148), .A2(new_n987), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  OR2_X1    g762(.A1(new_n821), .A2(new_n823), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n821), .A2(new_n823), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n767), .B(new_n1125), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n868), .B(new_n1110), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(G290), .B(G1986), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1187), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1185), .A2(new_n1194), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1187), .A2(KEYINPUT46), .A3(new_n1110), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT46), .B1(new_n1187), .B2(new_n1110), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1186), .B1(new_n1190), .B2(new_n745), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT47), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1192), .A2(new_n1187), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1186), .A2(G290), .A3(G1986), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT48), .Z(new_n1203));
  AOI21_X1  g778(.A(new_n1200), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1191), .A2(new_n1190), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1189), .B1(new_n1205), .B2(new_n1187), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n767), .A2(G2067), .ZN(new_n1207));
  OR3_X1    g782(.A1(new_n1206), .A2(KEYINPUT125), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(KEYINPUT125), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1208), .A2(new_n1187), .A3(new_n1209), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n1210), .A2(KEYINPUT126), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(KEYINPUT126), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1204), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1213), .B(KEYINPUT127), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1195), .A2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g790(.A(G319), .ZN(new_n1217));
  NOR4_X1   g791(.A1(G229), .A2(new_n1217), .A3(G401), .A4(G227), .ZN(new_n1218));
  OAI21_X1  g792(.A(new_n1218), .B1(new_n976), .B2(new_n977), .ZN(new_n1219));
  AND2_X1   g793(.A1(new_n894), .A2(new_n895), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n1219), .B1(new_n890), .B2(new_n1220), .ZN(G308));
  OAI211_X1 g795(.A(new_n896), .B(new_n1218), .C1(new_n976), .C2(new_n977), .ZN(G225));
endmodule


