//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  OR4_X1    g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  AND2_X1   g031(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n457));
  NOR2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  OAI22_X1  g041(.A1(new_n462), .A2(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n460), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n459), .A2(new_n461), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  MUX2_X1   g048(.A(G100), .B(G112), .S(G2105), .Z(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n459), .A2(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(G136), .B2(new_n477), .ZN(G162));
  OAI211_X1 g053(.A(G126), .B(G2105), .C1(new_n457), .C2(new_n458), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  OR2_X1    g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  MUX2_X1   g057(.A(G102), .B(G114), .S(G2105), .Z(new_n483));
  AOI22_X1  g058(.A1(new_n481), .A2(new_n482), .B1(G2104), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n461), .C1(new_n457), .C2(new_n458), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G164));
  INV_X1    g063(.A(G651), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT70), .B1(new_n489), .B2(KEYINPUT6), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G651), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(KEYINPUT6), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G88), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G50), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(new_n502), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  AND2_X1   g084(.A1(G75), .A2(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n501), .A2(new_n504), .A3(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  AND2_X1   g088(.A1(new_n494), .A2(new_n495), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(G89), .A3(new_n508), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(G51), .A3(G543), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT71), .B1(new_n497), .B2(new_n498), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n506), .A2(new_n518), .A3(new_n507), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n517), .A2(new_n519), .A3(G63), .A4(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  AND4_X1   g097(.A1(new_n515), .A2(new_n516), .A3(new_n520), .A4(new_n522), .ZN(G168));
  NAND2_X1  g098(.A1(new_n503), .A2(G52), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT72), .B(G90), .Z(new_n525));
  NAND2_X1  g100(.A1(new_n500), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n517), .A2(new_n519), .A3(G64), .ZN(new_n528));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n489), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(G171));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n517), .A2(new_n519), .A3(G56), .ZN(new_n533));
  NAND2_X1  g108(.A1(G68), .A2(G543), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n533), .A2(KEYINPUT73), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT73), .B1(new_n533), .B2(new_n534), .ZN(new_n536));
  NOR3_X1   g111(.A1(new_n535), .A2(new_n536), .A3(new_n489), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n514), .A2(G43), .A3(G543), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n514), .A2(G81), .A3(new_n508), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n532), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n536), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n533), .A2(KEYINPUT73), .A3(new_n534), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(G651), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n540), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT74), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND4_X1  g128(.A1(new_n494), .A2(G53), .A3(G543), .A4(new_n495), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n499), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n494), .A2(G91), .A3(new_n495), .A4(new_n508), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n555), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  NAND4_X1  g139(.A1(new_n515), .A2(new_n516), .A3(new_n520), .A4(new_n522), .ZN(G286));
  NAND4_X1  g140(.A1(new_n494), .A2(G49), .A3(G543), .A4(new_n495), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n494), .A2(G87), .A3(new_n495), .A4(new_n508), .ZN(new_n567));
  AOI21_X1  g142(.A(G74), .B1(new_n517), .B2(new_n519), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n489), .ZN(G288));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n514), .A2(new_n508), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n500), .A2(KEYINPUT76), .A3(G86), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT75), .B1(new_n499), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n508), .A2(new_n578), .A3(G61), .ZN(new_n579));
  INV_X1    g154(.A(G73), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n577), .B(new_n579), .C1(new_n580), .C2(new_n502), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n503), .B2(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n575), .A2(new_n582), .ZN(G305));
  NAND3_X1  g158(.A1(new_n517), .A2(new_n519), .A3(G60), .ZN(new_n584));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n589), .A3(G651), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT78), .B(G85), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(G47), .A2(new_n503), .B1(new_n500), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(G290));
  NAND4_X1  g170(.A1(new_n494), .A2(G92), .A3(new_n495), .A4(new_n508), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n489), .B1(new_n599), .B2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n503), .A2(G54), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n598), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g182(.A(new_n606), .B1(G868), .B2(G171), .ZN(G321));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  MUX2_X1   g184(.A(G286), .B(G299), .S(new_n609), .Z(G297));
  MUX2_X1   g185(.A(G286), .B(G299), .S(new_n609), .Z(G280));
  INV_X1    g186(.A(new_n605), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  OAI21_X1  g189(.A(KEYINPUT81), .B1(new_n547), .B2(G868), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n612), .A2(new_n616), .A3(new_n613), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT80), .B1(new_n605), .B2(G559), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  MUX2_X1   g195(.A(KEYINPUT81), .B(new_n615), .S(new_n620), .Z(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g197(.A1(new_n465), .A2(new_n459), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  MUX2_X1   g202(.A(G99), .B(G111), .S(G2105), .Z(new_n628));
  AOI22_X1  g203(.A1(new_n472), .A2(G123), .B1(G2104), .B2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G135), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n462), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT82), .Z(new_n632));
  INV_X1    g207(.A(G2096), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n627), .A2(new_n634), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2427), .ZN(new_n639));
  INV_X1    g214(.A(G2430), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n642), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT84), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  OR2_X1    g234(.A1(new_n654), .A2(new_n657), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n656), .B1(new_n660), .B2(KEYINPUT17), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n654), .B1(new_n663), .B2(new_n657), .ZN(new_n664));
  INV_X1    g239(.A(new_n657), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n664), .B1(new_n665), .B2(new_n662), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n659), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n633), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(G2100), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(G2100), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT87), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT86), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT20), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n673), .A2(new_n679), .A3(new_n675), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n673), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT88), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n681), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT89), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n690), .B(new_n694), .ZN(G229));
  MUX2_X1   g270(.A(G95), .B(G107), .S(G2105), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G2104), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT90), .Z(new_n698));
  AOI22_X1  g273(.A1(G119), .A2(new_n472), .B1(new_n477), .B2(G131), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G25), .B(new_n700), .S(G29), .Z(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G6), .B(G305), .S(G16), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G23), .ZN(new_n708));
  OR2_X1    g283(.A1(G288), .A2(KEYINPUT92), .ZN(new_n709));
  NAND2_X1  g284(.A1(G288), .A2(KEYINPUT92), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n708), .B1(new_n711), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT33), .B(G1976), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G16), .A2(G22), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G166), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n707), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n704), .B1(new_n719), .B2(KEYINPUT34), .ZN(new_n720));
  NOR2_X1   g295(.A1(G16), .A2(G24), .ZN(new_n721));
  INV_X1    g296(.A(G290), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G16), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT91), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1986), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n720), .B(new_n725), .C1(KEYINPUT34), .C2(new_n719), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT36), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT25), .ZN(new_n728));
  INV_X1    g303(.A(G103), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n464), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n477), .A2(G139), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n461), .B2(new_n733), .ZN(new_n734));
  MUX2_X1   g309(.A(G33), .B(new_n734), .S(G29), .Z(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G2072), .Z(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  NAND2_X1  g312(.A1(G160), .A2(G29), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  AND2_X1   g314(.A1(KEYINPUT24), .A2(G34), .ZN(new_n740));
  NOR2_X1   g315(.A1(KEYINPUT24), .A2(G34), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  AOI22_X1  g318(.A1(G129), .A2(new_n472), .B1(new_n477), .B2(G141), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT26), .Z(new_n746));
  INV_X1    g321(.A(G105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n746), .C1(new_n747), .C2(new_n465), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT95), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  MUX2_X1   g325(.A(G32), .B(new_n750), .S(G29), .Z(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT96), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n736), .B1(new_n737), .B2(new_n743), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT97), .ZN(new_n755));
  NOR2_X1   g330(.A1(G5), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G171), .B2(G16), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT100), .Z(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  NOR2_X1   g334(.A1(G16), .A2(G21), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G168), .B2(G16), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT98), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n758), .A2(new_n759), .B1(G1966), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G1966), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n751), .A2(new_n753), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n739), .A2(G27), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT101), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n487), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2078), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT29), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n765), .B(new_n769), .C1(G2090), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n739), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n477), .A2(G140), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n472), .A2(G128), .ZN(new_n777));
  MUX2_X1   g352(.A(G104), .B(G116), .S(G2105), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G2104), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(new_n739), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2067), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n743), .A2(new_n737), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT31), .B(G11), .Z(new_n785));
  XOR2_X1   g360(.A(KEYINPUT99), .B(G28), .Z(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT30), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n786), .B2(KEYINPUT30), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n784), .B(new_n789), .C1(new_n632), .C2(new_n739), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n773), .A2(new_n783), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G4), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n612), .B2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT93), .B(G1348), .Z(new_n794));
  XOR2_X1   g369(.A(new_n793), .B(new_n794), .Z(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n759), .B2(new_n758), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n755), .A2(new_n764), .A3(new_n791), .A4(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G16), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G19), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n547), .B2(new_n798), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT94), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1341), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n772), .A2(G2090), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n798), .A2(G20), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT23), .Z(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G299), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1956), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT102), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n797), .A2(new_n802), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n727), .A2(new_n810), .ZN(G150));
  INV_X1    g386(.A(G150), .ZN(G311));
  AOI22_X1  g387(.A1(G55), .A2(new_n503), .B1(new_n500), .B2(G93), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n517), .A2(new_n519), .A3(G67), .ZN(new_n814));
  AND2_X1   g389(.A1(G80), .A2(G543), .ZN(new_n815));
  OAI21_X1  g390(.A(G651), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G860), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n612), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n541), .A2(new_n546), .A3(new_n817), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n816), .B(new_n813), .C1(new_n537), .C2(new_n540), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n821), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT103), .Z(new_n827));
  INV_X1    g402(.A(G860), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n825), .B2(KEYINPUT39), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n819), .B1(new_n827), .B2(new_n829), .ZN(G145));
  MUX2_X1   g405(.A(G106), .B(G118), .S(G2105), .Z(new_n831));
  AOI22_X1  g406(.A1(new_n472), .A2(G130), .B1(G2104), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G142), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n462), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n625), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n700), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n750), .B(new_n780), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n487), .B(new_n734), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(G162), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n632), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  INV_X1    g422(.A(new_n845), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n841), .A2(new_n842), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n846), .A2(KEYINPUT104), .A3(new_n847), .A4(new_n849), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n852), .B2(new_n853), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(G395));
  INV_X1    g432(.A(KEYINPUT109), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT108), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(KEYINPUT42), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n709), .A2(new_n861), .A3(new_n710), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n709), .B2(new_n710), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n722), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n709), .A2(new_n710), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT106), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n709), .A2(new_n861), .A3(new_n710), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(G290), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G305), .B(G303), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT107), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT107), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n874), .A3(new_n870), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n871), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n859), .A2(KEYINPUT42), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n824), .B(new_n619), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n605), .A2(G299), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n601), .A2(new_n602), .B1(G54), .B2(new_n503), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n881), .A2(new_n562), .A3(new_n555), .A4(new_n598), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n824), .B(new_n619), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n880), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT41), .B1(new_n880), .B2(new_n882), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n878), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n876), .A2(new_n884), .A3(new_n877), .A4(new_n889), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n860), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n860), .A3(new_n892), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n609), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n817), .A2(G868), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n858), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n895), .ZN(new_n899));
  OAI21_X1  g474(.A(G868), .B1(new_n899), .B2(new_n893), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n900), .B(KEYINPUT109), .C1(G868), .C2(new_n817), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n898), .A2(new_n901), .ZN(G295));
  NOR2_X1   g477(.A1(new_n896), .A2(new_n897), .ZN(G331));
  AND2_X1   g478(.A1(new_n524), .A2(new_n526), .ZN(new_n904));
  INV_X1    g479(.A(new_n530), .ZN(new_n905));
  NAND3_X1  g480(.A1(G168), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(G286), .B1(new_n527), .B2(new_n530), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n822), .A2(new_n823), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n908), .B1(new_n822), .B2(new_n823), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n888), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n888), .B(KEYINPUT110), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT111), .ZN(new_n916));
  INV_X1    g491(.A(new_n908), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n824), .A2(KEYINPUT111), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n883), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n876), .ZN(new_n922));
  INV_X1    g497(.A(new_n871), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n869), .A2(new_n874), .A3(new_n870), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n874), .B1(new_n869), .B2(new_n870), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n915), .A2(new_n926), .A3(new_n920), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n847), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n824), .A2(new_n917), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n822), .A2(new_n823), .A3(new_n908), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(new_n888), .A3(new_n918), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n883), .A3(new_n933), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n876), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n927), .A2(new_n938), .A3(new_n847), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n930), .B1(new_n929), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n939), .A2(new_n943), .A3(KEYINPUT43), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(new_n939), .B2(KEYINPUT43), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT113), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT44), .B1(new_n928), .B2(KEYINPUT43), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT112), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n939), .A2(new_n943), .A3(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n922), .A2(new_n847), .A3(new_n927), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n941), .B1(new_n954), .B2(new_n929), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT113), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n942), .B1(new_n949), .B2(new_n956), .ZN(G397));
  NAND2_X1  g532(.A1(G160), .A2(G40), .ZN(new_n958));
  AOI21_X1  g533(.A(G1384), .B1(new_n484), .B2(new_n486), .ZN(new_n959));
  XOR2_X1   g534(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OR3_X1    g538(.A1(new_n963), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT46), .B1(new_n963), .B2(G1996), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n780), .B(G2067), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n750), .A2(new_n966), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n964), .A2(new_n965), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n962), .A2(new_n966), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT115), .Z(new_n971));
  XNOR2_X1  g546(.A(new_n750), .B(G1996), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n962), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n700), .A2(new_n703), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n780), .A2(G2067), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n963), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n702), .B1(new_n698), .B2(new_n699), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n962), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n973), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(G290), .A2(G1986), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n962), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT48), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n969), .B(new_n977), .C1(new_n980), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n581), .A2(G651), .ZN(new_n986));
  INV_X1    g561(.A(G48), .ZN(new_n987));
  INV_X1    g562(.A(new_n503), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n571), .A2(new_n572), .ZN(new_n990));
  OAI21_X1  g565(.A(G1981), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1981), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n575), .A2(new_n582), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n993), .A3(KEYINPUT49), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  INV_X1    g570(.A(G40), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n467), .A2(new_n470), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n995), .B1(new_n959), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n991), .A2(new_n993), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI211_X1 g578(.A(KEYINPUT118), .B(KEYINPUT49), .C1(new_n991), .C2(new_n993), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n999), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n998), .B1(new_n1006), .B2(new_n865), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT52), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n998), .B(new_n1009), .C1(new_n1006), .C2(new_n865), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1005), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G303), .A2(G8), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT55), .ZN(new_n1015));
  INV_X1    g590(.A(G1384), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n487), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n958), .B1(new_n1017), .B2(KEYINPUT50), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n959), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G2090), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n959), .A2(KEYINPUT117), .A3(new_n1019), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1018), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n997), .B1(new_n959), .B2(new_n961), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n717), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n995), .B(new_n1015), .C1(new_n1025), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1015), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1020), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n959), .A2(KEYINPUT119), .A3(new_n1019), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1018), .A2(new_n1033), .A3(new_n1023), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n1029), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1031), .B1(new_n1036), .B2(G8), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1013), .A2(new_n1030), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n997), .B1(new_n1017), .B2(new_n960), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n1042));
  OR4_X1    g617(.A1(new_n1040), .A2(new_n1041), .A3(G2078), .A4(new_n1042), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1040), .B1(new_n1044), .B2(G2078), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1018), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n759), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G171), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1018), .A2(new_n1022), .A3(new_n737), .A4(new_n1024), .ZN(new_n1051));
  INV_X1    g626(.A(G1966), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n995), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n1054), .B2(KEYINPUT125), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G168), .A2(new_n995), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G8), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1056), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(KEYINPUT125), .A3(KEYINPUT51), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1054), .A2(G286), .ZN(new_n1062));
  AND4_X1   g637(.A1(KEYINPUT62), .A2(new_n1057), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT62), .B1(new_n1064), .B2(new_n1057), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1050), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  OR4_X1    g641(.A1(new_n1040), .A2(new_n1027), .A3(new_n1028), .A4(G2078), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1045), .A2(new_n1067), .A3(G301), .A4(new_n1047), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1049), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT126), .B(KEYINPUT54), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1045), .A2(new_n1067), .A3(new_n1047), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(G171), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1043), .A2(new_n1045), .A3(G301), .A4(new_n1047), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1069), .A2(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1064), .A2(new_n1057), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT61), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1018), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G299), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT57), .ZN(new_n1082));
  XOR2_X1   g657(.A(new_n561), .B(KEYINPUT123), .Z(new_n1083));
  INV_X1    g658(.A(new_n555), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1082), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT56), .B(G2072), .Z(new_n1089));
  OR3_X1    g664(.A1(new_n1027), .A2(new_n1028), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1080), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1088), .B1(new_n1080), .B2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1077), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1080), .A2(new_n1090), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1088), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(KEYINPUT61), .A3(new_n1091), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1027), .A2(new_n1028), .A3(G1996), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1017), .A2(new_n958), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT58), .B(G1341), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n547), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT59), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n547), .B(new_n1105), .C1(new_n1099), .C2(new_n1102), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1017), .A2(new_n958), .A3(G2067), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1046), .B2(new_n794), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n605), .A2(KEYINPUT60), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1104), .A2(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1046), .A2(new_n794), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1107), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n605), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n612), .B(new_n1107), .C1(new_n1046), .C2(new_n794), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT60), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND4_X1   g690(.A1(new_n1094), .A2(new_n1098), .A3(new_n1110), .A4(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1091), .B1(new_n1093), .B2(new_n1113), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT124), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1119), .B(new_n1091), .C1(new_n1093), .C2(new_n1113), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1075), .B(new_n1076), .C1(new_n1116), .C2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1039), .B1(new_n1066), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n995), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1124), .A2(new_n1031), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1054), .A2(G168), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(KEYINPUT63), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1127), .A2(new_n1030), .A3(new_n1013), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT63), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT49), .B1(new_n991), .B2(new_n993), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(new_n1000), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1011), .B1(new_n1132), .B2(new_n999), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1037), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1124), .A2(new_n1031), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1126), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1130), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT120), .B1(new_n1038), .B2(new_n1126), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1129), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1038), .A2(KEYINPUT120), .A3(new_n1126), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1141), .A2(new_n1142), .A3(KEYINPUT121), .A4(new_n1130), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1128), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n993), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G288), .A2(G1976), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1005), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n998), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n1147), .A2(new_n1148), .B1(new_n1013), .B2(new_n1135), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1123), .A2(new_n1144), .A3(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(G290), .A2(G1986), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n962), .B1(new_n982), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n980), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT116), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n985), .B1(new_n1150), .B2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g730(.A1(new_n669), .A2(G319), .A3(new_n670), .ZN(new_n1157));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n1158));
  NOR2_X1   g732(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g733(.A1(new_n1159), .A2(G229), .A3(G401), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g736(.A(new_n1162), .B1(new_n852), .B2(new_n853), .ZN(new_n1163));
  AND2_X1   g737(.A1(new_n1163), .A2(new_n940), .ZN(G308));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n940), .ZN(G225));
endmodule


