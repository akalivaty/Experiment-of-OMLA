

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n640), .A2(n820), .ZN(n602) );
  NAND2_X1 U550 ( .A1(n699), .A2(n697), .ZN(n660) );
  NAND2_X1 U551 ( .A1(G8), .A2(n660), .ZN(n596) );
  XNOR2_X2 U552 ( .A(n516), .B(n515), .ZN(n531) );
  XNOR2_X2 U553 ( .A(KEYINPUT66), .B(G543), .ZN(n516) );
  NOR2_X1 U554 ( .A1(n650), .A2(n649), .ZN(n652) );
  NOR2_X2 U555 ( .A1(n553), .A2(n552), .ZN(G160) );
  XNOR2_X1 U556 ( .A(KEYINPUT90), .B(n700), .ZN(n513) );
  OR2_X1 U557 ( .A1(n745), .A2(n744), .ZN(n514) );
  INV_X1 U558 ( .A(KEYINPUT28), .ZN(n601) );
  INV_X1 U559 ( .A(KEYINPUT98), .ZN(n651) );
  INV_X1 U560 ( .A(KEYINPUT0), .ZN(n515) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n808) );
  AND2_X1 U562 ( .A1(n541), .A2(G2104), .ZN(n890) );
  XNOR2_X1 U563 ( .A(KEYINPUT64), .B(n519), .ZN(n812) );
  NOR2_X1 U564 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U565 ( .A(KEYINPUT72), .B(n530), .Z(G299) );
  NAND2_X1 U566 ( .A1(G91), .A2(n808), .ZN(n518) );
  INV_X1 U567 ( .A(G651), .ZN(n522) );
  NOR2_X1 U568 ( .A1(n522), .A2(n531), .ZN(n811) );
  NAND2_X1 U569 ( .A1(G78), .A2(n811), .ZN(n517) );
  NAND2_X1 U570 ( .A1(n518), .A2(n517), .ZN(n529) );
  NOR2_X1 U571 ( .A1(G651), .A2(n531), .ZN(n519) );
  NAND2_X1 U572 ( .A1(G53), .A2(n812), .ZN(n521) );
  INV_X1 U573 ( .A(KEYINPUT70), .ZN(n520) );
  XNOR2_X1 U574 ( .A(n521), .B(n520), .ZN(n526) );
  NOR2_X1 U575 ( .A1(G543), .A2(n522), .ZN(n523) );
  XOR2_X1 U576 ( .A(KEYINPUT1), .B(n523), .Z(n807) );
  NAND2_X1 U577 ( .A1(n807), .A2(G65), .ZN(n524) );
  XNOR2_X1 U578 ( .A(KEYINPUT69), .B(n524), .ZN(n525) );
  NOR2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U580 ( .A(n527), .B(KEYINPUT71), .ZN(n528) );
  NAND2_X1 U581 ( .A1(G87), .A2(n531), .ZN(n536) );
  NAND2_X1 U582 ( .A1(G651), .A2(G74), .ZN(n533) );
  NAND2_X1 U583 ( .A1(G49), .A2(n812), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U585 ( .A1(n807), .A2(n534), .ZN(n535) );
  NAND2_X1 U586 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U587 ( .A(KEYINPUT87), .B(n537), .Z(G288) );
  NOR2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n538) );
  XOR2_X1 U589 ( .A(KEYINPUT17), .B(n538), .Z(n889) );
  NAND2_X1 U590 ( .A1(G138), .A2(n889), .ZN(n540) );
  INV_X1 U591 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U592 ( .A1(G102), .A2(n890), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n545) );
  AND2_X1 U594 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U595 ( .A1(G114), .A2(n885), .ZN(n543) );
  NOR2_X1 U596 ( .A1(G2104), .A2(n541), .ZN(n886) );
  NAND2_X1 U597 ( .A1(G126), .A2(n886), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U599 ( .A1(n545), .A2(n544), .ZN(G164) );
  NAND2_X1 U600 ( .A1(G101), .A2(n890), .ZN(n546) );
  XNOR2_X1 U601 ( .A(n546), .B(KEYINPUT23), .ZN(n547) );
  XNOR2_X1 U602 ( .A(n547), .B(KEYINPUT65), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G113), .A2(n885), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U605 ( .A1(G125), .A2(n886), .ZN(n551) );
  NAND2_X1 U606 ( .A1(G137), .A2(n889), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G64), .A2(n807), .ZN(n554) );
  XNOR2_X1 U609 ( .A(n554), .B(KEYINPUT67), .ZN(n560) );
  NAND2_X1 U610 ( .A1(n808), .A2(G90), .ZN(n555) );
  XNOR2_X1 U611 ( .A(n555), .B(KEYINPUT68), .ZN(n557) );
  NAND2_X1 U612 ( .A1(G77), .A2(n811), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U614 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U616 ( .A1(G52), .A2(n812), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n562), .A2(n561), .ZN(G301) );
  XNOR2_X1 U618 ( .A(KEYINPUT7), .B(KEYINPUT80), .ZN(n574) );
  NAND2_X1 U619 ( .A1(n808), .A2(G89), .ZN(n563) );
  XNOR2_X1 U620 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G76), .A2(n811), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U623 ( .A(KEYINPUT5), .B(n566), .ZN(n572) );
  NAND2_X1 U624 ( .A1(n807), .A2(G63), .ZN(n567) );
  XOR2_X1 U625 ( .A(KEYINPUT79), .B(n567), .Z(n569) );
  NAND2_X1 U626 ( .A1(G51), .A2(n812), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U628 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U630 ( .A(n574), .B(n573), .ZN(G168) );
  NAND2_X1 U631 ( .A1(G62), .A2(n807), .ZN(n576) );
  NAND2_X1 U632 ( .A1(G50), .A2(n812), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U634 ( .A(KEYINPUT88), .B(n577), .Z(n581) );
  NAND2_X1 U635 ( .A1(G88), .A2(n808), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G75), .A2(n811), .ZN(n578) );
  AND2_X1 U637 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n581), .A2(n580), .ZN(G303) );
  INV_X1 U639 ( .A(G303), .ZN(G166) );
  XOR2_X1 U640 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U641 ( .A1(G61), .A2(n807), .ZN(n583) );
  NAND2_X1 U642 ( .A1(G86), .A2(n808), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U644 ( .A1(n811), .A2(G73), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT2), .B(n584), .Z(n585) );
  NOR2_X1 U646 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U647 ( .A1(G48), .A2(n812), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n588), .A2(n587), .ZN(G305) );
  NAND2_X1 U649 ( .A1(G60), .A2(n807), .ZN(n590) );
  NAND2_X1 U650 ( .A1(G85), .A2(n808), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U652 ( .A1(n811), .A2(G72), .ZN(n592) );
  NAND2_X1 U653 ( .A1(G47), .A2(n812), .ZN(n591) );
  NAND2_X1 U654 ( .A1(n592), .A2(n591), .ZN(n593) );
  OR2_X1 U655 ( .A1(n594), .A2(n593), .ZN(G290) );
  NOR2_X1 U656 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NOR2_X1 U657 ( .A1(G164), .A2(G1384), .ZN(n699) );
  NAND2_X1 U658 ( .A1(G40), .A2(G160), .ZN(n595) );
  XNOR2_X1 U659 ( .A(KEYINPUT89), .B(n595), .ZN(n697) );
  XOR2_X2 U660 ( .A(KEYINPUT95), .B(n596), .Z(n743) );
  INV_X1 U661 ( .A(n743), .ZN(n692) );
  NAND2_X1 U662 ( .A1(n687), .A2(n692), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n597), .A2(KEYINPUT33), .ZN(n695) );
  INV_X1 U664 ( .A(n660), .ZN(n646) );
  NAND2_X1 U665 ( .A1(n646), .A2(G2072), .ZN(n598) );
  XNOR2_X1 U666 ( .A(n598), .B(KEYINPUT27), .ZN(n600) );
  AND2_X1 U667 ( .A1(G1956), .A2(n660), .ZN(n599) );
  NOR2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n640) );
  INV_X1 U669 ( .A(G299), .ZN(n820) );
  XNOR2_X1 U670 ( .A(n602), .B(n601), .ZN(n644) );
  NAND2_X1 U671 ( .A1(n812), .A2(G54), .ZN(n610) );
  NAND2_X1 U672 ( .A1(G66), .A2(n807), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G92), .A2(n808), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U675 ( .A(KEYINPUT76), .B(n605), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n811), .A2(G79), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n606), .B(KEYINPUT77), .ZN(n607) );
  NOR2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(n612) );
  XOR2_X1 U680 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n611) );
  XNOR2_X2 U681 ( .A(n612), .B(n611), .ZN(n929) );
  NAND2_X1 U682 ( .A1(G1348), .A2(n660), .ZN(n614) );
  NAND2_X1 U683 ( .A1(G2067), .A2(n646), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U685 ( .A1(n929), .A2(n615), .ZN(n639) );
  XOR2_X1 U686 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n617) );
  NAND2_X1 U687 ( .A1(G56), .A2(n807), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n617), .B(n616), .ZN(n624) );
  NAND2_X1 U689 ( .A1(G81), .A2(n808), .ZN(n618) );
  XOR2_X1 U690 ( .A(KEYINPUT12), .B(n618), .Z(n619) );
  XNOR2_X1 U691 ( .A(n619), .B(KEYINPUT75), .ZN(n621) );
  NAND2_X1 U692 ( .A1(G68), .A2(n811), .ZN(n620) );
  NAND2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U694 ( .A(KEYINPUT13), .B(n622), .Z(n623) );
  NOR2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U696 ( .A1(G43), .A2(n812), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n921) );
  NAND2_X1 U698 ( .A1(n929), .A2(G1348), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n627), .A2(KEYINPUT26), .ZN(n628) );
  NOR2_X1 U700 ( .A1(G1341), .A2(n628), .ZN(n629) );
  NOR2_X1 U701 ( .A1(n646), .A2(n629), .ZN(n631) );
  NOR2_X1 U702 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n630) );
  NOR2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n636) );
  NAND2_X1 U704 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n929), .A2(G2067), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n646), .A2(n634), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U709 ( .A1(n921), .A2(n637), .ZN(n638) );
  NOR2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U711 ( .A1(n640), .A2(n820), .ZN(n641) );
  NAND2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n645), .B(KEYINPUT29), .ZN(n650) );
  XOR2_X1 U715 ( .A(G2078), .B(KEYINPUT25), .Z(n1012) );
  NOR2_X1 U716 ( .A1(n1012), .A2(n660), .ZN(n648) );
  NOR2_X1 U717 ( .A1(n646), .A2(G1961), .ZN(n647) );
  NOR2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n656) );
  NOR2_X1 U719 ( .A1(G301), .A2(n656), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n652), .B(n651), .ZN(n679) );
  NOR2_X1 U721 ( .A1(G1966), .A2(n743), .ZN(n680) );
  NOR2_X1 U722 ( .A1(G2084), .A2(n660), .ZN(n676) );
  NOR2_X1 U723 ( .A1(n680), .A2(n676), .ZN(n653) );
  NAND2_X1 U724 ( .A1(G8), .A2(n653), .ZN(n654) );
  XNOR2_X1 U725 ( .A(KEYINPUT30), .B(n654), .ZN(n655) );
  NOR2_X1 U726 ( .A1(G168), .A2(n655), .ZN(n658) );
  AND2_X1 U727 ( .A1(G301), .A2(n656), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U729 ( .A(KEYINPUT31), .B(n659), .Z(n678) );
  INV_X1 U730 ( .A(G8), .ZN(n666) );
  NOR2_X1 U731 ( .A1(G2090), .A2(n660), .ZN(n661) );
  XNOR2_X1 U732 ( .A(KEYINPUT99), .B(n661), .ZN(n664) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n743), .ZN(n662) );
  NOR2_X1 U734 ( .A1(G166), .A2(n662), .ZN(n663) );
  NAND2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  OR2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n668) );
  AND2_X1 U737 ( .A1(n678), .A2(n668), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n679), .A2(n667), .ZN(n672) );
  INV_X1 U739 ( .A(n668), .ZN(n670) );
  AND2_X1 U740 ( .A1(G286), .A2(G8), .ZN(n669) );
  OR2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n674) );
  XNOR2_X1 U743 ( .A(KEYINPUT100), .B(KEYINPUT32), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n674), .B(n673), .ZN(n735) );
  INV_X1 U745 ( .A(KEYINPUT33), .ZN(n675) );
  AND2_X1 U746 ( .A1(n735), .A2(n675), .ZN(n685) );
  NAND2_X1 U747 ( .A1(G8), .A2(n676), .ZN(n677) );
  XOR2_X1 U748 ( .A(KEYINPUT97), .B(n677), .Z(n683) );
  AND2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n681) );
  NOR2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n734) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n922) );
  AND2_X1 U753 ( .A1(n734), .A2(n922), .ZN(n684) );
  NAND2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n691) );
  INV_X1 U755 ( .A(n922), .ZN(n688) );
  NOR2_X1 U756 ( .A1(G1971), .A2(G303), .ZN(n686) );
  NOR2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n923) );
  OR2_X1 U758 ( .A1(n688), .A2(n923), .ZN(n689) );
  OR2_X1 U759 ( .A1(KEYINPUT33), .A2(n689), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n693) );
  NAND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U763 ( .A(KEYINPUT101), .B(n696), .Z(n732) );
  XOR2_X1 U764 ( .A(G1981), .B(G305), .Z(n939) );
  INV_X1 U765 ( .A(n697), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n761) );
  XNOR2_X1 U767 ( .A(G1986), .B(G290), .ZN(n928) );
  NAND2_X1 U768 ( .A1(n761), .A2(n928), .ZN(n700) );
  AND2_X1 U769 ( .A1(n939), .A2(n513), .ZN(n730) );
  XOR2_X1 U770 ( .A(KEYINPUT94), .B(KEYINPUT38), .Z(n702) );
  NAND2_X1 U771 ( .A1(G105), .A2(n890), .ZN(n701) );
  XNOR2_X1 U772 ( .A(n702), .B(n701), .ZN(n706) );
  NAND2_X1 U773 ( .A1(G117), .A2(n885), .ZN(n704) );
  NAND2_X1 U774 ( .A1(G129), .A2(n886), .ZN(n703) );
  NAND2_X1 U775 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U777 ( .A1(n889), .A2(G141), .ZN(n707) );
  NAND2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n882) );
  NAND2_X1 U779 ( .A1(G1996), .A2(n882), .ZN(n717) );
  NAND2_X1 U780 ( .A1(G107), .A2(n885), .ZN(n710) );
  NAND2_X1 U781 ( .A1(G131), .A2(n889), .ZN(n709) );
  NAND2_X1 U782 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U783 ( .A1(G119), .A2(n886), .ZN(n711) );
  XNOR2_X1 U784 ( .A(KEYINPUT93), .B(n711), .ZN(n712) );
  NOR2_X1 U785 ( .A1(n713), .A2(n712), .ZN(n715) );
  NAND2_X1 U786 ( .A1(n890), .A2(G95), .ZN(n714) );
  NAND2_X1 U787 ( .A1(n715), .A2(n714), .ZN(n883) );
  NAND2_X1 U788 ( .A1(G1991), .A2(n883), .ZN(n716) );
  NAND2_X1 U789 ( .A1(n717), .A2(n716), .ZN(n951) );
  NAND2_X1 U790 ( .A1(n951), .A2(n761), .ZN(n729) );
  XNOR2_X1 U791 ( .A(KEYINPUT37), .B(G2067), .ZN(n759) );
  NAND2_X1 U792 ( .A1(G116), .A2(n885), .ZN(n719) );
  NAND2_X1 U793 ( .A1(G128), .A2(n886), .ZN(n718) );
  NAND2_X1 U794 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U795 ( .A(KEYINPUT35), .B(n720), .Z(n727) );
  NAND2_X1 U796 ( .A1(G140), .A2(n889), .ZN(n722) );
  NAND2_X1 U797 ( .A1(G104), .A2(n890), .ZN(n721) );
  NAND2_X1 U798 ( .A1(n722), .A2(n721), .ZN(n725) );
  XNOR2_X1 U799 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n723) );
  XNOR2_X1 U800 ( .A(n723), .B(KEYINPUT34), .ZN(n724) );
  XOR2_X1 U801 ( .A(n725), .B(n724), .Z(n726) );
  NOR2_X1 U802 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U803 ( .A(KEYINPUT36), .B(n728), .ZN(n906) );
  NOR2_X1 U804 ( .A1(n759), .A2(n906), .ZN(n957) );
  NAND2_X1 U805 ( .A1(n957), .A2(n761), .ZN(n748) );
  AND2_X1 U806 ( .A1(n729), .A2(n748), .ZN(n733) );
  AND2_X1 U807 ( .A1(n730), .A2(n733), .ZN(n731) );
  NAND2_X1 U808 ( .A1(n732), .A2(n731), .ZN(n767) );
  INV_X1 U809 ( .A(n733), .ZN(n747) );
  NAND2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n738) );
  NOR2_X1 U811 ( .A1(G2090), .A2(G303), .ZN(n736) );
  NAND2_X1 U812 ( .A1(G8), .A2(n736), .ZN(n737) );
  NAND2_X1 U813 ( .A1(n738), .A2(n737), .ZN(n739) );
  AND2_X1 U814 ( .A1(n739), .A2(n743), .ZN(n745) );
  NOR2_X1 U815 ( .A1(G1981), .A2(G305), .ZN(n740) );
  XOR2_X1 U816 ( .A(n740), .B(KEYINPUT24), .Z(n741) );
  XNOR2_X1 U817 ( .A(KEYINPUT96), .B(n741), .ZN(n742) );
  NOR2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U819 ( .A1(n513), .A2(n514), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n765) );
  INV_X1 U821 ( .A(n748), .ZN(n758) );
  NOR2_X1 U822 ( .A1(n882), .A2(G1996), .ZN(n749) );
  XNOR2_X1 U823 ( .A(n749), .B(KEYINPUT102), .ZN(n960) );
  NOR2_X1 U824 ( .A1(n883), .A2(G1991), .ZN(n750) );
  XNOR2_X1 U825 ( .A(n750), .B(KEYINPUT104), .ZN(n952) );
  NOR2_X1 U826 ( .A1(G1986), .A2(G290), .ZN(n751) );
  XOR2_X1 U827 ( .A(n751), .B(KEYINPUT103), .Z(n752) );
  NOR2_X1 U828 ( .A1(n952), .A2(n752), .ZN(n753) );
  NOR2_X1 U829 ( .A1(n753), .A2(n951), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n960), .A2(n754), .ZN(n755) );
  XNOR2_X1 U831 ( .A(KEYINPUT39), .B(n755), .ZN(n756) );
  NAND2_X1 U832 ( .A1(n756), .A2(n761), .ZN(n757) );
  OR2_X1 U833 ( .A1(n758), .A2(n757), .ZN(n763) );
  NAND2_X1 U834 ( .A1(n906), .A2(n759), .ZN(n760) );
  XNOR2_X1 U835 ( .A(n760), .B(KEYINPUT105), .ZN(n965) );
  NAND2_X1 U836 ( .A1(n965), .A2(n761), .ZN(n762) );
  NAND2_X1 U837 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U838 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U839 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U840 ( .A(n768), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U841 ( .A(G2443), .B(G2446), .Z(n770) );
  XNOR2_X1 U842 ( .A(G2427), .B(G2451), .ZN(n769) );
  XNOR2_X1 U843 ( .A(n770), .B(n769), .ZN(n776) );
  XOR2_X1 U844 ( .A(G2430), .B(G2454), .Z(n772) );
  XNOR2_X1 U845 ( .A(G1348), .B(G1341), .ZN(n771) );
  XNOR2_X1 U846 ( .A(n772), .B(n771), .ZN(n774) );
  XOR2_X1 U847 ( .A(G2435), .B(G2438), .Z(n773) );
  XNOR2_X1 U848 ( .A(n774), .B(n773), .ZN(n775) );
  XOR2_X1 U849 ( .A(n776), .B(n775), .Z(n777) );
  AND2_X1 U850 ( .A1(G14), .A2(n777), .ZN(G401) );
  AND2_X1 U851 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U852 ( .A(G132), .ZN(G219) );
  INV_X1 U853 ( .A(G82), .ZN(G220) );
  NAND2_X1 U854 ( .A1(G7), .A2(G661), .ZN(n778) );
  XNOR2_X1 U855 ( .A(n778), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U856 ( .A(G223), .ZN(n843) );
  NAND2_X1 U857 ( .A1(n843), .A2(G567), .ZN(n779) );
  XOR2_X1 U858 ( .A(KEYINPUT11), .B(n779), .Z(G234) );
  INV_X1 U859 ( .A(G860), .ZN(n784) );
  OR2_X1 U860 ( .A1(n921), .A2(n784), .ZN(G153) );
  NOR2_X1 U861 ( .A1(n929), .A2(G868), .ZN(n781) );
  INV_X1 U862 ( .A(G868), .ZN(n827) );
  NOR2_X1 U863 ( .A1(n827), .A2(G301), .ZN(n780) );
  NOR2_X1 U864 ( .A1(n781), .A2(n780), .ZN(G284) );
  NAND2_X1 U865 ( .A1(G868), .A2(G286), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G299), .A2(n827), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n784), .A2(G559), .ZN(n785) );
  INV_X1 U869 ( .A(n929), .ZN(n805) );
  NAND2_X1 U870 ( .A1(n785), .A2(n805), .ZN(n786) );
  XNOR2_X1 U871 ( .A(n786), .B(KEYINPUT16), .ZN(n788) );
  XOR2_X1 U872 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n787) );
  XNOR2_X1 U873 ( .A(n788), .B(n787), .ZN(G148) );
  NOR2_X1 U874 ( .A1(n929), .A2(n827), .ZN(n789) );
  XOR2_X1 U875 ( .A(KEYINPUT84), .B(n789), .Z(n790) );
  NOR2_X1 U876 ( .A1(G559), .A2(n790), .ZN(n793) );
  NOR2_X1 U877 ( .A1(G868), .A2(n921), .ZN(n791) );
  XOR2_X1 U878 ( .A(KEYINPUT83), .B(n791), .Z(n792) );
  NOR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(G282) );
  NAND2_X1 U880 ( .A1(n886), .A2(G123), .ZN(n794) );
  XNOR2_X1 U881 ( .A(n794), .B(KEYINPUT18), .ZN(n796) );
  NAND2_X1 U882 ( .A1(G135), .A2(n889), .ZN(n795) );
  NAND2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(KEYINPUT85), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G99), .A2(n890), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U887 ( .A1(n885), .A2(G111), .ZN(n800) );
  XOR2_X1 U888 ( .A(KEYINPUT86), .B(n800), .Z(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n953) );
  XNOR2_X1 U890 ( .A(n953), .B(G2096), .ZN(n804) );
  INV_X1 U891 ( .A(G2100), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(G156) );
  NAND2_X1 U893 ( .A1(G559), .A2(n805), .ZN(n825) );
  XNOR2_X1 U894 ( .A(n921), .B(n825), .ZN(n806) );
  NOR2_X1 U895 ( .A1(n806), .A2(G860), .ZN(n817) );
  NAND2_X1 U896 ( .A1(G67), .A2(n807), .ZN(n810) );
  NAND2_X1 U897 ( .A1(G93), .A2(n808), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n810), .A2(n809), .ZN(n816) );
  NAND2_X1 U899 ( .A1(n811), .A2(G80), .ZN(n814) );
  NAND2_X1 U900 ( .A1(G55), .A2(n812), .ZN(n813) );
  NAND2_X1 U901 ( .A1(n814), .A2(n813), .ZN(n815) );
  OR2_X1 U902 ( .A1(n816), .A2(n815), .ZN(n828) );
  XOR2_X1 U903 ( .A(n817), .B(n828), .Z(G145) );
  XNOR2_X1 U904 ( .A(KEYINPUT19), .B(n828), .ZN(n818) );
  XNOR2_X1 U905 ( .A(G290), .B(n818), .ZN(n819) );
  XNOR2_X1 U906 ( .A(n819), .B(G305), .ZN(n823) );
  XNOR2_X1 U907 ( .A(n820), .B(n921), .ZN(n821) );
  XNOR2_X1 U908 ( .A(n821), .B(G288), .ZN(n822) );
  XNOR2_X1 U909 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U910 ( .A(G166), .B(n824), .ZN(n910) );
  XOR2_X1 U911 ( .A(n910), .B(n825), .Z(n826) );
  NOR2_X1 U912 ( .A1(n827), .A2(n826), .ZN(n830) );
  NOR2_X1 U913 ( .A1(G868), .A2(n828), .ZN(n829) );
  NOR2_X1 U914 ( .A1(n830), .A2(n829), .ZN(G295) );
  NAND2_X1 U915 ( .A1(G2084), .A2(G2078), .ZN(n831) );
  XOR2_X1 U916 ( .A(KEYINPUT20), .B(n831), .Z(n832) );
  NAND2_X1 U917 ( .A1(G2090), .A2(n832), .ZN(n833) );
  XNOR2_X1 U918 ( .A(KEYINPUT21), .B(n833), .ZN(n834) );
  NAND2_X1 U919 ( .A1(n834), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U920 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  XNOR2_X1 U921 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U922 ( .A1(G108), .A2(G120), .ZN(n835) );
  NOR2_X1 U923 ( .A1(G237), .A2(n835), .ZN(n836) );
  NAND2_X1 U924 ( .A1(G69), .A2(n836), .ZN(n919) );
  NAND2_X1 U925 ( .A1(n919), .A2(G567), .ZN(n841) );
  NOR2_X1 U926 ( .A1(G220), .A2(G219), .ZN(n837) );
  XOR2_X1 U927 ( .A(KEYINPUT22), .B(n837), .Z(n838) );
  NOR2_X1 U928 ( .A1(G218), .A2(n838), .ZN(n839) );
  NAND2_X1 U929 ( .A1(G96), .A2(n839), .ZN(n920) );
  NAND2_X1 U930 ( .A1(n920), .A2(G2106), .ZN(n840) );
  NAND2_X1 U931 ( .A1(n841), .A2(n840), .ZN(n847) );
  NAND2_X1 U932 ( .A1(G483), .A2(G661), .ZN(n842) );
  NOR2_X1 U933 ( .A1(n847), .A2(n842), .ZN(n846) );
  NAND2_X1 U934 ( .A1(n846), .A2(G36), .ZN(G176) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U937 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U939 ( .A1(n846), .A2(n845), .ZN(G188) );
  XOR2_X1 U940 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  INV_X1 U941 ( .A(n847), .ZN(G319) );
  XOR2_X1 U942 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n849) );
  XNOR2_X1 U943 ( .A(G2678), .B(KEYINPUT107), .ZN(n848) );
  XNOR2_X1 U944 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U945 ( .A(KEYINPUT43), .B(G2072), .Z(n851) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2090), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U948 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U949 ( .A(G2096), .B(G2100), .ZN(n854) );
  XNOR2_X1 U950 ( .A(n855), .B(n854), .ZN(n857) );
  XOR2_X1 U951 ( .A(G2084), .B(G2078), .Z(n856) );
  XNOR2_X1 U952 ( .A(n857), .B(n856), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1986), .B(G1976), .Z(n859) );
  XNOR2_X1 U954 ( .A(G1971), .B(G1961), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U956 ( .A(n860), .B(KEYINPUT41), .Z(n862) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n861) );
  XNOR2_X1 U958 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U959 ( .A(G2474), .B(G1981), .Z(n864) );
  XNOR2_X1 U960 ( .A(G1966), .B(G1956), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n866), .B(n865), .ZN(G229) );
  NAND2_X1 U963 ( .A1(G112), .A2(n885), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G100), .A2(n890), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U966 ( .A1(n886), .A2(G124), .ZN(n869) );
  XNOR2_X1 U967 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G136), .A2(n889), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U970 ( .A(KEYINPUT109), .B(n872), .Z(n873) );
  NOR2_X1 U971 ( .A1(n874), .A2(n873), .ZN(G162) );
  XNOR2_X1 U972 ( .A(G162), .B(n953), .ZN(n905) );
  NAND2_X1 U973 ( .A1(G139), .A2(n889), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G103), .A2(n890), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n881) );
  NAND2_X1 U976 ( .A1(G115), .A2(n885), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G127), .A2(n886), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n946) );
  XNOR2_X1 U981 ( .A(n946), .B(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n901) );
  XOR2_X1 U983 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n899) );
  NAND2_X1 U984 ( .A1(G118), .A2(n885), .ZN(n888) );
  NAND2_X1 U985 ( .A1(G130), .A2(n886), .ZN(n887) );
  NAND2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n896) );
  NAND2_X1 U987 ( .A1(G142), .A2(n889), .ZN(n892) );
  NAND2_X1 U988 ( .A1(G106), .A2(n890), .ZN(n891) );
  NAND2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U990 ( .A(KEYINPUT110), .B(n893), .Z(n894) );
  XNOR2_X1 U991 ( .A(KEYINPUT45), .B(n894), .ZN(n895) );
  NOR2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n897), .B(KEYINPUT48), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U995 ( .A(n901), .B(n900), .Z(n903) );
  XNOR2_X1 U996 ( .A(G164), .B(G160), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n907) );
  XOR2_X1 U999 ( .A(n907), .B(n906), .Z(n908) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n908), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(n929), .B(G286), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n909), .B(G301), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n913) );
  XOR2_X1 U1006 ( .A(KEYINPUT49), .B(n913), .Z(n914) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n914), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n915), .ZN(n916) );
  XNOR2_X1 U1009 ( .A(KEYINPUT112), .B(n916), .ZN(n918) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(G225) );
  XNOR2_X1 U1012 ( .A(KEYINPUT113), .B(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(G96), .ZN(G221) );
  INV_X1 U1016 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(G325) );
  INV_X1 U1018 ( .A(G325), .ZN(G261) );
  INV_X1 U1019 ( .A(G301), .ZN(G171) );
  XOR2_X1 U1020 ( .A(n921), .B(G1341), .Z(n938) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n925) );
  AND2_X1 U1022 ( .A1(G303), .A2(G1971), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(n926), .B(KEYINPUT119), .ZN(n935) );
  XNOR2_X1 U1025 ( .A(G1961), .B(G301), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(G299), .B(G1956), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n929), .B(G1348), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(KEYINPUT120), .B(n936), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n943) );
  XNOR2_X1 U1034 ( .A(G1966), .B(G168), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT57), .B(n941), .Z(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n945) );
  XOR2_X1 U1038 ( .A(KEYINPUT56), .B(G16), .Z(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n975) );
  XOR2_X1 U1040 ( .A(G2072), .B(n946), .Z(n948) );
  XOR2_X1 U1041 ( .A(G164), .B(G2078), .Z(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1043 ( .A(KEYINPUT50), .B(n949), .Z(n968) );
  XOR2_X1 U1044 ( .A(G160), .B(G2084), .Z(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n955) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(KEYINPUT114), .B(n958), .ZN(n963) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n959) );
  NOR2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1052 ( .A(KEYINPUT51), .B(n961), .Z(n962) );
  NAND2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1054 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(KEYINPUT115), .B(n966), .ZN(n967) );
  NOR2_X1 U1056 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(n969), .B(KEYINPUT52), .ZN(n971) );
  INV_X1 U1058 ( .A(KEYINPUT55), .ZN(n970) );
  NAND2_X1 U1059 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1060 ( .A1(G29), .A2(n972), .ZN(n973) );
  XOR2_X1 U1061 ( .A(KEYINPUT116), .B(n973), .Z(n974) );
  NOR2_X1 U1062 ( .A1(n975), .A2(n974), .ZN(n1029) );
  XOR2_X1 U1063 ( .A(G1961), .B(G5), .Z(n985) );
  XOR2_X1 U1064 ( .A(G1986), .B(G24), .Z(n980) );
  XNOR2_X1 U1065 ( .A(G1971), .B(G22), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(G1976), .B(G23), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(n978), .B(KEYINPUT124), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n983) );
  XNOR2_X1 U1070 ( .A(KEYINPUT58), .B(KEYINPUT126), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(n981), .B(KEYINPUT125), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(n983), .B(n982), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(n985), .A2(n984), .ZN(n1000) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G21), .ZN(n997) );
  XNOR2_X1 U1075 ( .A(KEYINPUT59), .B(KEYINPUT121), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(n986), .B(G4), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(G1348), .B(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(G1981), .B(G6), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G1956), .B(G20), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(G1341), .B(G19), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(KEYINPUT122), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(KEYINPUT60), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(n998), .B(KEYINPUT123), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(KEYINPUT61), .B(n1001), .Z(n1002) );
  NOR2_X1 U1090 ( .A1(G16), .A2(n1002), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(KEYINPUT127), .B(n1003), .Z(n1027) );
  XNOR2_X1 U1092 ( .A(G2067), .B(G26), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G1996), .B(G32), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1011) );
  XOR2_X1 U1095 ( .A(G2072), .B(G33), .Z(n1006) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(G28), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(G25), .B(G1991), .Z(n1007) );
  XNOR2_X1 U1098 ( .A(KEYINPUT117), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G27), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1103 ( .A(KEYINPUT53), .B(n1015), .Z(n1018) );
  XOR2_X1 U1104 ( .A(KEYINPUT54), .B(G34), .Z(n1016) );
  XNOR2_X1 U1105 ( .A(G2084), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G35), .B(G2090), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(n1021), .B(KEYINPUT55), .ZN(n1023) );
  INV_X1 U1110 ( .A(G29), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(G11), .A2(n1024), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(KEYINPUT118), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

