//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n531, new_n532, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n583, new_n586, new_n587, new_n589, new_n590, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  OR2_X1    g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  AOI21_X1  g034(.A(G2105), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n460), .A2(G137), .B1(G101), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G160));
  OAI21_X1  g042(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G112), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  XOR2_X1   g048(.A(new_n473), .B(KEYINPUT67), .Z(new_n474));
  AOI211_X1 g049(.A(new_n470), .B(new_n474), .C1(G136), .C2(new_n460), .ZN(G162));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  OAI211_X1 g052(.A(G126), .B(G2105), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G114), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT68), .ZN(new_n483));
  OAI211_X1 g058(.A(G138), .B(new_n461), .C1(new_n476), .C2(new_n477), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n464), .A2(new_n486), .A3(G138), .A4(new_n461), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n478), .A2(new_n481), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n483), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  OR2_X1    g067(.A1(KEYINPUT5), .A2(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT5), .A2(G543), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n495), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n496));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT6), .B(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G88), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OR2_X1    g079(.A1(new_n498), .A2(new_n504), .ZN(G303));
  INV_X1    g080(.A(G303), .ZN(G166));
  INV_X1    g081(.A(new_n502), .ZN(new_n507));
  AND2_X1   g082(.A1(G63), .A2(G651), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n507), .A2(G51), .B1(new_n495), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT69), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT7), .ZN(new_n512));
  INV_X1    g087(.A(G89), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(new_n500), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n509), .B1(new_n514), .B2(KEYINPUT70), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(KEYINPUT70), .B2(new_n514), .ZN(G168));
  AOI22_X1  g091(.A1(new_n495), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(new_n497), .ZN(new_n518));
  INV_X1    g093(.A(G90), .ZN(new_n519));
  INV_X1    g094(.A(G52), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n500), .A2(new_n519), .B1(new_n502), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(G171));
  AOI22_X1  g097(.A1(new_n495), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n497), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT71), .B(G81), .Z(new_n525));
  INV_X1    g100(.A(G43), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n500), .A2(new_n525), .B1(new_n502), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G860), .ZN(G153));
  NAND4_X1  g104(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g105(.A1(G1), .A2(G3), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT8), .ZN(new_n532));
  NAND4_X1  g107(.A1(G319), .A2(G483), .A3(G661), .A4(new_n532), .ZN(G188));
  NAND2_X1  g108(.A1(G78), .A2(G543), .ZN(new_n534));
  AND2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G65), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n495), .A2(new_n499), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G91), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n499), .A2(G53), .A3(G543), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n543), .A2(KEYINPUT9), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(KEYINPUT9), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n540), .B(new_n542), .C1(new_n544), .C2(new_n545), .ZN(G299));
  INV_X1    g121(.A(G171), .ZN(G301));
  OR2_X1    g122(.A1(new_n514), .A2(KEYINPUT70), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n514), .A2(KEYINPUT70), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(new_n549), .A3(new_n509), .ZN(G286));
  NAND2_X1  g125(.A1(new_n507), .A2(G49), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n541), .A2(G87), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n495), .B2(G74), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(G288));
  NAND2_X1  g129(.A1(new_n495), .A2(G61), .ZN(new_n555));
  NAND2_X1  g130(.A1(G73), .A2(G543), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n497), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n495), .A2(new_n499), .A3(G86), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n499), .A2(G48), .A3(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(G305));
  AOI22_X1  g137(.A1(new_n495), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n497), .ZN(new_n564));
  INV_X1    g139(.A(G85), .ZN(new_n565));
  INV_X1    g140(.A(G47), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n500), .A2(new_n565), .B1(new_n502), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G290));
  NAND2_X1  g144(.A1(G79), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G66), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n537), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(G54), .A2(new_n507), .B1(new_n572), .B2(G651), .ZN(new_n573));
  INV_X1    g148(.A(G92), .ZN(new_n574));
  XNOR2_X1  g149(.A(KEYINPUT72), .B(KEYINPUT10), .ZN(new_n575));
  OR3_X1    g150(.A1(new_n500), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n500), .B2(new_n574), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G868), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n579), .B2(G171), .ZN(G284));
  OAI21_X1  g156(.A(new_n580), .B1(new_n579), .B2(G171), .ZN(G321));
  NAND2_X1  g157(.A1(G299), .A2(new_n579), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(G168), .B2(new_n579), .ZN(G297));
  OAI21_X1  g159(.A(new_n583), .B1(G168), .B2(new_n579), .ZN(G280));
  INV_X1    g160(.A(new_n578), .ZN(new_n586));
  INV_X1    g161(.A(G559), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(G860), .ZN(G148));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G868), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(G868), .B2(new_n528), .ZN(G323));
  XNOR2_X1  g166(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g167(.A1(new_n464), .A2(new_n462), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT12), .ZN(new_n594));
  XNOR2_X1  g169(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G2100), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT74), .Z(new_n598));
  NAND2_X1  g173(.A1(new_n460), .A2(G135), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n461), .A2(G111), .ZN(new_n600));
  OAI21_X1  g175(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n601));
  INV_X1    g176(.A(G123), .ZN(new_n602));
  OAI221_X1 g177(.A(new_n599), .B1(new_n600), .B2(new_n601), .C1(new_n602), .C2(new_n471), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT75), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(G2096), .Z(new_n605));
  OAI211_X1 g180(.A(new_n598), .B(new_n605), .C1(G2100), .C2(new_n596), .ZN(G156));
  INV_X1    g181(.A(KEYINPUT14), .ZN(new_n607));
  XNOR2_X1  g182(.A(G2427), .B(G2438), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2430), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT15), .B(G2435), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n610), .B2(new_n609), .ZN(new_n612));
  XNOR2_X1  g187(.A(G2451), .B(G2454), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT16), .ZN(new_n614));
  XOR2_X1   g189(.A(G1341), .B(G1348), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n612), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(G2443), .B(G2446), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n617), .A2(new_n619), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(G14), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT76), .Z(G401));
  XOR2_X1   g198(.A(KEYINPUT77), .B(KEYINPUT18), .Z(new_n624));
  XOR2_X1   g199(.A(G2084), .B(G2090), .Z(new_n625));
  XNOR2_X1  g200(.A(G2067), .B(G2678), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT17), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n625), .A2(new_n626), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT78), .Z(new_n631));
  XOR2_X1   g206(.A(G2072), .B(G2078), .Z(new_n632));
  INV_X1    g207(.A(new_n624), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n632), .B1(new_n627), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2096), .B(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(G227));
  XOR2_X1   g212(.A(G1991), .B(G1996), .Z(new_n638));
  XNOR2_X1  g213(.A(G1961), .B(G1966), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT79), .ZN(new_n640));
  XOR2_X1   g215(.A(G1956), .B(G2474), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1971), .B(G1976), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT19), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n641), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n644), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n647), .A2(KEYINPUT20), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(KEYINPUT20), .ZN(new_n649));
  OAI221_X1 g224(.A(new_n646), .B1(new_n644), .B2(new_n642), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n652), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n638), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n650), .A2(new_n652), .ZN(new_n656));
  INV_X1    g231(.A(new_n638), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n650), .A2(new_n652), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1981), .B(G1986), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n655), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n660), .B1(new_n655), .B2(new_n659), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(G229));
  INV_X1    g238(.A(G16), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G22), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(G166), .B2(new_n664), .ZN(new_n666));
  INV_X1    g241(.A(G1971), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(G6), .A2(G16), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n561), .B2(G16), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT32), .B(G1981), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n664), .A2(G23), .ZN(new_n673));
  INV_X1    g248(.A(G288), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n673), .B1(new_n674), .B2(new_n664), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT33), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n668), .A2(new_n672), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT34), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n460), .A2(G131), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT80), .Z(new_n681));
  OAI21_X1  g256(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n682));
  INV_X1    g257(.A(G107), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(G2105), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n472), .B2(G119), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  MUX2_X1   g261(.A(G25), .B(new_n686), .S(G29), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT35), .B(G1991), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n664), .A2(G24), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT81), .Z(new_n692));
  NOR2_X1   g267(.A1(G290), .A2(KEYINPUT82), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n694));
  OAI21_X1  g269(.A(G16), .B1(new_n568), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n692), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n690), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n679), .B(new_n700), .C1(new_n699), .C2(new_n698), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT84), .B(KEYINPUT36), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n664), .A2(G4), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n586), .B2(new_n664), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT85), .B(G1348), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n664), .A2(G19), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n528), .B2(new_n664), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G1341), .Z(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G26), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT86), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  OR2_X1    g289(.A1(G104), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n716));
  OAI211_X1 g291(.A(G140), .B(new_n461), .C1(new_n476), .C2(new_n477), .ZN(new_n717));
  OAI211_X1 g292(.A(G128), .B(G2105), .C1(new_n476), .C2(new_n477), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n711), .B2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(G2067), .Z(new_n722));
  NAND3_X1  g297(.A1(new_n707), .A2(new_n710), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT87), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n711), .A2(G35), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G162), .B2(new_n711), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n727));
  INV_X1    g302(.A(G2090), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n726), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G29), .A2(G33), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT88), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT25), .Z(new_n734));
  INV_X1    g309(.A(G139), .ZN(new_n735));
  INV_X1    g310(.A(new_n460), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n464), .A2(G127), .ZN(new_n738));
  NAND2_X1  g313(.A1(G115), .A2(G2104), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n461), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n732), .B1(new_n741), .B2(new_n711), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G2072), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n664), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n664), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1961), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT31), .B(G11), .ZN(new_n747));
  INV_X1    g322(.A(G28), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n748), .B2(KEYINPUT30), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(KEYINPUT92), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n751));
  OR3_X1    g326(.A1(new_n751), .A2(new_n748), .A3(KEYINPUT30), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n749), .A2(KEYINPUT92), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n751), .B1(new_n748), .B2(KEYINPUT30), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT24), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n711), .B1(new_n756), .B2(G34), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n756), .A2(G34), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n466), .A2(new_n711), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n747), .B1(new_n750), .B2(new_n755), .C1(new_n763), .C2(G2084), .ZN(new_n764));
  OR3_X1    g339(.A1(new_n743), .A2(new_n746), .A3(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n462), .A2(G105), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n460), .A2(G141), .ZN(new_n771));
  INV_X1    g346(.A(G129), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n471), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(new_n711), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n711), .B2(G32), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n776), .A2(new_n777), .B1(G2084), .B2(new_n763), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n778), .B1(new_n711), .B2(new_n604), .C1(new_n776), .C2(new_n777), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n711), .A2(G27), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G164), .B2(new_n711), .ZN(new_n781));
  INV_X1    g356(.A(G2078), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n664), .A2(G20), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT23), .Z(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G299), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1956), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n730), .A2(new_n765), .A3(new_n779), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n664), .A2(G21), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G168), .B2(new_n664), .ZN(new_n791));
  INV_X1    g366(.A(G1966), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AND4_X1   g368(.A1(new_n703), .A2(new_n724), .A3(new_n789), .A4(new_n793), .ZN(G311));
  NAND4_X1  g369(.A1(new_n703), .A2(new_n724), .A3(new_n789), .A4(new_n793), .ZN(G150));
  AOI22_X1  g370(.A1(new_n495), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(new_n497), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT94), .B(G55), .Z(new_n798));
  NAND3_X1  g373(.A1(new_n798), .A2(G543), .A3(new_n499), .ZN(new_n799));
  INV_X1    g374(.A(G93), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n500), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT95), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n541), .A2(G93), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n799), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n797), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G860), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT37), .Z(new_n808));
  INV_X1    g383(.A(G860), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n578), .A2(new_n587), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT96), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT38), .ZN(new_n812));
  INV_X1    g387(.A(new_n528), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n804), .A2(new_n803), .A3(new_n799), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n817), .A2(new_n528), .A3(new_n797), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n812), .B(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n809), .B1(new_n821), .B2(KEYINPUT39), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n812), .B(new_n819), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n824));
  OR3_X1    g399(.A1(new_n823), .A2(KEYINPUT97), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT97), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI211_X1 g404(.A(KEYINPUT98), .B(new_n822), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n808), .B1(new_n829), .B2(new_n830), .ZN(G145));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n686), .B(new_n594), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n472), .A2(G130), .B1(G142), .B2(new_n460), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n836));
  INV_X1    g411(.A(G118), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n835), .A2(new_n836), .B1(new_n837), .B2(G2105), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n836), .B2(new_n835), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n833), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n482), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n485), .A2(new_n487), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n485), .B2(new_n487), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n720), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n842), .B(new_n719), .C1(new_n844), .C2(new_n845), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n847), .A2(new_n774), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n774), .B1(new_n847), .B2(new_n848), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT101), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n774), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n488), .A2(KEYINPUT100), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n485), .A2(new_n487), .A3(new_n843), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n719), .B1(new_n855), .B2(new_n842), .ZN(new_n856));
  INV_X1    g431(.A(new_n848), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n847), .A2(new_n774), .A3(new_n848), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  INV_X1    g437(.A(new_n741), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n851), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n851), .A2(new_n863), .A3(new_n861), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n858), .A2(new_n741), .A3(new_n860), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT102), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n841), .B(new_n864), .C1(new_n865), .C2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT106), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n841), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n858), .A2(new_n860), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n741), .B1(new_n872), .B2(KEYINPUT101), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n867), .B1(new_n873), .B2(new_n861), .ZN(new_n874));
  INV_X1    g449(.A(new_n864), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n466), .B(KEYINPUT99), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n604), .B(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G162), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n851), .A2(new_n863), .A3(new_n861), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(KEYINPUT102), .A3(new_n866), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n881), .A2(KEYINPUT106), .A3(new_n841), .A4(new_n864), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n870), .A2(new_n876), .A3(new_n879), .A4(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n876), .A2(new_n887), .A3(new_n868), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n881), .A2(KEYINPUT104), .A3(new_n841), .A4(new_n864), .ZN(new_n889));
  INV_X1    g464(.A(new_n879), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n886), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n876), .A2(new_n887), .A3(new_n868), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n893), .A2(KEYINPUT105), .A3(new_n890), .A4(new_n889), .ZN(new_n894));
  AOI211_X1 g469(.A(new_n832), .B(new_n885), .C1(new_n892), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n894), .ZN(new_n896));
  INV_X1    g471(.A(new_n885), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT40), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n895), .A2(new_n898), .ZN(G395));
  XNOR2_X1  g474(.A(new_n819), .B(new_n589), .ZN(new_n900));
  INV_X1    g475(.A(G299), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n576), .A2(new_n577), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n573), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n578), .A2(G299), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT41), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(new_n907), .A3(new_n904), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n900), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n905), .B2(new_n900), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n674), .B(G303), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n568), .B(new_n561), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n913), .B2(new_n914), .ZN(new_n919));
  OAI21_X1  g494(.A(G868), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n806), .A2(new_n579), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(G295));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n921), .ZN(G331));
  INV_X1    g498(.A(new_n818), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n528), .B1(new_n817), .B2(new_n797), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n924), .A2(G171), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(G301), .B1(new_n814), .B2(new_n818), .ZN(new_n927));
  OAI21_X1  g502(.A(G286), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(G171), .B1(new_n924), .B2(new_n925), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n814), .A2(G301), .A3(new_n818), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(G168), .A3(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n928), .A2(new_n909), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n905), .B1(new_n928), .B2(new_n931), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n932), .A2(new_n933), .A3(KEYINPUT107), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n935));
  INV_X1    g510(.A(new_n905), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n926), .A2(new_n927), .A3(G286), .ZN(new_n937));
  AOI21_X1  g512(.A(G168), .B1(new_n929), .B2(new_n930), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n928), .A2(new_n909), .A3(new_n931), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n917), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n934), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(new_n942), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n884), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT43), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  INV_X1    g522(.A(new_n945), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n908), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n903), .A2(KEYINPUT108), .A3(new_n907), .A4(new_n904), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n906), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n928), .A2(new_n952), .A3(new_n953), .A4(new_n931), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n954), .A2(new_n917), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n928), .A2(new_n952), .A3(new_n931), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n939), .A2(KEYINPUT109), .A3(new_n956), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n955), .A2(new_n957), .A3(KEYINPUT110), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT110), .B1(new_n955), .B2(new_n957), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n947), .B(new_n948), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n946), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n947), .B1(new_n943), .B2(new_n945), .ZN(new_n962));
  OAI211_X1 g537(.A(KEYINPUT43), .B(new_n948), .C1(new_n958), .C2(new_n959), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  MUX2_X1   g539(.A(new_n961), .B(new_n964), .S(KEYINPUT44), .Z(G397));
  OAI211_X1 g540(.A(new_n463), .B(G40), .C1(new_n461), .C2(new_n465), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n491), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n846), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n971));
  AOI21_X1  g546(.A(G1971), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n966), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n975));
  XOR2_X1   g550(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n846), .B2(new_n967), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n973), .B1(G2090), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G8), .ZN(new_n980));
  NAND2_X1  g555(.A1(G303), .A2(G8), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(G1981), .B1(new_n557), .B2(new_n560), .ZN(new_n986));
  INV_X1    g561(.A(G61), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n493), .B2(new_n494), .ZN(new_n988));
  INV_X1    g563(.A(new_n556), .ZN(new_n989));
  OAI21_X1  g564(.A(G651), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1981), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n558), .A4(new_n559), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n986), .A2(KEYINPUT114), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n995), .B(G1981), .C1(new_n557), .C2(new_n560), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n994), .B1(new_n993), .B2(new_n996), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n846), .A2(new_n974), .A3(new_n967), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1001), .A2(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n674), .A2(G1976), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(G8), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1000), .A2(new_n1002), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n966), .B1(new_n968), .B2(KEYINPUT50), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n846), .A2(new_n967), .A3(new_n976), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1009), .A2(new_n728), .A3(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n983), .B(G8), .C1(new_n1011), .C2(new_n972), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1004), .A2(KEYINPUT113), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1001), .A2(new_n1014), .A3(G8), .A4(new_n1003), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(KEYINPUT52), .A3(new_n1015), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1008), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2084), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1009), .A2(new_n1018), .A3(new_n1010), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n974), .B1(new_n968), .B2(new_n969), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT45), .B1(new_n846), .B2(new_n967), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n792), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1009), .A2(KEYINPUT115), .A3(new_n1010), .A4(new_n1018), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G286), .A2(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1026), .A2(KEYINPUT116), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT116), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n985), .B(new_n1017), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1030), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1026), .A2(KEYINPUT116), .A3(new_n1028), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(G8), .B1(new_n1011), .B2(new_n972), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n984), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT63), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1008), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1031), .A2(new_n1033), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g617(.A(G1976), .B(G288), .C1(new_n1000), .C2(new_n1002), .ZN(new_n1043));
  INV_X1    g618(.A(new_n992), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1002), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1012), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(new_n1016), .A3(new_n1008), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT118), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n970), .A2(new_n782), .A3(new_n971), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1052));
  INV_X1    g627(.A(G1961), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1050), .A2(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(KEYINPUT53), .A3(new_n782), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(G301), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT126), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n465), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n465), .A2(new_n1059), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(G2105), .A3(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n463), .A2(G40), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT53), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1064), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1023), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n971), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1054), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT126), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1054), .A2(new_n1075), .A3(G301), .A4(new_n1056), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1058), .A2(new_n1074), .A3(KEYINPUT54), .A4(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n983), .B1(new_n979), .B2(G8), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(new_n1040), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1054), .A2(new_n1072), .A3(G301), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1081), .A2(KEYINPUT125), .B1(new_n1082), .B2(G171), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1054), .A2(new_n1072), .A3(new_n1084), .A4(G301), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT54), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1956), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n975), .B2(new_n977), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1090), .A2(KEYINPUT57), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(KEYINPUT57), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n901), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(G299), .A2(new_n1090), .A3(KEYINPUT57), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n970), .A2(new_n971), .A3(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1089), .A2(new_n1093), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1001), .A2(G2067), .ZN(new_n1098));
  INV_X1    g673(.A(new_n706), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1097), .B(new_n586), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1089), .A2(new_n1096), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1097), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT121), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1104), .A2(new_n1109), .A3(KEYINPUT61), .A4(new_n1097), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1100), .A2(new_n1098), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n578), .B1(new_n1112), .B2(KEYINPUT60), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n1114));
  NOR4_X1   g689(.A1(new_n1100), .A2(new_n1098), .A3(new_n1114), .A4(new_n586), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n1113), .A2(new_n1115), .B1(KEYINPUT60), .B2(new_n1112), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1117));
  INV_X1    g692(.A(G1996), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n970), .A2(new_n1118), .A3(new_n971), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT58), .B(G1341), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1001), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n813), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1116), .A2(new_n1117), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1105), .B1(new_n1111), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(G8), .B1(new_n1026), .B2(G286), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1127), .A2(KEYINPUT51), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1026), .A2(G286), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT51), .B1(new_n1129), .B2(new_n1127), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1087), .A2(new_n1126), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(KEYINPUT62), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1128), .A2(new_n1130), .A3(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1079), .A2(G171), .A3(new_n1082), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1048), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1032), .B1(new_n1036), .B2(new_n1079), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1017), .A2(KEYINPUT63), .A3(new_n1038), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1138), .B(new_n1139), .C1(new_n1140), .C2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1049), .A2(new_n1132), .A3(new_n1137), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1023), .A2(new_n974), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1146), .A2(new_n1118), .A3(new_n774), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT111), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1146), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n719), .B(G2067), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n852), .A2(G1996), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n688), .B1(new_n681), .B2(new_n685), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n686), .A2(new_n689), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1149), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n568), .A2(new_n697), .ZN(new_n1158));
  NAND2_X1  g733(.A1(G290), .A2(G1986), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1146), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1145), .A2(new_n1161), .ZN(new_n1162));
  OR3_X1    g737(.A1(new_n1146), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT46), .B1(new_n1146), .B2(G1996), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n852), .A2(new_n1150), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1163), .A2(new_n1164), .B1(new_n1149), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT47), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n719), .A2(G2067), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1146), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1157), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1146), .A2(new_n1158), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1172), .B(KEYINPUT48), .Z(new_n1173));
  AOI211_X1 g748(.A(new_n1167), .B(new_n1170), .C1(new_n1171), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1162), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g750(.A1(new_n896), .A2(new_n897), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n622), .A2(G319), .ZN(new_n1178));
  NOR2_X1   g752(.A1(G227), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1179), .B1(new_n661), .B2(new_n662), .ZN(new_n1180));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n1181));
  XNOR2_X1  g755(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  AND3_X1   g756(.A1(new_n1177), .A2(new_n961), .A3(new_n1182), .ZN(G308));
  NAND3_X1  g757(.A1(new_n1177), .A2(new_n961), .A3(new_n1182), .ZN(G225));
endmodule


