//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  XOR2_X1   g000(.A(KEYINPUT74), .B(G217), .Z(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT78), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n191), .A2(new_n193), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G146), .ZN(new_n200));
  XNOR2_X1  g014(.A(G125), .B(G140), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(KEYINPUT78), .A3(new_n202), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n197), .A2(G146), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT75), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT75), .A3(G119), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT24), .B(G110), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n206), .B2(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n216));
  INV_X1    g030(.A(G110), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n208), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n213), .A2(KEYINPUT77), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT77), .B1(new_n213), .B2(new_n218), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n204), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n215), .A2(new_n216), .A3(new_n208), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G110), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT76), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n225), .A3(G110), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n211), .A2(new_n212), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n196), .A2(new_n202), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n194), .A2(new_n195), .A3(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G137), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(G221), .A3(G234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n233), .B(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n221), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(new_n221), .B2(new_n232), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT25), .B1(new_n239), .B2(new_n188), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n221), .A2(new_n232), .ZN(new_n241));
  INV_X1    g055(.A(new_n236), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n221), .A2(new_n232), .A3(new_n236), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n243), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n189), .B1(new_n240), .B2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n189), .A2(G902), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n239), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n189), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n243), .A2(new_n188), .A3(new_n244), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT25), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n252), .B1(new_n255), .B2(new_n245), .ZN(new_n256));
  INV_X1    g070(.A(new_n249), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT79), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(G119), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n206), .A2(KEYINPUT70), .A3(G116), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(G119), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n267));
  INV_X1    g081(.A(G113), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n269), .A2(new_n270), .B1(KEYINPUT2), .B2(G113), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(KEYINPUT2), .A2(G113), .ZN(new_n273));
  INV_X1    g087(.A(new_n270), .ZN(new_n274));
  NOR3_X1   g088(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n280));
  INV_X1    g094(.A(G143), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n202), .A2(G143), .ZN(new_n283));
  OAI22_X1  g097(.A1(new_n280), .A2(new_n282), .B1(new_n283), .B2(G128), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n286));
  XNOR2_X1  g100(.A(G143), .B(G146), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n280), .ZN(new_n288));
  AND4_X1   g102(.A1(new_n286), .A2(new_n280), .A3(new_n282), .A4(new_n283), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT11), .ZN(new_n291));
  INV_X1    g105(.A(G134), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(G137), .ZN(new_n293));
  INV_X1    g107(.A(G137), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT11), .A3(G134), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(G137), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT66), .B(G131), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(G134), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n296), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n297), .A2(new_n298), .B1(G131), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G131), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n298), .A2(new_n293), .A3(new_n295), .A4(new_n296), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g119(.A1(KEYINPUT0), .A2(G128), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n282), .A2(new_n283), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT0), .B(G128), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n287), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n290), .A2(new_n301), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT30), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n287), .A2(new_n286), .A3(new_n280), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n284), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n300), .A2(G131), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n304), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT68), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT68), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n290), .A2(new_n320), .A3(new_n301), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n307), .B(KEYINPUT65), .C1(new_n287), .C2(new_n308), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n306), .ZN(new_n324));
  OR2_X1    g138(.A1(KEYINPUT0), .A2(G128), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n202), .A2(G143), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n281), .A2(G146), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT65), .B1(new_n328), .B2(new_n307), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n319), .A2(new_n321), .B1(new_n330), .B2(new_n305), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n279), .B(new_n312), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT31), .ZN(new_n335));
  INV_X1    g149(.A(new_n279), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n311), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT26), .B(G101), .ZN(new_n338));
  NOR2_X1   g152(.A1(G237), .A2(G953), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G210), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n338), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n334), .A2(new_n335), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n335), .B1(new_n334), .B2(new_n344), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n311), .A2(KEYINPUT28), .A3(new_n336), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT28), .B1(new_n311), .B2(new_n336), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n319), .A2(new_n321), .ZN(new_n350));
  INV_X1    g164(.A(new_n305), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n351), .A2(new_n323), .A3(new_n329), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n279), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n343), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n345), .A2(new_n346), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(G472), .A2(G902), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT32), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n355), .A2(KEYINPUT73), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT73), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n334), .A2(new_n344), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT31), .ZN(new_n361));
  INV_X1    g175(.A(new_n343), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT28), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n337), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n311), .A2(KEYINPUT28), .A3(new_n336), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n331), .A2(new_n336), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n362), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n334), .A2(new_n335), .A3(new_n344), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n361), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n357), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n359), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n358), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n343), .B1(new_n366), .B2(new_n367), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n334), .A2(new_n362), .A3(new_n337), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n337), .A2(KEYINPUT72), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n311), .A2(new_n336), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT72), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n311), .A2(new_n381), .A3(new_n336), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n348), .B1(new_n383), .B2(KEYINPUT28), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n343), .A2(KEYINPUT29), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n378), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n370), .A2(new_n356), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT32), .ZN(new_n390));
  AOI22_X1  g204(.A1(G472), .A2(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n259), .B1(new_n373), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT9), .B(G234), .ZN(new_n393));
  OAI21_X1  g207(.A(G221), .B1(new_n393), .B2(G902), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(KEYINPUT80), .ZN(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT3), .B1(new_n396), .B2(G107), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n398));
  INV_X1    g212(.A(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(G104), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(G107), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G101), .ZN(new_n403));
  INV_X1    g217(.A(G101), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n397), .A2(new_n400), .A3(new_n404), .A4(new_n401), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(KEYINPUT4), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n404), .A2(KEYINPUT4), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT81), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n402), .A2(KEYINPUT81), .A3(new_n407), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n406), .B(new_n310), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT10), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n396), .A2(G107), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n399), .A2(G104), .ZN(new_n413));
  OAI21_X1  g227(.A(G101), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n411), .B1(new_n316), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n415), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n290), .A2(KEYINPUT10), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n410), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n305), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n410), .A2(new_n416), .A3(new_n418), .A4(new_n351), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G110), .B(G140), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n234), .A2(G227), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n314), .A2(new_n315), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n428), .A2(new_n415), .A3(new_n285), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n415), .B1(new_n428), .B2(new_n285), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n305), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT12), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(KEYINPUT12), .B(new_n305), .C1(new_n429), .C2(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT82), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n421), .A2(new_n436), .A3(new_n425), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n421), .B2(new_n425), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n427), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G469), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n188), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT83), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n421), .A2(new_n425), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT82), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n435), .A3(new_n437), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n446), .B2(new_n427), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n441), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n435), .A2(new_n421), .ZN(new_n451));
  INV_X1    g265(.A(new_n444), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n451), .A2(new_n426), .B1(new_n452), .B2(new_n420), .ZN(new_n453));
  OAI21_X1  g267(.A(G469), .B1(new_n453), .B2(G902), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n395), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G214), .B1(G237), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G122), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT84), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT5), .A4(new_n264), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n261), .A2(G119), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT5), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n268), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n417), .A2(new_n272), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n265), .A2(new_n271), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n276), .A2(new_n277), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n402), .A2(G101), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n405), .A2(KEYINPUT4), .ZN(new_n470));
  OAI22_X1  g284(.A1(new_n467), .A2(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n409), .A2(new_n408), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n460), .B(new_n466), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT85), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n279), .B(new_n406), .C1(new_n408), .C2(new_n409), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n475), .A2(new_n476), .A3(new_n460), .A4(new_n466), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n234), .A2(G224), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n316), .A2(new_n192), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n309), .A2(G125), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n465), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n415), .B1(new_n489), .B2(new_n468), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n491), .A2(new_n464), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n405), .B(new_n414), .C1(new_n276), .C2(new_n277), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n459), .B(KEYINPUT8), .Z(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n483), .A2(new_n484), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n481), .A3(new_n480), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n488), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n188), .B1(new_n479), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n475), .A2(new_n466), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n504), .B2(new_n459), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n494), .A2(new_n489), .ZN(new_n506));
  INV_X1    g320(.A(new_n470), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n507), .A2(new_n403), .B1(new_n272), .B2(new_n278), .ZN(new_n508));
  INV_X1    g322(.A(new_n408), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n402), .A2(KEYINPUT81), .A3(new_n407), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n506), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n476), .B1(new_n512), .B2(new_n460), .ZN(new_n513));
  INV_X1    g327(.A(new_n477), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n505), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n486), .A2(new_n487), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n512), .A2(KEYINPUT6), .A3(new_n460), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AND4_X1   g332(.A1(KEYINPUT86), .A2(new_n515), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n478), .B2(new_n505), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT86), .B1(new_n520), .B2(new_n516), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n502), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(G210), .B1(G237), .B2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT86), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n520), .A2(KEYINPUT86), .A3(new_n516), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n523), .A3(new_n502), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n457), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT90), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT66), .B(G131), .Z(new_n534));
  INV_X1    g348(.A(G237), .ZN(new_n535));
  AND4_X1   g349(.A1(G143), .A2(new_n535), .A3(new_n234), .A4(G214), .ZN(new_n536));
  AOI21_X1  g350(.A(G143), .B1(new_n339), .B2(G214), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n534), .B(KEYINPUT88), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n234), .A3(G214), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n281), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n339), .A2(G143), .A3(G214), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT88), .B1(new_n543), .B2(new_n534), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT17), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n231), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT88), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n541), .A2(new_n298), .A3(new_n542), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n538), .A4(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n545), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(G113), .B(G122), .Z(new_n554));
  XOR2_X1   g368(.A(KEYINPUT89), .B(G104), .Z(new_n555));
  XOR2_X1   g369(.A(new_n554), .B(new_n555), .Z(new_n556));
  NAND2_X1  g370(.A1(new_n200), .A2(new_n203), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n199), .A2(G146), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(KEYINPUT18), .A2(G131), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n543), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n543), .A2(new_n560), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n556), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n549), .A2(new_n538), .A3(new_n551), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT19), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n199), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n201), .A2(KEYINPUT19), .ZN(new_n568));
  AOI21_X1  g382(.A(G146), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n230), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n563), .ZN(new_n573));
  INV_X1    g387(.A(new_n556), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n533), .B1(new_n564), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n556), .B1(new_n572), .B2(new_n563), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n549), .A2(new_n538), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n231), .B1(new_n578), .B2(KEYINPUT17), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n561), .A2(new_n562), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n579), .A2(new_n552), .B1(new_n559), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n577), .B1(new_n581), .B2(new_n556), .ZN(new_n582));
  NOR2_X1   g396(.A1(G475), .A2(G902), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI22_X1  g398(.A1(new_n576), .A2(KEYINPUT20), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n564), .A2(new_n575), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT20), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n586), .A2(new_n533), .A3(new_n587), .A4(new_n583), .ZN(new_n588));
  INV_X1    g402(.A(new_n564), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n556), .B1(new_n553), .B2(new_n563), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n188), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n585), .A2(new_n588), .B1(G475), .B2(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n187), .A2(G953), .A3(new_n393), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n281), .B2(G128), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n209), .A2(KEYINPUT92), .A3(G143), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n281), .A2(G128), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n598), .A2(new_n292), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G122), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G116), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(G116), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G107), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n399), .A3(new_n605), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g424(.A1(KEYINPUT91), .A2(KEYINPUT13), .ZN(new_n611));
  NAND2_X1  g425(.A1(KEYINPUT91), .A2(KEYINPUT13), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n599), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n598), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n611), .A2(new_n612), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n617), .A2(new_n599), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n598), .A2(new_n613), .A3(KEYINPUT93), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n610), .B1(new_n620), .B2(G134), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n292), .B1(new_n598), .B2(new_n599), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n608), .B1(new_n600), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT94), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n604), .B2(KEYINPUT14), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT14), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n603), .A2(KEYINPUT94), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n604), .A2(KEYINPUT14), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n625), .A2(new_n605), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n623), .B1(G107), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n594), .B1(new_n621), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(G107), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n632), .B(new_n608), .C1(new_n600), .C2(new_n622), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n620), .A2(G134), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n633), .B(new_n593), .C1(new_n634), .C2(new_n610), .ZN(new_n635));
  AOI21_X1  g449(.A(G902), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G478), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(KEYINPUT15), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  AOI211_X1 g454(.A(G902), .B(new_n638), .C1(new_n631), .C2(new_n635), .ZN(new_n641));
  NAND2_X1  g455(.A1(G234), .A2(G237), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(G952), .A3(new_n234), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(G902), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n234), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT21), .B(G898), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n640), .A2(new_n641), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n592), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n392), .A2(new_n455), .A3(new_n532), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G101), .ZN(G3));
  NAND2_X1  g466(.A1(KEYINPUT95), .A2(G472), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n370), .A2(new_n188), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n653), .B1(new_n370), .B2(new_n188), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n259), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n455), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n631), .A2(new_n635), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT33), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT33), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n631), .A2(new_n635), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n659), .A2(G478), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n637), .A2(new_n188), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n636), .B2(new_n637), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n592), .A2(new_n665), .A3(new_n648), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n523), .B1(new_n530), .B2(new_n502), .ZN(new_n667));
  AOI211_X1 g481(.A(new_n524), .B(new_n501), .C1(new_n528), .C2(new_n529), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n456), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n657), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT34), .B(G104), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  XNOR2_X1  g486(.A(new_n636), .B(new_n639), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n584), .B1(new_n564), .B2(new_n575), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n587), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n591), .A2(G475), .ZN(new_n676));
  INV_X1    g490(.A(new_n648), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n673), .A2(new_n675), .A3(new_n676), .A4(new_n677), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n457), .B(new_n678), .C1(new_n525), .C2(new_n531), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n455), .A3(new_n656), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT96), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT35), .B(G107), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  NOR2_X1   g497(.A1(new_n242), .A2(KEYINPUT36), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n241), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n248), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n247), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n592), .A3(new_n649), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n688), .A2(new_n654), .A3(new_n655), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n532), .A2(new_n689), .A3(new_n455), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT37), .B(G110), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  NAND2_X1  g506(.A1(new_n389), .A2(new_n390), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n384), .A2(new_n386), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n188), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT29), .B1(new_n374), .B2(new_n375), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT73), .B1(new_n355), .B2(new_n357), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n370), .A2(new_n359), .A3(new_n371), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n693), .A2(new_n697), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n645), .A2(G900), .A3(new_n234), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT97), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n643), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n673), .A2(new_n675), .A3(new_n676), .A4(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n687), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n455), .A2(new_n532), .A3(new_n700), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n209), .ZN(G30));
  NAND2_X1  g524(.A1(new_n525), .A2(new_n531), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT38), .Z(new_n712));
  AOI21_X1  g526(.A(new_n362), .B1(new_n334), .B2(new_n337), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n188), .B1(new_n383), .B2(new_n343), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n693), .A2(new_n698), .A3(new_n699), .A4(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n716), .A2(new_n707), .ZN(new_n717));
  INV_X1    g531(.A(new_n673), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n592), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n717), .A2(new_n456), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n705), .B(KEYINPUT39), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n455), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n712), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  INV_X1    g541(.A(new_n592), .ZN(new_n728));
  INV_X1    g542(.A(new_n665), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n705), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n707), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n532), .A2(new_n455), .A3(new_n700), .A4(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT98), .B(G146), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G48));
  NAND2_X1  g548(.A1(new_n440), .A2(new_n188), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n395), .B1(new_n735), .B2(G469), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n448), .A2(new_n440), .A3(new_n441), .A4(new_n188), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n448), .B1(new_n447), .B2(new_n441), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n736), .B(KEYINPUT99), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT99), .B1(new_n450), .B2(new_n736), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n669), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n392), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  OAI21_X1  g560(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT99), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n679), .A2(new_n392), .A3(new_n749), .A4(new_n739), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  AOI21_X1  g565(.A(new_n688), .B1(new_n373), .B2(new_n391), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n532), .A3(new_n749), .A4(new_n739), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT100), .B(G119), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G21));
  OAI21_X1  g569(.A(G472), .B1(new_n355), .B2(G902), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n361), .A2(new_n369), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n384), .A2(new_n343), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n356), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT101), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n247), .B2(new_n249), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT101), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(new_n749), .A3(new_n677), .A4(new_n739), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT102), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n711), .A2(new_n767), .A3(new_n456), .A4(new_n719), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n456), .B(new_n719), .C1(new_n667), .C2(new_n668), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT102), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n766), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n602), .ZN(G24));
  NAND3_X1  g586(.A1(new_n756), .A2(new_n687), .A3(new_n759), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n730), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n742), .A2(KEYINPUT103), .A3(new_n532), .A4(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n774), .A2(new_n532), .A3(new_n749), .A4(new_n739), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT103), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT32), .B1(new_n370), .B2(new_n356), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT107), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n355), .B2(new_n357), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n370), .A2(KEYINPUT106), .A3(new_n371), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n697), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n730), .B(new_n764), .C1(new_n783), .C2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n395), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n525), .A2(new_n531), .A3(new_n789), .A4(new_n456), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n737), .A2(new_n738), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n453), .A2(G469), .ZN(new_n792));
  NAND2_X1  g606(.A1(G469), .A2(G902), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT104), .Z(new_n794));
  OR2_X1    g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT105), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT105), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n792), .A2(new_n794), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n450), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n790), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n781), .B1(new_n788), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n730), .A2(KEYINPUT42), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n392), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(G131), .Z(G33));
  NAND2_X1  g620(.A1(new_n796), .A2(new_n799), .ZN(new_n807));
  INV_X1    g621(.A(new_n706), .ZN(new_n808));
  INV_X1    g622(.A(new_n790), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n392), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT108), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT108), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n800), .A2(new_n812), .A3(new_n392), .A4(new_n808), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G134), .ZN(G36));
  OR2_X1    g629(.A1(new_n453), .A2(KEYINPUT45), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n453), .A2(KEYINPUT45), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(G469), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT109), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n794), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n450), .B1(new_n820), .B2(KEYINPUT46), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(KEYINPUT46), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n395), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n721), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n711), .A2(new_n457), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n728), .A2(new_n665), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT43), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n829), .B(new_n687), .C1(new_n654), .C2(new_n655), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n827), .B1(new_n831), .B2(KEYINPUT44), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(KEYINPUT44), .B2(new_n831), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n825), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n294), .ZN(G39));
  INV_X1    g649(.A(KEYINPUT47), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT111), .B1(new_n824), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n823), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n789), .B1(new_n838), .B2(new_n821), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT47), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n824), .A2(new_n842), .A3(new_n836), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT110), .B1(new_n839), .B2(KEYINPUT47), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n837), .A2(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n259), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n700), .A2(new_n846), .A3(new_n730), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n826), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(KEYINPUT112), .B(G140), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n848), .B(new_n849), .ZN(G42));
  AND3_X1   g664(.A1(new_n829), .A2(new_n644), .A3(new_n765), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n791), .B1(G469), .B2(new_n735), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n852), .A2(new_n395), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n826), .B(new_n851), .C1(new_n845), .C2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n773), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n742), .A2(new_n644), .A3(new_n826), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n829), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n716), .A2(new_n259), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n728), .A2(new_n729), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n855), .A2(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n851), .A2(new_n712), .A3(new_n457), .A4(new_n742), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT50), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT117), .Z(new_n865));
  NAND3_X1  g679(.A1(new_n854), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT118), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n800), .A2(new_n774), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n675), .A2(new_n676), .ZN(new_n871));
  INV_X1    g685(.A(new_n705), .ZN(new_n872));
  NOR4_X1   g686(.A1(new_n707), .A2(new_n871), .A3(new_n673), .A4(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n826), .A2(new_n455), .A3(new_n700), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n814), .A2(new_n802), .A3(new_n876), .A4(new_n804), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT113), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n744), .A2(new_n750), .A3(new_n753), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n878), .B1(new_n879), .B2(new_n771), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT114), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n532), .A2(new_n455), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n700), .A2(new_n846), .A3(new_n650), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n690), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n728), .A2(new_n729), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n592), .A2(new_n673), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n648), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n532), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n657), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n881), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n887), .A2(new_n532), .A3(new_n656), .A4(new_n455), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n651), .A2(KEYINPUT114), .A3(new_n690), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n766), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n770), .A2(new_n768), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n742), .B(new_n392), .C1(new_n743), .C2(new_n679), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(KEYINPUT113), .A3(new_n753), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n880), .A2(new_n893), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n709), .B1(new_n775), .B2(new_n778), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n872), .A2(new_n395), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n716), .A2(new_n707), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n796), .B2(new_n799), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n903), .A2(new_n895), .A3(KEYINPUT115), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT115), .B1(new_n903), .B2(new_n895), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n900), .B(new_n732), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT52), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n770), .A2(new_n768), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n807), .A2(new_n717), .A3(new_n901), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n903), .A2(new_n895), .A3(KEYINPUT115), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(KEYINPUT52), .A3(new_n732), .A4(new_n900), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n877), .B(new_n899), .C1(new_n908), .C2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(KEYINPUT116), .A3(KEYINPUT53), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT116), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n908), .A2(new_n915), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n899), .A2(new_n877), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT53), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT53), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n917), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n879), .A2(new_n771), .A3(new_n922), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n893), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(new_n877), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT54), .B1(new_n919), .B2(new_n929), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n926), .A2(KEYINPUT54), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n864), .A2(new_n867), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n854), .A2(new_n862), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n764), .B1(new_n783), .B2(new_n787), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n858), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT48), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n851), .A2(new_n532), .A3(new_n742), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(G952), .A3(new_n234), .ZN(new_n938));
  INV_X1    g752(.A(new_n885), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(new_n860), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT119), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n869), .A2(new_n931), .A3(new_n933), .A4(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(G952), .A2(G953), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n852), .B(KEYINPUT49), .ZN(new_n946));
  INV_X1    g760(.A(new_n828), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n789), .A2(new_n456), .ZN(new_n948));
  NOR4_X1   g762(.A1(new_n947), .A2(new_n716), .A3(new_n764), .A4(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n946), .A2(new_n712), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n945), .A2(new_n950), .ZN(G75));
  NOR2_X1   g765(.A1(new_n234), .A2(G952), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n919), .A2(new_n929), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n188), .B1(new_n925), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT56), .B1(new_n955), .B2(G210), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n520), .B(new_n516), .ZN(new_n957));
  XOR2_X1   g771(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n953), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n956), .B2(new_n959), .ZN(G51));
  NAND2_X1  g775(.A1(new_n955), .A2(new_n819), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n440), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n794), .B(KEYINPUT57), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT121), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n930), .C1(new_n916), .C2(KEYINPUT53), .ZN(new_n967));
  INV_X1    g781(.A(new_n804), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n801), .A2(new_n968), .A3(new_n875), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n969), .A2(new_n814), .A3(new_n927), .A4(new_n893), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n908), .B2(new_n915), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT54), .B1(new_n924), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n966), .B1(new_n925), .B2(new_n930), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n965), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT122), .ZN(new_n976));
  INV_X1    g790(.A(new_n930), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT121), .B1(new_n977), .B2(new_n924), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n967), .A3(new_n972), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT122), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n980), .A3(new_n965), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n964), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n963), .B1(new_n982), .B2(KEYINPUT123), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n975), .A2(KEYINPUT122), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n980), .B1(new_n979), .B2(new_n965), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n440), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT123), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n952), .B1(new_n983), .B2(new_n988), .ZN(G54));
  NAND3_X1  g803(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n990), .A2(new_n582), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n582), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n991), .A2(new_n992), .A3(new_n952), .ZN(G60));
  AND2_X1   g807(.A1(new_n659), .A2(new_n661), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n663), .B(KEYINPUT59), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n994), .B1(new_n931), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n952), .B1(new_n979), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT124), .ZN(G63));
  NAND2_X1  g814(.A1(G217), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT60), .Z(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n924), .B2(new_n971), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT125), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n952), .B1(new_n1004), .B2(new_n685), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1005), .B1(new_n239), .B2(new_n1004), .ZN(new_n1006));
  AOI21_X1  g820(.A(KEYINPUT126), .B1(new_n1004), .B2(new_n685), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1007), .A2(KEYINPUT61), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1006), .B(new_n1008), .ZN(G66));
  INV_X1    g823(.A(G224), .ZN(new_n1010));
  OAI21_X1  g824(.A(G953), .B1(new_n647), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n899), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1011), .B1(new_n1012), .B2(G953), .ZN(new_n1013));
  INV_X1    g827(.A(new_n520), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1014), .B1(G898), .B2(new_n234), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1013), .B(new_n1015), .ZN(G69));
  AND2_X1   g830(.A1(new_n900), .A2(new_n732), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n726), .ZN(new_n1018));
  OR2_X1    g832(.A1(new_n1018), .A2(KEYINPUT62), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(KEYINPUT62), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n885), .A2(new_n886), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n826), .A2(new_n392), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1022), .A2(new_n722), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n834), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n848), .A2(new_n1019), .A3(new_n1020), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n234), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n312), .B1(new_n331), .B2(new_n333), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n567), .A2(new_n568), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n234), .A2(G900), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n895), .A2(new_n934), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n825), .B1(new_n833), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1033), .A2(new_n805), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n848), .A2(new_n814), .A3(new_n1017), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1031), .B1(new_n1035), .B2(new_n234), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1030), .B1(new_n1036), .B2(new_n1029), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n234), .B1(G227), .B2(G900), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1037), .B(new_n1038), .ZN(G72));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT63), .Z(new_n1041));
  XNOR2_X1  g855(.A(new_n1041), .B(KEYINPUT127), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1042), .B1(new_n1025), .B2(new_n899), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n713), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1042), .B1(new_n1035), .B2(new_n899), .ZN(new_n1045));
  INV_X1    g859(.A(new_n375), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1044), .A2(new_n1047), .A3(new_n953), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1041), .ZN(new_n1049));
  NOR3_X1   g863(.A1(new_n1046), .A2(new_n713), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1048), .B1(new_n926), .B2(new_n1050), .ZN(G57));
endmodule


