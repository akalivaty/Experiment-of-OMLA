//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  INV_X1    g030(.A(G2104), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n456), .A2(G2105), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n457), .A2(G101), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n460), .A2(new_n461), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT65), .A3(G137), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n458), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n471), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT68), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n467), .A2(new_n463), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(G124), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n487), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n464), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n468), .A2(KEYINPUT4), .A3(G138), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n486), .A2(G126), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT5), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT70), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n509), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  OAI211_X1 g090(.A(G62), .B(new_n508), .C1(new_n511), .C2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(G543), .B1(new_n512), .B2(new_n513), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT72), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n507), .B1(new_n520), .B2(new_n514), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT73), .A3(G62), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n518), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT6), .B(G651), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  AOI211_X1 g102(.A(new_n507), .B(new_n527), .C1(new_n520), .C2(new_n514), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n527), .A2(new_n505), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G50), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n525), .A2(new_n533), .A3(KEYINPUT74), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  INV_X1    g111(.A(new_n523), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n516), .B2(new_n517), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n536), .B1(new_n538), .B2(new_n522), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n535), .B1(new_n539), .B2(new_n532), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n534), .A2(new_n540), .ZN(G166));
  NAND3_X1  g116(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n530), .A2(G51), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT75), .B(G89), .Z(new_n548));
  NAND2_X1  g123(.A1(new_n528), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  AOI22_X1  g126(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n536), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n530), .A2(G52), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n521), .A2(new_n526), .ZN(new_n555));
  INV_X1    g130(.A(G90), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(G171));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n520), .A2(new_n514), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(new_n508), .ZN(new_n561));
  INV_X1    g136(.A(G56), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n560), .A2(G81), .A3(new_n508), .A4(new_n526), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n530), .A2(G43), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n566), .B1(new_n565), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  NAND4_X1  g147(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  NAND2_X1  g151(.A1(new_n530), .A2(G53), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n530), .A2(new_n579), .A3(G53), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n528), .A2(G91), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n581), .B(new_n582), .C1(new_n583), .C2(new_n536), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  INV_X1    g160(.A(G166), .ZN(G303));
  AOI22_X1  g161(.A1(new_n528), .A2(G87), .B1(G49), .B2(new_n530), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G288));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n521), .B2(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n590), .B1(new_n593), .B2(new_n536), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n521), .A2(G86), .A3(new_n526), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n526), .A2(G48), .A3(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  AOI211_X1 g175(.A(new_n600), .B(new_n507), .C1(new_n520), .C2(new_n514), .ZN(new_n601));
  OAI211_X1 g176(.A(KEYINPUT77), .B(G651), .C1(new_n601), .C2(new_n592), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n594), .A2(new_n599), .A3(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n536), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n530), .A2(G47), .ZN(new_n606));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n555), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n561), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n560), .A2(G92), .A3(new_n508), .A4(new_n526), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT79), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT10), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT79), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n521), .A2(new_n619), .A3(G92), .A4(new_n526), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n618), .B1(new_n617), .B2(new_n620), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n611), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n611), .B1(new_n624), .B2(G868), .ZN(G321));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(G299), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G168), .B2(new_n627), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(G168), .B2(new_n627), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  NAND2_X1  g207(.A1(new_n624), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n571), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n462), .A2(new_n457), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n486), .A2(G123), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n463), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  INV_X1    g219(.A(G135), .ZN(new_n645));
  OAI221_X1 g220(.A(new_n642), .B1(new_n643), .B2(new_n644), .C1(new_n491), .C2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n640), .A2(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(G2096), .ZN(new_n649));
  NAND4_X1  g224(.A1(new_n641), .A2(new_n647), .A3(new_n648), .A4(new_n649), .ZN(G156));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n654), .B(new_n660), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(G14), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n662), .ZN(G401));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT17), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n669), .B2(new_n667), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT80), .Z(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n669), .A3(new_n667), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n673), .A2(new_n669), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n668), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2096), .B(G2100), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT81), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT20), .Z(new_n693));
  NOR2_X1   g268(.A1(new_n686), .A2(new_n688), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n695), .A2(new_n691), .A3(new_n689), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n693), .B(new_n696), .C1(new_n691), .C2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT82), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n705));
  NAND2_X1  g280(.A1(G166), .A2(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G16), .B2(G22), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(KEYINPUT85), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(KEYINPUT85), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G1971), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(G288), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT33), .ZN(new_n716));
  INV_X1    g291(.A(G1976), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G6), .B(G305), .S(G16), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT32), .B(G1981), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT84), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n719), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G1971), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n708), .A2(new_n724), .A3(new_n709), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n711), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(KEYINPUT34), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n486), .A2(G119), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n463), .A2(G107), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n730));
  INV_X1    g305(.A(G131), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n728), .B1(new_n729), .B2(new_n730), .C1(new_n491), .C2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(G25), .B(new_n732), .S(G29), .Z(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n712), .A2(G24), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT83), .Z(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G290), .B2(G16), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G1986), .Z(new_n740));
  NOR3_X1   g315(.A1(new_n727), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n726), .A2(KEYINPUT34), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n705), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n705), .A3(new_n742), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G27), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G164), .B2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(G2078), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n750), .A2(KEYINPUT94), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n746), .A2(G32), .ZN(new_n752));
  INV_X1    g327(.A(new_n491), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G141), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT26), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n457), .A2(G105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT93), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n756), .B(new_n758), .C1(G129), .C2(new_n486), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n752), .B1(new_n760), .B2(new_n746), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT27), .B(G1996), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n750), .A2(KEYINPUT94), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT31), .B(G11), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n766), .A2(G28), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n746), .B1(new_n766), .B2(G28), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n765), .B1(new_n767), .B2(new_n768), .C1(new_n646), .C2(new_n746), .ZN(new_n769));
  NOR4_X1   g344(.A1(new_n751), .A2(new_n763), .A3(new_n764), .A4(new_n769), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(new_n463), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT89), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n753), .A2(G139), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n775));
  NAND3_X1  g350(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n773), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT90), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(new_n746), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n746), .B2(G33), .ZN(new_n781));
  INV_X1    g356(.A(G2072), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n712), .A2(G21), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G168), .B2(new_n712), .ZN(new_n785));
  INV_X1    g360(.A(G1966), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G34), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(KEYINPUT24), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n788), .B2(KEYINPUT24), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(KEYINPUT91), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(KEYINPUT91), .B2(new_n790), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n480), .B2(new_n746), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT92), .B(G2084), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n781), .B2(new_n782), .ZN(new_n796));
  AND4_X1   g371(.A1(new_n770), .A2(new_n783), .A3(new_n787), .A4(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT95), .B(KEYINPUT23), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n712), .A2(G20), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G299), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n712), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT96), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1956), .ZN(new_n804));
  NOR2_X1   g379(.A1(G29), .A2(G35), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G162), .B2(G29), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT29), .ZN(new_n807));
  INV_X1    g382(.A(G2090), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n712), .A2(G5), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G171), .B2(new_n712), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1961), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n746), .A2(G26), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT28), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n815));
  INV_X1    g390(.A(G116), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G2105), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n486), .B2(G128), .ZN(new_n818));
  INV_X1    g393(.A(G140), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n491), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT87), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n814), .B1(new_n822), .B2(new_n746), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G2067), .ZN(new_n824));
  AOI211_X1 g399(.A(new_n812), .B(new_n824), .C1(new_n793), .C2(new_n794), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n797), .A2(new_n804), .A3(new_n809), .A4(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT97), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n624), .A2(G16), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G4), .B2(G16), .ZN(new_n829));
  INV_X1    g404(.A(G1348), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n712), .A2(G19), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT86), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n571), .B2(new_n712), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G1341), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n831), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  OR3_X1    g413(.A1(new_n826), .A2(new_n827), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n827), .B1(new_n826), .B2(new_n838), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n744), .A2(new_n745), .B1(new_n839), .B2(new_n840), .ZN(G311));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  INV_X1    g417(.A(new_n745), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n743), .B2(new_n843), .ZN(G150));
  NOR2_X1   g419(.A1(new_n623), .A2(new_n631), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT38), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n847));
  INV_X1    g422(.A(G67), .ZN(new_n848));
  AOI211_X1 g423(.A(new_n848), .B(new_n507), .C1(new_n520), .C2(new_n514), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n847), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n560), .A2(G67), .A3(new_n508), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n853), .A2(KEYINPUT98), .A3(new_n850), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(G651), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n528), .A2(G93), .B1(G55), .B2(new_n530), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n570), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n565), .A2(new_n567), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT76), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n862), .A2(new_n564), .A3(new_n855), .A4(new_n856), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n846), .B(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n866), .A2(new_n867), .A3(G860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n857), .A2(G860), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT99), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  OR2_X1    g446(.A1(new_n868), .A2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(G160), .B(G162), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n646), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n486), .A2(G130), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n463), .A2(G118), .ZN(new_n876));
  OAI21_X1  g451(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n877));
  INV_X1    g452(.A(G142), .ZN(new_n878));
  OAI221_X1 g453(.A(new_n875), .B1(new_n876), .B2(new_n877), .C1(new_n491), .C2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n638), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(new_n732), .Z(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(KEYINPUT100), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n822), .B(G164), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n760), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n822), .B(new_n501), .ZN(new_n885));
  INV_X1    g460(.A(new_n760), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n779), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(new_n887), .A3(new_n778), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n882), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(KEYINPUT100), .A3(new_n881), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n881), .A2(KEYINPUT100), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n882), .A2(new_n889), .A3(new_n893), .A4(new_n890), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n874), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(G37), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n874), .A3(new_n894), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n897), .A2(KEYINPUT101), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(KEYINPUT101), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g476(.A(new_n633), .B(new_n864), .Z(new_n902));
  NAND2_X1  g477(.A1(new_n623), .A2(new_n801), .ZN(new_n903));
  OAI211_X1 g478(.A(G299), .B(new_n615), .C1(new_n621), .C2(new_n622), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n617), .A2(new_n620), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT10), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G299), .B1(new_n912), .B2(new_n615), .ZN(new_n913));
  INV_X1    g488(.A(new_n904), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT103), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n902), .A2(new_n908), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n905), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n903), .A2(KEYINPUT102), .A3(new_n904), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n918), .B(KEYINPUT104), .C1(new_n902), .C2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(KEYINPUT104), .B2(new_n918), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n595), .A2(new_n598), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n521), .A2(G61), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n536), .B1(new_n927), .B2(new_n591), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n928), .B2(KEYINPUT77), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT105), .B1(new_n587), .B2(new_n588), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n521), .A2(G87), .A3(new_n526), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n530), .A2(G49), .ZN(new_n932));
  AND4_X1   g507(.A1(KEYINPUT105), .A2(new_n588), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n594), .B(new_n929), .C1(new_n930), .C2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n931), .A2(new_n932), .ZN(new_n936));
  INV_X1    g511(.A(new_n588), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n587), .A2(KEYINPUT105), .A3(new_n588), .ZN(new_n939));
  NAND3_X1  g514(.A1(G305), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n534), .A2(new_n540), .A3(G290), .ZN(new_n942));
  AOI21_X1  g517(.A(G290), .B1(new_n534), .B2(new_n540), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT74), .B1(new_n525), .B2(new_n533), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n539), .A2(new_n535), .A3(new_n532), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n609), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n534), .A2(new_n540), .A3(G290), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n940), .A4(new_n934), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n944), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT107), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n942), .A2(new_n941), .A3(new_n943), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n947), .A2(new_n948), .B1(new_n940), .B2(new_n934), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n944), .A2(new_n949), .A3(KEYINPUT106), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n952), .B1(new_n950), .B2(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n925), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n925), .A2(new_n959), .ZN(new_n961));
  OAI21_X1  g536(.A(G868), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n857), .A2(new_n627), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(G295));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n963), .ZN(G331));
  NOR2_X1   g540(.A1(new_n857), .A2(new_n570), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n862), .A2(new_n564), .B1(new_n855), .B2(new_n856), .ZN(new_n967));
  OAI21_X1  g542(.A(G171), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n858), .A2(new_n863), .A3(G301), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(G168), .A3(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n858), .A2(new_n863), .A3(G301), .ZN(new_n971));
  AOI21_X1  g546(.A(G301), .B1(new_n858), .B2(new_n863), .ZN(new_n972));
  OAI21_X1  g547(.A(G286), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n917), .A2(new_n908), .A3(new_n970), .A4(new_n973), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n971), .A2(new_n972), .A3(G286), .ZN(new_n975));
  AOI21_X1  g550(.A(G168), .B1(new_n968), .B2(new_n969), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n905), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n977), .A3(KEYINPUT108), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n975), .A2(new_n976), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n908), .A4(new_n917), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n958), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n973), .A2(new_n970), .B1(new_n921), .B2(new_n920), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n985), .A2(new_n986), .B1(new_n956), .B2(new_n957), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n915), .A2(new_n916), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(new_n973), .A3(new_n970), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT111), .B(new_n989), .C1(new_n979), .C2(new_n923), .ZN(new_n990));
  AOI21_X1  g565(.A(G37), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n984), .A2(new_n991), .A3(KEYINPUT112), .A4(new_n992), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n956), .B2(new_n957), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n978), .A2(new_n1000), .A3(new_n981), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n978), .B2(new_n981), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n1001), .A2(new_n1002), .A3(G37), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n998), .B1(new_n1003), .B2(new_n992), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1002), .A2(G37), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n1005), .C2(new_n1001), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n997), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n984), .A2(KEYINPUT43), .A3(new_n991), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT44), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(G397));
  INV_X1    g588(.A(G2067), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n822), .B(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n470), .A2(new_n471), .ZN(new_n1016));
  OAI211_X1 g591(.A(G40), .B(new_n479), .C1(new_n1016), .C2(new_n472), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT45), .B1(new_n501), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1015), .A2(KEYINPUT113), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT113), .B1(new_n1015), .B2(new_n1021), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1021), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n760), .B(G1996), .ZN(new_n1025));
  OAI22_X1  g600(.A1(new_n1022), .A2(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1026), .B(KEYINPUT114), .Z(new_n1027));
  XNOR2_X1  g602(.A(new_n732), .B(new_n734), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g604(.A(new_n609), .B(G1986), .Z(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1021), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G305), .A2(G1981), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G305), .A2(G1981), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1035), .ZN(new_n1039));
  INV_X1    g614(.A(G8), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1017), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n501), .A2(new_n1018), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT116), .B1(new_n501), .B2(new_n1018), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1040), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1038), .A2(new_n1039), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n717), .A3(new_n714), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1034), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1042), .A2(KEYINPUT50), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1041), .B(new_n1052), .C1(new_n1053), .C2(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1054), .B2(G2090), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n1018), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1020), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1041), .A2(KEYINPUT115), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1020), .A2(new_n1056), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1017), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n724), .A3(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n475), .A2(G40), .A3(new_n1052), .A4(new_n479), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1044), .A2(new_n1045), .A3(KEYINPUT50), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(KEYINPUT117), .A3(new_n808), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1055), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1067), .A2(G8), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1047), .B1(new_n717), .B2(G288), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT52), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n717), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1047), .B(new_n1077), .C1(new_n717), .C2(G288), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1048), .A2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1050), .A2(new_n1047), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G286), .A2(G8), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT51), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  XOR2_X1   g659(.A(new_n1056), .B(KEYINPUT119), .Z(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n1041), .C1(KEYINPUT45), .C2(new_n1046), .ZN(new_n1086));
  INV_X1    g661(.A(G2084), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1086), .A2(new_n786), .B1(new_n1065), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(G8), .B(new_n1084), .C1(new_n1089), .C2(G286), .ZN(new_n1090));
  OAI221_X1 g665(.A(new_n1082), .B1(new_n1083), .B2(KEYINPUT51), .C1(new_n1088), .C2(new_n1040), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1088), .A2(new_n1082), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1961), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1054), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n749), .A2(KEYINPUT53), .ZN(new_n1096));
  AOI21_X1  g671(.A(G2078), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1097));
  OAI221_X1 g672(.A(new_n1095), .B1(new_n1086), .B2(new_n1096), .C1(new_n1097), .C2(KEYINPUT53), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G171), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1093), .B1(KEYINPUT62), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1042), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT50), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1041), .B(new_n1103), .C1(new_n1046), .C2(new_n1102), .ZN(new_n1104));
  INV_X1    g679(.A(G1956), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1017), .A2(new_n1060), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1104), .A2(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n582), .B1(new_n583), .B2(new_n536), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n581), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(KEYINPUT122), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1113), .B2(G299), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT122), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1108), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n830), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1041), .A2(new_n1014), .A3(new_n1046), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n623), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1108), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1117), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT60), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT60), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n624), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT60), .B(new_n623), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1996), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1106), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1053), .B2(new_n1017), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n570), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1124), .A2(KEYINPUT61), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1108), .B(new_n1139), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1125), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1097), .A2(KEYINPUT53), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n1094), .B2(new_n1054), .ZN(new_n1144));
  XOR2_X1   g719(.A(G171), .B(KEYINPUT54), .Z(new_n1145));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n1146));
  AOI211_X1 g721(.A(new_n1096), .B(new_n1060), .C1(new_n1146), .C2(new_n1017), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1041), .A2(KEYINPUT125), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1145), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1144), .A2(new_n1149), .B1(new_n1098), .B2(new_n1145), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1100), .B1(new_n1142), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1098), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1152), .A2(new_n1090), .A3(new_n1092), .A4(new_n1091), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1062), .B1(new_n1104), .B2(G2090), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(G8), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1153), .A2(new_n1156), .A3(new_n1080), .A4(new_n1073), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1081), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1080), .A2(new_n1073), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1072), .B1(new_n1067), .B2(G8), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1089), .A2(G8), .A3(G168), .ZN(new_n1162));
  NOR4_X1   g737(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1156), .A2(new_n1073), .A3(new_n1048), .A4(new_n1079), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1164), .A2(KEYINPUT120), .A3(new_n1162), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1165), .A2(KEYINPUT63), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT120), .B1(new_n1164), .B2(new_n1162), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1163), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1031), .B1(new_n1158), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1021), .B1(new_n1015), .B2(new_n886), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1021), .A2(KEYINPUT46), .A3(new_n1131), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT46), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1024), .B2(G1996), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT47), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1024), .A2(G1986), .A3(G290), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT48), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1175), .B1(new_n1029), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n732), .A2(new_n735), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1027), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n822), .A2(new_n1014), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1024), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1169), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g759(.A1(new_n683), .A2(G319), .ZN(new_n1186));
  XOR2_X1   g760(.A(new_n1186), .B(KEYINPUT126), .Z(new_n1187));
  NOR3_X1   g761(.A1(G229), .A2(G401), .A3(new_n1187), .ZN(new_n1188));
  AND3_X1   g762(.A1(new_n1007), .A2(new_n900), .A3(new_n1188), .ZN(G308));
  NAND3_X1  g763(.A1(new_n1007), .A2(new_n900), .A3(new_n1188), .ZN(G225));
endmodule


