//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0004(.A(G50), .B1(G58), .B2(G68), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT64), .Z(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n211), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n210), .B(new_n214), .C1(new_n221), .C2(KEYINPUT1), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT2), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G226), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n227), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G87), .B(G97), .ZN(new_n234));
  INV_X1    g0034(.A(G107), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  INV_X1    g0037(.A(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  OAI21_X1  g0044(.A(new_n207), .B1(new_n211), .B2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n208), .A2(G33), .ZN(new_n247));
  OAI22_X1  g0047(.A1(new_n247), .A2(new_n202), .B1(new_n208), .B2(G68), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT74), .ZN(new_n249));
  OR2_X1    g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n248), .A2(new_n249), .B1(G50), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n246), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT11), .ZN(new_n254));
  INV_X1    g0054(.A(G68), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT70), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT70), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n259), .A2(new_n256), .A3(G13), .A4(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n261), .B(new_n246), .C1(G1), .C2(new_n208), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n262), .A2(KEYINPUT12), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n254), .B1(new_n255), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n258), .A2(new_n260), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(KEYINPUT12), .A3(new_n255), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n266), .B1(KEYINPUT12), .B2(new_n265), .C1(new_n253), .C2(KEYINPUT11), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT75), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT14), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT67), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G1), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT68), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n276), .A2(new_n281), .A3(new_n278), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n271), .B2(new_n275), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n280), .A2(new_n282), .B1(new_n285), .B2(G238), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT13), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OR2_X1    g0090(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G226), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G232), .A2(G1698), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G97), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n283), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n286), .A2(new_n287), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n287), .B1(new_n286), .B2(new_n298), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n270), .B(G169), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n301), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(G179), .A3(new_n299), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n299), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n270), .B1(new_n306), .B2(G169), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n269), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(G169), .B1(new_n300), .B2(new_n301), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT14), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n310), .A2(KEYINPUT75), .A3(new_n304), .A4(new_n302), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n268), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n268), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n303), .B2(new_n299), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n280), .A2(new_n282), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n285), .A2(G232), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n291), .A2(G223), .A3(new_n292), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G226), .A2(G1698), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n290), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G87), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n244), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n283), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(G200), .B1(new_n322), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n244), .ZN(new_n334));
  NAND2_X1  g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n332), .B1(new_n336), .B2(G20), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n255), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n208), .A2(new_n244), .ZN(new_n340));
  INV_X1    g0140(.A(G159), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT76), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT76), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n251), .A2(new_n343), .A3(G159), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(G58), .B(G68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G20), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n331), .B1(new_n339), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT7), .B1(new_n290), .B2(new_n208), .ZN(new_n350));
  NOR4_X1   g0150(.A1(new_n288), .A2(new_n289), .A3(new_n332), .A4(G20), .ZN(new_n351));
  OAI21_X1  g0151(.A(G68), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n342), .A2(new_n344), .B1(G20), .B2(new_n346), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(KEYINPUT16), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n349), .A2(new_n245), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT8), .B(G58), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n261), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n262), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(new_n357), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n328), .A2(new_n320), .A3(G190), .A4(new_n321), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n330), .A2(new_n355), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT17), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n362), .B(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(G169), .B1(new_n322), .B2(new_n329), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n328), .A2(new_n320), .A3(G179), .A4(new_n321), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n355), .A2(new_n360), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT18), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n364), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n207), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n244), .B2(new_n271), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n202), .B2(new_n290), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G223), .A2(G1698), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n291), .A2(new_n292), .ZN(new_n379));
  INV_X1    g0179(.A(G222), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n336), .B(new_n378), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n377), .A2(new_n381), .B1(G226), .B2(new_n285), .ZN(new_n382));
  INV_X1    g0182(.A(G179), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n383), .A3(new_n320), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n359), .A2(G50), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n251), .A2(G150), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n388), .B1(new_n201), .B2(new_n208), .C1(new_n356), .C2(new_n247), .ZN(new_n389));
  INV_X1    g0189(.A(G50), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n389), .A2(new_n245), .B1(new_n265), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n382), .A2(new_n320), .ZN(new_n393));
  INV_X1    g0193(.A(G169), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n386), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n385), .B2(new_n384), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n387), .A2(KEYINPUT9), .A3(new_n391), .ZN(new_n398));
  XOR2_X1   g0198(.A(new_n398), .B(KEYINPUT73), .Z(new_n399));
  NOR2_X1   g0199(.A1(new_n393), .A2(new_n313), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(G200), .B2(new_n393), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT9), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n392), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OR3_X1    g0204(.A1(new_n399), .A2(new_n404), .A3(KEYINPUT10), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT10), .B1(new_n399), .B2(new_n404), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n397), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n285), .A2(G244), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n320), .A2(new_n408), .ZN(new_n409));
  XOR2_X1   g0209(.A(KEYINPUT69), .B(G1698), .Z(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(G232), .A3(new_n336), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT72), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G238), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n334), .B2(new_n335), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(G1698), .B1(new_n290), .B2(G107), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n409), .B1(new_n417), .B2(new_n283), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n383), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G20), .A2(G77), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT15), .B(G87), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n420), .B1(new_n356), .B2(new_n340), .C1(new_n247), .C2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n245), .B1(new_n202), .B2(new_n265), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n202), .B2(new_n262), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n418), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n394), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n426), .B2(G200), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n418), .A2(G190), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n319), .A2(new_n374), .A3(new_n407), .A4(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT5), .B1(new_n272), .B2(new_n274), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT5), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n256), .B(G45), .C1(new_n435), .C2(G41), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n283), .A2(new_n277), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(KEYINPUT85), .A2(G294), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT85), .A2(G294), .ZN(new_n441));
  OAI21_X1  g0241(.A(G33), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(G257), .A2(G1698), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n288), .B2(new_n289), .ZN(new_n444));
  OAI21_X1  g0244(.A(G250), .B1(new_n288), .B2(new_n289), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n442), .B(new_n444), .C1(new_n445), .C2(new_n379), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n283), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n376), .B(G264), .C1(new_n434), .C2(new_n436), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n447), .A2(KEYINPUT86), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT86), .B1(new_n447), .B2(new_n448), .ZN(new_n450));
  OAI211_X1 g0250(.A(G179), .B(new_n439), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT87), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n447), .A2(new_n448), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT86), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n447), .A2(KEYINPUT86), .A3(new_n448), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n458), .A2(KEYINPUT87), .A3(G179), .A4(new_n439), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n447), .A2(new_n439), .A3(new_n448), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G169), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n453), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(new_n235), .A3(G20), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G116), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT84), .ZN(new_n467));
  OAI221_X1 g0267(.A(new_n464), .B1(G20), .B2(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n336), .A2(new_n208), .A3(G87), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n471), .A2(KEYINPUT22), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(KEYINPUT22), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT24), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT24), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n470), .B(new_n476), .C1(new_n472), .C2(new_n473), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n246), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n256), .A2(G33), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n261), .A2(new_n246), .A3(new_n479), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n480), .A2(new_n235), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT25), .B1(new_n261), .B2(G107), .ZN(new_n482));
  OR3_X1    g0282(.A1(new_n261), .A2(KEYINPUT25), .A3(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n462), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n449), .A2(new_n450), .ZN(new_n487));
  INV_X1    g0287(.A(new_n439), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n316), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n460), .A2(G190), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n478), .A2(new_n484), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n265), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n480), .B2(new_n495), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(G107), .B1(new_n350), .B2(new_n351), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  AND2_X1   g0300(.A1(G97), .A2(G107), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n235), .A2(KEYINPUT6), .A3(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n505), .A2(G20), .B1(G77), .B2(new_n251), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n246), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT77), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI211_X1 g0309(.A(KEYINPUT77), .B(new_n246), .C1(new_n499), .C2(new_n506), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n498), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g0312(.A(G244), .B1(new_n288), .B2(new_n289), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n379), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT78), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT78), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n512), .C1(new_n513), .C2(new_n379), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G244), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n334), .B2(new_n335), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(new_n410), .A3(KEYINPUT4), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n336), .A2(G250), .A3(G1698), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n283), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n437), .A2(new_n283), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n488), .B1(G257), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n383), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n376), .B1(new_n518), .B2(new_n524), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n527), .A2(G257), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n439), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n394), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n511), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n251), .A2(G77), .ZN(new_n535));
  INV_X1    g0335(.A(new_n504), .ZN(new_n536));
  XNOR2_X1  g0336(.A(G97), .B(G107), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n500), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n535), .B1(new_n538), .B2(new_n208), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n235), .B1(new_n337), .B2(new_n338), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n245), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT77), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n507), .A2(new_n508), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n497), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n526), .A2(G190), .A3(new_n528), .ZN(new_n545));
  OAI21_X1  g0345(.A(G200), .B1(new_n530), .B2(new_n532), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n534), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n265), .A2(new_n238), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n522), .B(new_n208), .C1(G33), .C2(new_n495), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n550), .B(new_n245), .C1(new_n208), .C2(G116), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT20), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n480), .A2(new_n238), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G264), .A2(G1698), .ZN(new_n558));
  INV_X1    g0358(.A(G257), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n336), .B(new_n558), .C1(new_n379), .C2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n560), .B(new_n283), .C1(G303), .C2(new_n336), .ZN(new_n561));
  OAI211_X1 g0361(.A(G270), .B(new_n376), .C1(new_n434), .C2(new_n436), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n439), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n557), .B(new_n564), .C1(new_n313), .C2(new_n563), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(G169), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n557), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n563), .A2(new_n383), .ZN(new_n569));
  OAI221_X1 g0369(.A(new_n549), .B1(new_n480), .B2(new_n238), .C1(new_n553), .C2(new_n554), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n570), .A2(KEYINPUT21), .A3(G169), .A4(new_n563), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n565), .A2(new_n568), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(G250), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n275), .B2(G1), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n256), .A2(new_n277), .A3(G45), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n376), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G238), .B1(new_n288), .B2(new_n289), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n465), .B1(new_n579), .B2(new_n379), .ZN(new_n580));
  OAI211_X1 g0380(.A(G244), .B(G1698), .C1(new_n288), .C2(new_n289), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT79), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT79), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n520), .A2(new_n583), .A3(G1698), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n580), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT80), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n283), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n415), .A2(new_n410), .B1(G33), .B2(G116), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n583), .B1(new_n520), .B2(G1698), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n581), .A2(KEYINPUT79), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n588), .B(new_n586), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n578), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n394), .ZN(new_n594));
  INV_X1    g0394(.A(new_n578), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n376), .B1(new_n596), .B2(KEYINPUT80), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n595), .B1(new_n597), .B2(new_n591), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n383), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT82), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n326), .A2(new_n495), .A3(new_n235), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n296), .A2(new_n208), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT19), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n208), .B(G68), .C1(new_n288), .C2(new_n289), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n247), .B2(new_n495), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n245), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n265), .A2(new_n421), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT81), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(KEYINPUT81), .A3(new_n609), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n480), .A2(new_n421), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n600), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n608), .A2(KEYINPUT81), .A3(new_n609), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT81), .B1(new_n608), .B2(new_n609), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n615), .B(new_n600), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n594), .B(new_n599), .C1(new_n616), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n593), .A2(G200), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n480), .A2(new_n326), .ZN(new_n623));
  XOR2_X1   g0423(.A(new_n623), .B(KEYINPUT83), .Z(new_n624));
  NAND2_X1  g0424(.A1(new_n596), .A2(KEYINPUT80), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n283), .A3(new_n591), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(G190), .A3(new_n578), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n622), .A2(new_n614), .A3(new_n624), .A4(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n548), .A2(new_n574), .A3(new_n621), .A4(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n433), .A2(new_n494), .A3(new_n629), .ZN(G372));
  XNOR2_X1  g0430(.A(new_n362), .B(KEYINPUT17), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n428), .A2(new_n318), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n312), .B2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n371), .B1(new_n367), .B2(new_n368), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n405), .A2(new_n406), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n397), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n621), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n511), .A2(new_n529), .A3(new_n533), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n621), .A2(new_n641), .A3(new_n628), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n621), .A2(new_n641), .A3(new_n628), .A4(KEYINPUT26), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND4_X1   g0446(.A1(new_n534), .A2(new_n621), .A3(new_n547), .A4(new_n628), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT88), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n451), .A2(new_n452), .B1(G169), .B2(new_n460), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n492), .B1(new_n649), .B2(new_n459), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n651), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n486), .A2(KEYINPUT88), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n647), .A2(new_n652), .A3(new_n654), .A4(new_n493), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n646), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n639), .B1(new_n433), .B2(new_n656), .ZN(G369));
  NAND3_X1  g0457(.A1(new_n256), .A2(new_n208), .A3(G13), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  XOR2_X1   g0459(.A(new_n659), .B(KEYINPUT89), .Z(new_n660));
  INV_X1    g0460(.A(G213), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n658), .B2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n486), .B(new_n493), .C1(new_n492), .C2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n650), .A2(new_n665), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n666), .A2(new_n557), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n651), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n573), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G330), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n494), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n653), .A2(new_n665), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n677), .A2(new_n678), .B1(new_n650), .B2(new_n666), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n212), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n272), .A2(new_n274), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n601), .A2(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n205), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT90), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT91), .B1(new_n593), .B2(new_n487), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n530), .A2(new_n532), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT91), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n458), .A2(new_n626), .A3(new_n693), .A4(new_n578), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n691), .A2(new_n569), .A3(new_n692), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT92), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  INV_X1    g0497(.A(new_n569), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n458), .A2(new_n626), .A3(new_n578), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(KEYINPUT91), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(new_n692), .A4(new_n694), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n530), .A2(new_n532), .A3(new_n697), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n691), .A2(new_n569), .A3(new_n694), .A4(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT94), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n700), .A2(KEYINPUT94), .A3(new_n694), .A4(new_n704), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT93), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n563), .A2(new_n383), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n598), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n593), .A2(KEYINPUT93), .A3(new_n383), .A4(new_n563), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n458), .A2(new_n439), .B1(new_n526), .B2(new_n528), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT95), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT95), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n712), .A2(new_n713), .A3(new_n717), .A4(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n703), .A2(new_n709), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n665), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n703), .A2(new_n709), .A3(new_n715), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n666), .A2(new_n722), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n629), .A2(new_n494), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n666), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n690), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n486), .A2(new_n653), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n647), .A2(new_n493), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n665), .B1(new_n646), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n665), .B1(new_n646), .B2(new_n655), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(KEYINPUT29), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n729), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n689), .B1(new_n737), .B2(G1), .ZN(G364));
  INV_X1    g0538(.A(new_n673), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n690), .ZN(new_n740));
  INV_X1    g0540(.A(G13), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G45), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n684), .A2(G1), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n674), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT96), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n207), .B1(G20), .B2(new_n394), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT98), .Z(new_n752));
  NOR2_X1   g0552(.A1(new_n681), .A2(new_n336), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n275), .B2(new_n206), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(KEYINPUT97), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(G45), .B2(new_n242), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n755), .A2(KEYINPUT97), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n681), .A2(new_n290), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n760), .A2(G355), .B1(new_n238), .B2(new_n681), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n752), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n750), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n208), .B1(new_n764), .B2(G190), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n495), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n313), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n767), .B1(new_n770), .B2(new_n390), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n768), .A2(G190), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n771), .B1(G68), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n208), .A2(G190), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(new_n383), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT99), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G107), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n774), .A2(new_n764), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n341), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n208), .A2(new_n313), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n383), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G58), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n774), .A2(new_n786), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n202), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n785), .A2(new_n383), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n326), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n790), .A2(new_n792), .A3(new_n290), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n773), .A2(new_n781), .A3(new_n784), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n780), .A2(G283), .ZN(new_n795));
  INV_X1    g0595(.A(G303), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n290), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G326), .B2(new_n769), .ZN(new_n798));
  INV_X1    g0598(.A(new_n765), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n440), .A2(new_n441), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n799), .A2(new_n801), .B1(new_n772), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n787), .A2(new_n804), .B1(new_n789), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n782), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G329), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n795), .A2(new_n798), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n763), .B1(new_n794), .B2(new_n809), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n762), .A2(new_n744), .A3(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT100), .Z(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n739), .B2(new_n749), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n746), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NOR2_X1   g0615(.A1(new_n750), .A2(new_n747), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n744), .B1(new_n202), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT101), .ZN(new_n818));
  INV_X1    g0618(.A(new_n772), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n767), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n780), .A2(G87), .ZN(new_n822));
  INV_X1    g0622(.A(new_n787), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G294), .A2(new_n823), .B1(new_n807), .B2(G311), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(new_n238), .C2(new_n789), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n821), .B(new_n825), .C1(G303), .C2(new_n769), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n290), .B1(new_n791), .B2(new_n235), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT102), .ZN(new_n828));
  INV_X1    g0628(.A(new_n789), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G143), .A2(new_n823), .B1(new_n829), .B2(G159), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  INV_X1    g0631(.A(G150), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n770), .B2(new_n831), .C1(new_n832), .C2(new_n819), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n779), .A2(new_n255), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n765), .A2(new_n788), .ZN(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n336), .B1(new_n782), .B2(new_n839), .C1(new_n791), .C2(new_n390), .ZN(new_n840));
  NOR4_X1   g0640(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n826), .A2(new_n828), .B1(new_n835), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n425), .A2(new_n427), .A3(new_n666), .ZN(new_n843));
  INV_X1    g0643(.A(new_n428), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n429), .A2(new_n430), .B1(new_n424), .B2(new_n665), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n818), .B1(new_n763), .B2(new_n842), .C1(new_n847), .C2(new_n748), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n734), .B(new_n847), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n729), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n744), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n729), .A2(new_n849), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(G384));
  NOR2_X1   g0653(.A1(new_n742), .A2(new_n256), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n308), .A2(new_n311), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n315), .ZN(new_n856));
  INV_X1    g0656(.A(new_n318), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n315), .A2(new_n665), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n855), .A2(new_n315), .A3(new_n665), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n846), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT40), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n368), .A2(KEYINPUT103), .ZN(new_n863));
  INV_X1    g0663(.A(new_n663), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT103), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n355), .A2(new_n865), .A3(new_n360), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n364), .B2(new_n373), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  INV_X1    g0670(.A(new_n362), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n355), .A2(new_n865), .A3(new_n360), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n865), .B1(new_n355), .B2(new_n360), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n871), .B1(new_n874), .B2(new_n367), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n870), .B1(new_n875), .B2(new_n867), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n368), .A2(new_n864), .ZN(new_n877));
  AND4_X1   g0677(.A1(new_n870), .A2(new_n369), .A3(new_n877), .A4(new_n362), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT38), .B(new_n869), .C1(new_n876), .C2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n369), .A2(new_n877), .A3(new_n362), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(new_n870), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n877), .B1(new_n631), .B2(new_n636), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n862), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n720), .A2(new_n725), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n726), .A2(new_n666), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT31), .B1(new_n720), .B2(new_n665), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n861), .B(new_n885), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT105), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n707), .A2(new_n708), .B1(new_n716), .B2(new_n718), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n666), .B1(new_n893), .B2(new_n703), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n886), .B(new_n887), .C1(new_n894), .C2(KEYINPUT31), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n895), .A2(KEYINPUT105), .A3(new_n861), .A4(new_n885), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n863), .A2(new_n367), .A3(new_n866), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n867), .A2(new_n898), .A3(new_n362), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n878), .B1(new_n899), .B2(KEYINPUT37), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n901), .A2(KEYINPUT104), .A3(KEYINPUT38), .A4(new_n869), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n867), .B1(new_n631), .B2(new_n636), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n880), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n879), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n895), .A2(new_n861), .A3(new_n902), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n862), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n720), .A2(new_n725), .B1(new_n726), .B2(new_n666), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n433), .B1(new_n723), .B2(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n897), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(new_n897), .B2(new_n908), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n911), .A2(new_n912), .A3(new_n690), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT106), .Z(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n859), .A2(new_n860), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n734), .A2(new_n847), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n918), .B2(new_n843), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n906), .A2(new_n902), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n919), .A2(new_n920), .B1(new_n373), .B2(new_n663), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n906), .A2(KEYINPUT39), .A3(new_n902), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n879), .A2(new_n884), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n312), .A2(new_n666), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n433), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n733), .B(new_n930), .C1(KEYINPUT29), .C2(new_n734), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n639), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n929), .B(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n854), .B1(new_n915), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n915), .B2(new_n933), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n936), .A2(G116), .A3(new_n209), .A4(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT36), .ZN(new_n939));
  OAI21_X1  g0739(.A(G77), .B1(new_n788), .B2(new_n255), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n940), .A2(new_n205), .B1(G50), .B2(new_n255), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G1), .A3(new_n741), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n935), .A2(new_n939), .A3(new_n942), .ZN(G367));
  NAND2_X1  g0743(.A1(new_n624), .A2(new_n614), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n665), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n621), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n621), .A2(new_n628), .A3(new_n945), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n749), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n751), .B1(new_n212), .B2(new_n421), .C1(new_n232), .C2(new_n754), .ZN(new_n953));
  INV_X1    g0753(.A(new_n744), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n780), .A2(G77), .ZN(new_n956));
  INV_X1    g0756(.A(new_n791), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n957), .A2(G58), .B1(new_n807), .B2(G137), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n956), .B(new_n958), .C1(new_n390), .C2(new_n789), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n765), .A2(new_n255), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n290), .B(new_n960), .C1(G150), .C2(new_n823), .ZN(new_n961));
  INV_X1    g0761(.A(G143), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n961), .B1(new_n962), .B2(new_n770), .C1(new_n341), .C2(new_n819), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n780), .A2(G97), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n336), .B1(new_n829), .B2(G283), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G303), .A2(new_n823), .B1(new_n807), .B2(G317), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n957), .A2(G116), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT46), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n967), .A2(new_n968), .B1(new_n772), .B2(new_n801), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n769), .A2(G311), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n235), .B2(new_n765), .C1(new_n967), .C2(new_n968), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n959), .A2(new_n963), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n955), .B1(new_n750), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n952), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n743), .A2(G1), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT111), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n669), .B2(new_n678), .ZN(new_n979));
  INV_X1    g0779(.A(new_n678), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n667), .A2(new_n980), .A3(KEYINPUT111), .A4(new_n668), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n674), .A2(KEYINPUT112), .B1(new_n677), .B2(new_n678), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n674), .A2(KEYINPUT112), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n984), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n979), .A2(new_n986), .A3(new_n981), .A4(new_n982), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n988), .A2(new_n729), .A3(new_n735), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT113), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n677), .A2(new_n678), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n650), .A2(new_n666), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n534), .B(new_n547), .C1(new_n544), .C2(new_n666), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n641), .A2(new_n665), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AND4_X1   g0796(.A1(KEYINPUT45), .A2(new_n992), .A3(new_n993), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT45), .B1(new_n679), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n992), .A2(new_n993), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n996), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1002), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n679), .B2(new_n996), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n675), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT45), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n679), .A2(KEYINPUT45), .A3(new_n996), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1011), .A2(new_n676), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n988), .A2(new_n729), .A3(KEYINPUT113), .A4(new_n735), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n991), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT114), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT114), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1013), .B1(new_n989), .B2(new_n990), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n1015), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n737), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n683), .B(KEYINPUT41), .Z(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n977), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n677), .A2(new_n996), .A3(new_n678), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT42), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n534), .B1(new_n994), .B2(new_n486), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n666), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT108), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT43), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1027), .A2(new_n1028), .B1(new_n666), .B2(new_n1030), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT43), .B1(new_n1036), .B2(KEYINPUT108), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1037), .A3(new_n950), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1035), .A2(new_n1037), .B1(new_n950), .B2(new_n1032), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1039), .A2(new_n1040), .A3(KEYINPUT109), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT109), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1032), .A2(new_n950), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1045), .B2(new_n1038), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1041), .A2(new_n1046), .B1(new_n676), .B2(new_n1001), .ZN(new_n1047));
  OAI21_X1  g0847(.A(KEYINPUT109), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1045), .A2(new_n1042), .A3(new_n1038), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n676), .A2(new_n1001), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n976), .B1(new_n1024), .B2(new_n1052), .ZN(G387));
  NAND2_X1  g0853(.A1(new_n989), .A2(new_n683), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n988), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1054), .A2(KEYINPUT115), .B1(new_n736), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(KEYINPUT115), .B2(new_n1054), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n670), .A2(new_n749), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n791), .A2(new_n800), .B1(new_n765), .B2(new_n820), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G317), .A2(new_n823), .B1(new_n829), .B2(G303), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n770), .B2(new_n804), .C1(new_n805), .C2(new_n819), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1061), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n779), .A2(new_n238), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n336), .B(new_n1068), .C1(G326), .C2(new_n807), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n765), .A2(new_n421), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n290), .B(new_n1071), .C1(G50), .C2(new_n823), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n357), .A2(new_n772), .B1(G159), .B2(new_n769), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n791), .A2(new_n202), .B1(new_n789), .B2(new_n255), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G150), .B2(new_n807), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n964), .A2(new_n1072), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n763), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n752), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n357), .A2(new_n390), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT50), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n685), .B(new_n275), .C1(new_n255), .C2(new_n202), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n753), .B1(new_n1080), .B2(new_n1081), .C1(new_n227), .C2(new_n275), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n760), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1082), .B1(G107), .B2(new_n212), .C1(new_n685), .C2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n744), .B(new_n1077), .C1(new_n1078), .C2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n988), .A2(new_n977), .B1(new_n1058), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1057), .A2(new_n1086), .ZN(G393));
  AOI21_X1  g0887(.A(new_n684), .B1(new_n1013), .B2(new_n989), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n239), .A2(new_n753), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n750), .B(new_n749), .C1(G97), .C2(new_n681), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n744), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n823), .A2(G311), .B1(G317), .B2(new_n769), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT52), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n336), .B1(new_n957), .B2(G283), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n829), .A2(G294), .B1(new_n807), .B2(G322), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n799), .A2(G116), .B1(G303), .B2(new_n772), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n781), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n290), .B1(new_n957), .B2(G68), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n789), .A2(new_n356), .B1(new_n782), .B2(new_n962), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n765), .A2(new_n202), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n772), .B2(G50), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n822), .A2(new_n1099), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n770), .A2(new_n832), .B1(new_n787), .B2(new_n341), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1094), .A2(new_n1098), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n750), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1092), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n1001), .B2(new_n749), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1014), .B2(new_n977), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1089), .A2(new_n1112), .ZN(G390));
  NAND2_X1  g0913(.A1(new_n918), .A2(new_n843), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n916), .B1(new_n728), .B2(new_n847), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n847), .A2(G330), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n895), .A2(new_n916), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1114), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n728), .A2(new_n847), .A3(new_n916), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n895), .A2(new_n1117), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n917), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n843), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n845), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n428), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n732), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1120), .A2(new_n1122), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1119), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n910), .A2(G330), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT117), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n910), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n932), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n665), .B(new_n846), .C1(new_n646), .C2(new_n655), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n916), .B1(new_n1135), .B2(new_n1123), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n925), .B1(new_n926), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n879), .A2(new_n884), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n926), .C1(new_n1126), .C2(new_n917), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1118), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n919), .A2(new_n927), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1139), .B(new_n1120), .C1(new_n1142), .C2(new_n925), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1134), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1128), .A2(new_n1141), .A3(new_n1133), .A4(new_n1143), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n683), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1141), .A2(new_n1143), .A3(new_n977), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n816), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n954), .B1(new_n357), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n837), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n819), .A2(new_n235), .B1(new_n770), .B2(new_n820), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1152), .A2(new_n792), .A3(new_n336), .A4(new_n1102), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n823), .A2(G116), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n829), .A2(G97), .B1(new_n807), .B2(G294), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT120), .Z(new_n1157));
  NOR2_X1   g0957(.A1(new_n765), .A2(new_n341), .ZN(new_n1158));
  INV_X1    g0958(.A(G125), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n787), .A2(new_n839), .B1(new_n782), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(G128), .C2(new_n769), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT54), .B(G143), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n819), .A2(new_n831), .B1(new_n789), .B2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT118), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n791), .A2(new_n832), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT53), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1161), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n336), .B1(new_n779), .B2(new_n390), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT119), .Z(new_n1169));
  OAI21_X1  g0969(.A(new_n1157), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1150), .B1(new_n1170), .B2(new_n750), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n925), .B2(new_n748), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1148), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT121), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT121), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1148), .A2(new_n1175), .A3(new_n1172), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1147), .A2(new_n1174), .A3(new_n1176), .ZN(G378));
  AOI21_X1  g0977(.A(new_n690), .B1(new_n907), .B2(new_n862), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n407), .B(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n392), .A2(new_n864), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n897), .A2(new_n1178), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n897), .B2(new_n1178), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n929), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n897), .A2(new_n1178), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1182), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n929), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n897), .A2(new_n1178), .A3(new_n1183), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1186), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1182), .A2(new_n747), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n954), .B1(G50), .B2(new_n1149), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n290), .A2(new_n272), .A3(new_n274), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G77), .B2(new_n957), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT122), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n770), .A2(new_n238), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n960), .B(new_n1198), .C1(G97), .C2(new_n772), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n780), .A2(G58), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n789), .A2(new_n421), .B1(new_n782), .B2(new_n820), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G107), .B2(new_n823), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT58), .ZN(new_n1204));
  AOI21_X1  g1004(.A(G50), .B1(new_n244), .B2(new_n271), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1203), .A2(new_n1204), .B1(new_n1195), .B2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n807), .C2(G124), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n770), .A2(new_n1159), .B1(new_n765), .B2(new_n832), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1162), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n957), .A2(new_n1209), .B1(new_n823), .B2(G128), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n831), .B2(new_n789), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1208), .B(new_n1211), .C1(G132), .C2(new_n772), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT59), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1207), .B1(new_n341), .B2(new_n779), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1212), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1206), .B1(new_n1204), .B2(new_n1203), .C1(new_n1214), .C2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1194), .B1(new_n1217), .B2(new_n750), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1192), .A2(new_n977), .B1(new_n1193), .B2(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1191), .A2(new_n1186), .B1(new_n1146), .B2(new_n1133), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n683), .B1(new_n1220), .B2(KEYINPUT57), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1146), .A2(new_n1133), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1192), .A2(KEYINPUT57), .A3(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1219), .B1(new_n1221), .B2(new_n1223), .ZN(G375));
  XNOR2_X1  g1024(.A(new_n1022), .B(KEYINPUT123), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n910), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT117), .B1(new_n910), .B2(G330), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n639), .B(new_n931), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n1119), .A3(new_n1127), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1226), .A2(new_n1230), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n336), .B(new_n1071), .C1(G97), .C2(new_n957), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G116), .A2(new_n772), .B1(new_n769), .B2(G294), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n787), .A2(new_n820), .B1(new_n782), .B2(new_n796), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G107), .B2(new_n829), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n956), .A2(new_n1232), .A3(new_n1233), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(G128), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n787), .A2(new_n831), .B1(new_n782), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G159), .B2(new_n957), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n336), .B1(new_n789), .B2(new_n832), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G50), .B2(new_n799), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1209), .A2(new_n772), .B1(G132), .B2(new_n769), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1200), .A2(new_n1239), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n763), .B1(new_n1236), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n954), .B1(G68), .B2(new_n1149), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n917), .C2(new_n747), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1128), .B2(new_n977), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1231), .A2(new_n1247), .ZN(G381));
  INV_X1    g1048(.A(new_n977), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1016), .A2(KEYINPUT114), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1019), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n736), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1249), .B1(new_n1252), .B2(new_n1022), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(G390), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n976), .A3(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1057), .A2(new_n814), .A3(new_n1086), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(new_n1257), .A2(G384), .A3(G381), .A4(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(G375), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1147), .A2(new_n1148), .A3(new_n1172), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(G407));
  NOR2_X1   g1062(.A1(new_n1259), .A2(new_n664), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1264));
  OAI21_X1  g1064(.A(G213), .B1(new_n1263), .B2(new_n1264), .ZN(G409));
  NAND2_X1  g1065(.A1(G393), .A2(G396), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1258), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1255), .A2(new_n976), .A3(new_n1256), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1256), .B1(new_n1255), .B2(new_n976), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1268), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G387), .A2(G390), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(new_n1257), .A3(new_n1267), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G378), .B(new_n1219), .C1(new_n1221), .C2(new_n1223), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1192), .A2(new_n1222), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(new_n1225), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1192), .A2(new_n977), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1193), .A2(new_n1218), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1261), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1275), .A2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n661), .A2(G343), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1229), .A2(KEYINPUT60), .A3(new_n1119), .A4(new_n1127), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1134), .A3(new_n683), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1128), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT60), .B1(new_n1287), .B2(new_n1229), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G384), .B(new_n1247), .C1(new_n1286), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT60), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1230), .A2(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1292), .A2(new_n683), .A3(new_n1134), .A4(new_n1285), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G384), .B1(new_n1293), .B2(new_n1247), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1284), .B1(new_n1290), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1247), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1296));
  INV_X1    g1096(.A(G384), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(KEYINPUT125), .A3(new_n1289), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1295), .A2(KEYINPUT62), .A3(new_n1299), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1282), .A2(new_n1283), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1295), .A2(new_n1299), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1283), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1275), .A2(KEYINPUT124), .A3(new_n1281), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT124), .B1(new_n1275), .B2(new_n1281), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1303), .B(new_n1304), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1301), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1298), .A2(new_n1289), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1283), .A2(G2897), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n1302), .B2(new_n1313), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1310), .B1(new_n1311), .B2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1274), .B1(new_n1309), .B2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1271), .A2(new_n1310), .A3(new_n1273), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT126), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1302), .A2(new_n1320), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1318), .A2(new_n1319), .B1(new_n1311), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1307), .A2(new_n1320), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1304), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1315), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1271), .A2(new_n1273), .A3(KEYINPUT126), .A4(new_n1310), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1322), .A2(new_n1323), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1317), .A2(new_n1328), .ZN(G405));
  NAND2_X1  g1129(.A1(G375), .A2(new_n1261), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT127), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(G375), .A2(KEYINPUT127), .A3(new_n1261), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(new_n1275), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1303), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1332), .A2(new_n1312), .A3(new_n1275), .A4(new_n1333), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1335), .A2(new_n1274), .A3(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1274), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


