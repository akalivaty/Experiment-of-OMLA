

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579;

  XNOR2_X1 U320 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n466) );
  XNOR2_X1 U321 ( .A(KEYINPUT38), .B(n452), .ZN(n500) );
  XOR2_X1 U322 ( .A(n470), .B(KEYINPUT28), .Z(n520) );
  XNOR2_X1 U323 ( .A(n346), .B(n363), .ZN(n517) );
  XOR2_X1 U324 ( .A(G218GAT), .B(G92GAT), .Z(n288) );
  XOR2_X1 U325 ( .A(n469), .B(KEYINPUT54), .Z(n289) );
  INV_X1 U326 ( .A(KEYINPUT101), .ZN(n333) );
  XNOR2_X1 U327 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U328 ( .A(n397), .B(n335), .ZN(n340) );
  XNOR2_X1 U329 ( .A(n471), .B(KEYINPUT119), .ZN(n472) );
  NOR2_X1 U330 ( .A1(n520), .A2(n540), .ZN(n525) );
  NOR2_X1 U331 ( .A1(n414), .A2(n576), .ZN(n415) );
  XNOR2_X1 U332 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U333 ( .A(n467), .B(n466), .ZN(n541) );
  XOR2_X1 U334 ( .A(n363), .B(n362), .Z(n526) );
  XNOR2_X1 U335 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n453) );
  XNOR2_X1 U337 ( .A(n479), .B(n478), .ZN(G1351GAT) );
  XNOR2_X1 U338 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n291) );
  XNOR2_X1 U340 ( .A(KEYINPUT84), .B(KEYINPUT14), .ZN(n290) );
  XNOR2_X1 U341 ( .A(n291), .B(n290), .ZN(n309) );
  XOR2_X1 U342 ( .A(G78GAT), .B(G64GAT), .Z(n293) );
  XNOR2_X1 U343 ( .A(G8GAT), .B(G1GAT), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U345 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n295) );
  XNOR2_X1 U346 ( .A(KEYINPUT15), .B(KEYINPUT82), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U348 ( .A(n297), .B(n296), .Z(n302) );
  XOR2_X1 U349 ( .A(KEYINPUT83), .B(G211GAT), .Z(n299) );
  NAND2_X1 U350 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U352 ( .A(G183GAT), .B(n300), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U354 ( .A(G22GAT), .B(G155GAT), .Z(n366) );
  XOR2_X1 U355 ( .A(n303), .B(n366), .Z(n307) );
  XOR2_X1 U356 ( .A(G15GAT), .B(G127GAT), .Z(n353) );
  XOR2_X1 U357 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n305) );
  XNOR2_X1 U358 ( .A(G71GAT), .B(G57GAT), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n422) );
  XNOR2_X1 U360 ( .A(n353), .B(n422), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n573) );
  XOR2_X1 U363 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n311) );
  XNOR2_X1 U364 ( .A(G141GAT), .B(KEYINPUT96), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n371) );
  XOR2_X1 U366 ( .A(n371), .B(G85GAT), .Z(n313) );
  XOR2_X1 U367 ( .A(G113GAT), .B(G1GAT), .Z(n442) );
  XNOR2_X1 U368 ( .A(G29GAT), .B(n442), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n326) );
  XOR2_X1 U370 ( .A(G155GAT), .B(G148GAT), .Z(n315) );
  XNOR2_X1 U371 ( .A(G162GAT), .B(G57GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U373 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n317) );
  XNOR2_X1 U374 ( .A(G127GAT), .B(KEYINPUT6), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U376 ( .A(n319), .B(n318), .Z(n324) );
  XOR2_X1 U377 ( .A(KEYINPUT100), .B(KEYINPUT1), .Z(n321) );
  NAND2_X1 U378 ( .A1(G225GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U380 ( .A(KEYINPUT4), .B(n322), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n331) );
  XOR2_X1 U383 ( .A(G120GAT), .B(G134GAT), .Z(n328) );
  XNOR2_X1 U384 ( .A(KEYINPUT0), .B(KEYINPUT87), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U386 ( .A(KEYINPUT88), .B(n329), .Z(n357) );
  INV_X1 U387 ( .A(n357), .ZN(n330) );
  XOR2_X1 U388 ( .A(n331), .B(n330), .Z(n390) );
  XNOR2_X1 U389 ( .A(G36GAT), .B(G190GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n288), .B(n332), .ZN(n397) );
  NAND2_X1 U391 ( .A1(G226GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U392 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n336), .B(KEYINPUT95), .ZN(n337) );
  XOR2_X1 U394 ( .A(n337), .B(KEYINPUT94), .Z(n339) );
  XNOR2_X1 U395 ( .A(G197GAT), .B(G204GAT), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n378) );
  XOR2_X1 U397 ( .A(n340), .B(n378), .Z(n342) );
  XOR2_X1 U398 ( .A(G169GAT), .B(G8GAT), .Z(n443) );
  XOR2_X1 U399 ( .A(G176GAT), .B(G64GAT), .Z(n423) );
  XNOR2_X1 U400 ( .A(n443), .B(n423), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U402 ( .A(KEYINPUT17), .B(G183GAT), .Z(n344) );
  XNOR2_X1 U403 ( .A(KEYINPUT19), .B(KEYINPUT90), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U405 ( .A(KEYINPUT18), .B(n345), .Z(n363) );
  XOR2_X1 U406 ( .A(KEYINPUT89), .B(KEYINPUT66), .Z(n348) );
  XNOR2_X1 U407 ( .A(G113GAT), .B(KEYINPUT91), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U409 ( .A(G176GAT), .B(G71GAT), .Z(n350) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(G43GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n361) );
  XOR2_X1 U413 ( .A(G190GAT), .B(G99GAT), .Z(n355) );
  XNOR2_X1 U414 ( .A(n353), .B(KEYINPUT20), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U416 ( .A(n357), .B(n356), .Z(n359) );
  NAND2_X1 U417 ( .A1(G227GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n362) );
  NAND2_X1 U420 ( .A1(n517), .A2(n526), .ZN(n381) );
  XOR2_X1 U421 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n365) );
  XNOR2_X1 U422 ( .A(KEYINPUT98), .B(KEYINPUT23), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n367) );
  XOR2_X1 U424 ( .A(n367), .B(n366), .Z(n369) );
  XNOR2_X1 U425 ( .A(G106GAT), .B(G218GAT), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U427 ( .A(G50GAT), .B(G162GAT), .Z(n396) );
  XOR2_X1 U428 ( .A(n370), .B(n396), .Z(n373) );
  XOR2_X1 U429 ( .A(G148GAT), .B(G78GAT), .Z(n429) );
  XNOR2_X1 U430 ( .A(n371), .B(n429), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U432 ( .A(KEYINPUT97), .B(KEYINPUT24), .Z(n375) );
  NAND2_X1 U433 ( .A1(G228GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U435 ( .A(n377), .B(n376), .Z(n380) );
  XNOR2_X1 U436 ( .A(n378), .B(KEYINPUT22), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n470) );
  NAND2_X1 U438 ( .A1(n381), .A2(n470), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n382), .B(KEYINPUT105), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n383), .B(KEYINPUT25), .ZN(n388) );
  XNOR2_X1 U441 ( .A(KEYINPUT104), .B(KEYINPUT26), .ZN(n385) );
  NOR2_X1 U442 ( .A1(n526), .A2(n470), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n563) );
  XNOR2_X1 U444 ( .A(n517), .B(KEYINPUT102), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n386), .B(KEYINPUT27), .ZN(n391) );
  NAND2_X1 U446 ( .A1(n563), .A2(n391), .ZN(n387) );
  NAND2_X1 U447 ( .A1(n388), .A2(n387), .ZN(n389) );
  NAND2_X1 U448 ( .A1(n390), .A2(n389), .ZN(n394) );
  INV_X1 U449 ( .A(n390), .ZN(n515) );
  NAND2_X1 U450 ( .A1(n391), .A2(n515), .ZN(n392) );
  XOR2_X1 U451 ( .A(KEYINPUT103), .B(n392), .Z(n540) );
  INV_X1 U452 ( .A(n526), .ZN(n475) );
  NAND2_X1 U453 ( .A1(n525), .A2(n475), .ZN(n393) );
  NAND2_X1 U454 ( .A1(n394), .A2(n393), .ZN(n484) );
  NAND2_X1 U455 ( .A1(n573), .A2(n484), .ZN(n395) );
  XOR2_X1 U456 ( .A(KEYINPUT109), .B(n395), .Z(n414) );
  XOR2_X1 U457 ( .A(KEYINPUT10), .B(n396), .Z(n399) );
  XNOR2_X1 U458 ( .A(n397), .B(G134GAT), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n405) );
  XNOR2_X1 U460 ( .A(G99GAT), .B(G85GAT), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n400), .B(G106GAT), .ZN(n418) );
  INV_X1 U462 ( .A(KEYINPUT67), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n418), .B(n401), .ZN(n403) );
  NAND2_X1 U464 ( .A1(G232GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U466 ( .A(n405), .B(n404), .Z(n413) );
  XOR2_X1 U467 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n407) );
  XNOR2_X1 U468 ( .A(G43GAT), .B(G29GAT), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U470 ( .A(KEYINPUT71), .B(n408), .Z(n439) );
  XOR2_X1 U471 ( .A(KEYINPUT79), .B(KEYINPUT11), .Z(n410) );
  XNOR2_X1 U472 ( .A(KEYINPUT9), .B(KEYINPUT65), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n439), .B(n411), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n552) );
  XNOR2_X1 U476 ( .A(n552), .B(KEYINPUT80), .ZN(n536) );
  XOR2_X1 U477 ( .A(KEYINPUT36), .B(n536), .Z(n576) );
  XNOR2_X1 U478 ( .A(KEYINPUT37), .B(n415), .ZN(n514) );
  XOR2_X1 U479 ( .A(G204GAT), .B(KEYINPUT33), .Z(n421) );
  XOR2_X1 U480 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n417) );
  XNOR2_X1 U481 ( .A(KEYINPUT31), .B(KEYINPUT77), .ZN(n416) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n435) );
  XOR2_X1 U485 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U486 ( .A1(G230GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n433) );
  XOR2_X1 U488 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n427) );
  XNOR2_X1 U489 ( .A(KEYINPUT73), .B(KEYINPUT78), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n428), .B(G92GAT), .ZN(n431) );
  XOR2_X1 U492 ( .A(G120GAT), .B(n429), .Z(n430) );
  XOR2_X1 U493 ( .A(n431), .B(n430), .Z(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U495 ( .A(n435), .B(n434), .Z(n569) );
  XOR2_X1 U496 ( .A(G197GAT), .B(G141GAT), .Z(n437) );
  XNOR2_X1 U497 ( .A(G15GAT), .B(KEYINPUT29), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n451) );
  XOR2_X1 U500 ( .A(G22GAT), .B(KEYINPUT70), .Z(n441) );
  XNOR2_X1 U501 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n447) );
  XOR2_X1 U503 ( .A(G50GAT), .B(G36GAT), .Z(n445) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U506 ( .A(n447), .B(n446), .Z(n449) );
  NAND2_X1 U507 ( .A1(G229GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n565) );
  INV_X1 U510 ( .A(n565), .ZN(n555) );
  NAND2_X1 U511 ( .A1(n569), .A2(n555), .ZN(n487) );
  NOR2_X1 U512 ( .A1(n514), .A2(n487), .ZN(n452) );
  NAND2_X1 U513 ( .A1(n500), .A2(n526), .ZN(n454) );
  XNOR2_X1 U514 ( .A(KEYINPUT41), .B(n569), .ZN(n455) );
  INV_X1 U515 ( .A(n455), .ZN(n544) );
  NOR2_X1 U516 ( .A1(n544), .A2(n565), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n456), .B(KEYINPUT46), .ZN(n457) );
  NOR2_X1 U518 ( .A1(n552), .A2(n457), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n458), .A2(n573), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n459), .B(KEYINPUT47), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n573), .A2(n576), .ZN(n461) );
  XNOR2_X1 U522 ( .A(KEYINPUT68), .B(KEYINPUT45), .ZN(n460) );
  XNOR2_X1 U523 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U524 ( .A1(n569), .A2(n462), .ZN(n463) );
  NOR2_X1 U525 ( .A1(n555), .A2(n463), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n465), .A2(n464), .ZN(n467) );
  XOR2_X1 U527 ( .A(n517), .B(KEYINPUT118), .Z(n468) );
  NOR2_X1 U528 ( .A1(n541), .A2(n468), .ZN(n469) );
  NOR2_X1 U529 ( .A1(n515), .A2(n289), .ZN(n564) );
  AND2_X1 U530 ( .A1(n470), .A2(n564), .ZN(n473) );
  INV_X1 U531 ( .A(KEYINPUT55), .ZN(n471) );
  NOR2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n560) );
  NAND2_X1 U533 ( .A1(n560), .A2(n536), .ZN(n479) );
  XOR2_X1 U534 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n477) );
  INV_X1 U535 ( .A(G190GAT), .ZN(n476) );
  INV_X1 U536 ( .A(n573), .ZN(n533) );
  NAND2_X1 U537 ( .A1(n560), .A2(n533), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(G183GAT), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(G1350GAT) );
  XNOR2_X1 U541 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n489) );
  NOR2_X1 U542 ( .A1(n536), .A2(n573), .ZN(n483) );
  XNOR2_X1 U543 ( .A(KEYINPUT16), .B(n483), .ZN(n485) );
  NAND2_X1 U544 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(KEYINPUT106), .ZN(n502) );
  NOR2_X1 U546 ( .A1(n502), .A2(n487), .ZN(n495) );
  NAND2_X1 U547 ( .A1(n495), .A2(n515), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(G1324GAT) );
  XOR2_X1 U549 ( .A(G8GAT), .B(KEYINPUT107), .Z(n491) );
  NAND2_X1 U550 ( .A1(n495), .A2(n517), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT108), .B(KEYINPUT35), .Z(n493) );
  NAND2_X1 U553 ( .A1(n495), .A2(n526), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G15GAT), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n495), .A2(n520), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  NAND2_X1 U559 ( .A1(n500), .A2(n515), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U561 ( .A1(n500), .A2(n517), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U563 ( .A1(n500), .A2(n520), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT110), .Z(n505) );
  NAND2_X1 U566 ( .A1(n565), .A2(n455), .ZN(n513) );
  NOR2_X1 U567 ( .A1(n502), .A2(n513), .ZN(n503) );
  XOR2_X1 U568 ( .A(KEYINPUT111), .B(n503), .Z(n510) );
  NAND2_X1 U569 ( .A1(n510), .A2(n515), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n507) );
  XOR2_X1 U571 ( .A(KEYINPUT42), .B(KEYINPUT112), .Z(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n517), .A2(n510), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n526), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n509), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U578 ( .A1(n510), .A2(n520), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n521), .A2(n515), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n517), .A2(n521), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n526), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n523) );
  NAND2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n541), .A2(n527), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n555), .A2(n537), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n530) );
  NAND2_X1 U596 ( .A1(n537), .A2(n455), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n532) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT114), .Z(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NAND2_X1 U600 ( .A1(n537), .A2(n533), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n563), .A2(n542), .ZN(n551) );
  NOR2_X1 U608 ( .A1(n565), .A2(n551), .ZN(n543) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  NOR2_X1 U610 ( .A1(n544), .A2(n551), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(KEYINPUT53), .B(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n573), .A2(n551), .ZN(n550) );
  XOR2_X1 U617 ( .A(G155GAT), .B(n550), .Z(G1346GAT) );
  INV_X1 U618 ( .A(n551), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n560), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n556), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n558) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(n559), .Z(n562) );
  NAND2_X1 U627 ( .A1(n560), .A2(n455), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n575) );
  NOR2_X1 U630 ( .A1(n565), .A2(n575), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n575), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n575), .ZN(n574) );
  XOR2_X1 U639 ( .A(G211GAT), .B(n574), .Z(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(G218GAT), .B(n579), .Z(G1355GAT) );
endmodule

