//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n594, new_n595,
    new_n596, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT67), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(new_n467), .A3(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  AND2_X1   g049(.A1(new_n465), .A2(new_n467), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT68), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n465), .A2(new_n467), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n463), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT69), .Z(new_n483));
  NOR2_X1   g058(.A1(new_n480), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n483), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND3_X1  g064(.A1(new_n475), .A2(G126), .A3(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT70), .B1(new_n463), .B2(G114), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n493), .A2(new_n494), .A3(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n491), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  AOI211_X1 g074(.A(KEYINPUT71), .B(new_n497), .C1(new_n492), .C2(new_n495), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n490), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n463), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n504), .B(KEYINPUT4), .ZN(new_n505));
  OAI211_X1 g080(.A(KEYINPUT72), .B(new_n490), .C1(new_n499), .C2(new_n500), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT73), .A3(G651), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(new_n513), .B1(KEYINPUT6), .B2(new_n510), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(G62), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n514), .A2(new_n521), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n517), .A2(new_n525), .ZN(G166));
  NAND2_X1  g101(.A1(new_n511), .A2(new_n513), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n527), .A2(G543), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n514), .B2(G543), .ZN(new_n532));
  OAI21_X1  g107(.A(G51), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n514), .A2(G89), .A3(new_n521), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n514), .A2(new_n531), .A3(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G52), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n510), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n527), .A2(new_n528), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n518), .A2(new_n520), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G90), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n544), .A2(new_n546), .A3(new_n550), .ZN(G171));
  NAND2_X1  g126(.A1(new_n543), .A2(G43), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n523), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n541), .B2(new_n542), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT75), .B1(new_n559), .B2(new_n555), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(new_n510), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  NAND4_X1  g146(.A1(new_n527), .A2(G53), .A3(G543), .A4(new_n528), .ZN(new_n572));
  AND2_X1   g147(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n574), .A2(new_n575), .B1(G91), .B2(new_n549), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n548), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n518), .A2(new_n520), .A3(KEYINPUT78), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n579), .A2(G65), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT77), .Z(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n577), .B1(new_n584), .B2(G651), .ZN(new_n585));
  AOI211_X1 g160(.A(KEYINPUT79), .B(new_n510), .C1(new_n581), .C2(new_n583), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n576), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n576), .B(KEYINPUT80), .C1(new_n585), .C2(new_n586), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G299));
  NAND3_X1  g166(.A1(new_n544), .A2(new_n546), .A3(new_n550), .ZN(G301));
  NAND3_X1  g167(.A1(new_n533), .A2(KEYINPUT81), .A3(new_n538), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(KEYINPUT81), .B1(new_n533), .B2(new_n538), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G286));
  OR2_X1    g172(.A1(new_n517), .A2(new_n525), .ZN(G303));
  NAND2_X1  g173(.A1(new_n549), .A2(G87), .ZN(new_n599));
  INV_X1    g174(.A(new_n529), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G49), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(G288));
  AOI22_X1  g178(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(new_n510), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n549), .A2(G86), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n600), .A2(G48), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(G305));
  XNOR2_X1  g183(.A(KEYINPUT82), .B(G47), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n541), .B2(new_n542), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G85), .ZN(new_n612));
  OAI22_X1  g187(.A1(new_n611), .A2(new_n510), .B1(new_n523), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n514), .A2(G92), .A3(new_n521), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT10), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n543), .A2(G54), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n579), .A2(G66), .A3(new_n580), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT83), .Z(new_n622));
  OAI21_X1  g197(.A(G651), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n618), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n616), .B1(new_n625), .B2(G868), .ZN(G321));
  XOR2_X1   g201(.A(G321), .B(KEYINPUT84), .Z(G284));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(G299), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(new_n596), .ZN(G297));
  OAI21_X1  g205(.A(new_n629), .B1(new_n628), .B2(new_n596), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n625), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g212(.A(new_n481), .ZN(new_n638));
  INV_X1    g213(.A(G123), .ZN(new_n639));
  OR3_X1    g214(.A1(new_n638), .A2(KEYINPUT85), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n484), .A2(G135), .ZN(new_n641));
  OR2_X1    g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n642), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n643));
  OAI21_X1  g218(.A(KEYINPUT85), .B1(new_n638), .B2(new_n639), .ZN(new_n644));
  NAND4_X1  g219(.A1(new_n640), .A2(new_n641), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT12), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT13), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n646), .A2(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2435), .ZN(new_n653));
  XOR2_X1   g228(.A(G2427), .B(G2438), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT14), .ZN(new_n656));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n661), .B(new_n662), .Z(new_n663));
  AND2_X1   g238(.A1(new_n663), .A2(G14), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2067), .B(G2678), .Z(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT17), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT86), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT87), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(G1986), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT22), .B(G1981), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  NAND2_X1  g272(.A1(new_n481), .A2(G129), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT94), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT96), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT26), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT95), .ZN(new_n705));
  AOI211_X1 g280(.A(new_n703), .B(new_n705), .C1(new_n484), .C2(G141), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n700), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n701), .B1(new_n700), .B2(new_n706), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G32), .B(new_n710), .S(G29), .Z(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT28), .ZN(new_n714));
  INV_X1    g289(.A(G26), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G29), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n484), .A2(G140), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n481), .A2(G128), .ZN(new_n721));
  OR2_X1    g296(.A1(G104), .A2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n722), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n717), .B1(new_n724), .B2(G29), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n716), .B1(new_n725), .B2(new_n714), .ZN(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G19), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n565), .B2(G16), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n726), .A2(G2067), .B1(G1341), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G2067), .B2(new_n726), .ZN(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G20), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT99), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT23), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G299), .B2(G16), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1956), .ZN(new_n736));
  NAND2_X1  g311(.A1(G171), .A2(G16), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G5), .B2(G16), .ZN(new_n738));
  INV_X1    g313(.A(G1961), .ZN(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G21), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G168), .B2(G16), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n738), .A2(new_n739), .B1(G1966), .B2(new_n741), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n736), .B(new_n742), .C1(G1341), .C2(new_n728), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT30), .B(G28), .Z(new_n744));
  OAI22_X1  g319(.A1(new_n741), .A2(G1966), .B1(G29), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G27), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G164), .B2(new_n746), .ZN(new_n748));
  MUX2_X1   g323(.A(new_n747), .B(new_n748), .S(KEYINPUT97), .Z(new_n749));
  AOI21_X1  g324(.A(new_n745), .B1(new_n749), .B2(G2078), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(G33), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n484), .A2(G139), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(new_n463), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT25), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n751), .B1(new_n758), .B2(new_n746), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT93), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G2072), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n645), .A2(new_n746), .ZN(new_n762));
  INV_X1    g337(.A(G34), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(KEYINPUT24), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(KEYINPUT24), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n746), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G160), .B2(new_n746), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G2084), .Z(new_n768));
  NAND4_X1  g343(.A1(new_n750), .A2(new_n761), .A3(new_n762), .A4(new_n768), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n730), .A2(new_n743), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n771));
  OAI22_X1  g346(.A1(new_n738), .A2(new_n739), .B1(new_n771), .B2(G11), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n760), .A2(G2072), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n772), .B(new_n773), .C1(new_n771), .C2(G11), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n625), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G4), .B2(G16), .ZN(new_n776));
  INV_X1    g351(.A(G1348), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AND4_X1   g353(.A1(new_n713), .A2(new_n770), .A3(new_n774), .A4(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n746), .A2(G25), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n481), .A2(G119), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n484), .A2(G131), .ZN(new_n782));
  OR2_X1    g357(.A1(G95), .A2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n783), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n780), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT35), .B(G1991), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n731), .A2(G24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n614), .B2(new_n731), .ZN(new_n790));
  INV_X1    g365(.A(G1986), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n731), .A2(G6), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n731), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT32), .B(G1981), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G22), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT90), .B1(new_n798), .B2(G16), .ZN(new_n799));
  OR3_X1    g374(.A1(new_n798), .A2(KEYINPUT90), .A3(G16), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n799), .B(new_n800), .C1(G166), .C2(new_n731), .ZN(new_n801));
  INV_X1    g376(.A(G1971), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT89), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G16), .B2(G23), .ZN(new_n805));
  OR3_X1    g380(.A1(new_n804), .A2(G16), .A3(G23), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n805), .B(new_n806), .C1(G288), .C2(new_n731), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT33), .B(G1976), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n797), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT88), .B(KEYINPUT34), .Z(new_n811));
  OAI211_X1 g386(.A(new_n788), .B(new_n792), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT91), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT36), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n814), .A2(new_n818), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n746), .A2(G35), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G162), .B2(new_n746), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2090), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n776), .A2(new_n777), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n779), .A2(new_n820), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n749), .A2(G2078), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n827), .A2(new_n829), .ZN(G311));
  OR2_X1    g405(.A1(new_n827), .A2(new_n829), .ZN(G150));
  AOI22_X1  g406(.A1(new_n543), .A2(G55), .B1(G93), .B2(new_n549), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(new_n510), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  AOI21_X1  g412(.A(new_n835), .B1(new_n561), .B2(new_n563), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n561), .A2(new_n563), .A3(new_n835), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n624), .A2(new_n632), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n837), .B1(new_n845), .B2(G860), .ZN(G145));
  INV_X1    g421(.A(G126), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n477), .A2(new_n847), .A3(new_n463), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n496), .A2(new_n498), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(KEYINPUT71), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n496), .A2(new_n491), .A3(new_n498), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n853), .A3(new_n505), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT4), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n504), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT100), .B1(new_n501), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n724), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n724), .A2(new_n858), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n700), .A2(new_n706), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT96), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n757), .B1(new_n862), .B2(new_n707), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n757), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n859), .B(new_n860), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n724), .B(new_n858), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n758), .B1(new_n708), .B2(new_n709), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n868), .A3(new_n864), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n481), .A2(G130), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n484), .A2(G142), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n874), .B(new_n875), .C1(G118), .C2(new_n463), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n870), .A2(new_n871), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n648), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n785), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n866), .A2(new_n869), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n866), .B2(new_n869), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n866), .A2(new_n869), .A3(KEYINPUT102), .A4(new_n879), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n645), .B(G160), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G162), .ZN(new_n887));
  AOI21_X1  g462(.A(G37), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(KEYINPUT103), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(new_n881), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(KEYINPUT103), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n880), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g469(.A1(new_n835), .A2(new_n628), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n841), .B(new_n634), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n589), .A2(new_n625), .A3(new_n590), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n625), .B1(new_n589), .B2(new_n590), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(G299), .A2(new_n624), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n899), .A2(new_n900), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(new_n896), .ZN(new_n907));
  NAND2_X1  g482(.A1(G303), .A2(KEYINPUT104), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n517), .A2(new_n525), .A3(KEYINPUT104), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(G305), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n912));
  NOR2_X1   g487(.A1(G166), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n794), .B1(new_n913), .B2(new_n909), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n614), .A2(G288), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n614), .A2(G288), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n915), .A2(KEYINPUT105), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  INV_X1    g495(.A(new_n918), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n916), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(KEYINPUT105), .A3(new_n918), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n914), .A4(new_n911), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT42), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n919), .A2(new_n924), .A3(KEYINPUT106), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT106), .B1(new_n919), .B2(new_n924), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n928), .B2(KEYINPUT42), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n907), .B(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n895), .B1(new_n930), .B2(new_n628), .ZN(G295));
  OAI21_X1  g506(.A(new_n895), .B1(new_n930), .B2(new_n628), .ZN(G331));
  NAND2_X1  g507(.A1(G168), .A2(G301), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n596), .B2(G301), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n839), .A2(new_n934), .A3(new_n840), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT81), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n539), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G301), .B1(new_n937), .B2(new_n593), .ZN(new_n938));
  NOR2_X1   g513(.A1(G171), .A2(new_n539), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n840), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n940), .B1(new_n941), .B2(new_n838), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n901), .A2(new_n903), .A3(new_n935), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT107), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n935), .A2(new_n942), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n901), .A4(new_n903), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n935), .A2(new_n942), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n906), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n944), .A2(new_n947), .A3(new_n928), .A4(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n943), .A2(new_n949), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n926), .B2(new_n927), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n950), .A2(new_n951), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n943), .A2(KEYINPUT107), .B1(new_n906), .B2(new_n948), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n928), .B1(new_n959), .B2(new_n947), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT43), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n950), .A2(new_n956), .A3(new_n954), .A4(new_n951), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT108), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n957), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n952), .A2(KEYINPUT43), .A3(new_n956), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n954), .B1(new_n958), .B2(new_n960), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(G397));
  AOI21_X1  g546(.A(G1384), .B1(new_n854), .B2(new_n857), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT109), .B(G40), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n470), .A2(new_n473), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n972), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT110), .Z(new_n977));
  XNOR2_X1  g552(.A(new_n724), .B(G2067), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n977), .B1(new_n978), .B2(new_n861), .ZN(new_n979));
  INV_X1    g554(.A(G1996), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT46), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n983), .B(KEYINPUT47), .Z(new_n984));
  NAND3_X1  g559(.A1(new_n977), .A2(G1996), .A3(new_n861), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(KEYINPUT111), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n710), .A2(new_n981), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n977), .B2(new_n978), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n785), .A2(new_n787), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n785), .A2(new_n787), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n977), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n985), .A2(KEYINPUT111), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n986), .A2(new_n988), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n976), .A2(new_n791), .A3(new_n614), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n994), .B(KEYINPUT48), .Z(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n986), .A2(new_n988), .A3(new_n989), .A4(new_n992), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G2067), .B2(new_n724), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n984), .B(new_n996), .C1(new_n977), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT63), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(G1384), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n507), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(new_n501), .B2(new_n856), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n974), .B1(new_n1004), .B2(KEYINPUT50), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1003), .A2(G2084), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n1002), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n975), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1966), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(G8), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1011), .A2(G286), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G303), .A2(G8), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n1015), .B(KEYINPUT55), .Z(new_n1016));
  AOI21_X1  g591(.A(new_n975), .B1(new_n972), .B2(KEYINPUT45), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n507), .A2(new_n1002), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n1008), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n802), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n507), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n974), .A3(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1024), .A2(G2090), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1016), .B1(new_n1026), .B2(G8), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n974), .B(new_n1002), .C1(new_n501), .C2(new_n856), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n599), .A2(new_n601), .A3(G1976), .A4(new_n602), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(G8), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(KEYINPUT112), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(KEYINPUT112), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(KEYINPUT52), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT114), .B(G1981), .Z(new_n1037));
  NOR2_X1   g612(.A1(G305), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1034), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G305), .A2(G1981), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(KEYINPUT49), .C1(G305), .C2(new_n1037), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1028), .A2(G8), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1044), .B1(new_n1047), .B2(new_n1030), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1042), .A2(KEYINPUT113), .A3(new_n1029), .A4(new_n1046), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1033), .A2(new_n1043), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1971), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1003), .A2(G2090), .A3(new_n1005), .ZN(new_n1053));
  OAI211_X1 g628(.A(G8), .B(new_n1016), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1027), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1000), .B1(new_n1014), .B2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1012), .B(KEYINPUT116), .ZN(new_n1058));
  OAI21_X1  g633(.A(G8), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1016), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1000), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1055), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1058), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT126), .ZN(new_n1065));
  INV_X1    g640(.A(G2078), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n858), .A2(KEYINPUT45), .A3(new_n1002), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1019), .A2(new_n1066), .A3(new_n974), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1018), .A2(KEYINPUT50), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1005), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT125), .B(G1961), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1068), .A2(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1007), .A2(new_n1066), .A3(new_n1009), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1007), .A2(KEYINPUT124), .A3(new_n1066), .A4(new_n1009), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(KEYINPUT53), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1065), .B1(new_n1080), .B2(G171), .ZN(new_n1081));
  AOI211_X1 g656(.A(KEYINPUT126), .B(G301), .C1(new_n1074), .C2(new_n1079), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n539), .A2(G8), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT122), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(new_n1086), .C1(new_n1006), .C2(new_n1010), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT51), .B1(new_n1085), .B2(KEYINPUT123), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1011), .A2(new_n1085), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n1011), .B2(new_n1085), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT62), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1027), .A2(new_n1055), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1091), .B(new_n1098), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1084), .A2(new_n1096), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G288), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1043), .A2(new_n1045), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1042), .B1(new_n1102), .B2(new_n1038), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1051), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(new_n1054), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT115), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1064), .A2(new_n1100), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1024), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1019), .A2(new_n974), .A3(new_n1067), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n587), .B(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1110), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1019), .A2(new_n980), .A3(new_n974), .A4(new_n1067), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1028), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1028), .A2(new_n1121), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT58), .B(G1341), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n565), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT59), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1130), .A3(new_n565), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1108), .A2(new_n1119), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1110), .A2(new_n1112), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1116), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1110), .A2(new_n1112), .A3(new_n1137), .A4(new_n1115), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1138), .A2(KEYINPUT61), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1118), .A2(KEYINPUT119), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n777), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1142));
  INV_X1    g717(.A(G2067), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1122), .A2(new_n1123), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1145), .A2(KEYINPUT120), .A3(new_n624), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT60), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT120), .B1(new_n1145), .B2(new_n624), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1147), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1154), .B2(new_n625), .ZN(new_n1155));
  OAI22_X1  g730(.A1(new_n1155), .A2(new_n1146), .B1(new_n1149), .B2(new_n1148), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1132), .A2(new_n1141), .A3(new_n1152), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1118), .A2(new_n625), .A3(new_n1148), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1136), .A2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1158), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n972), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1069), .B1(new_n1164), .B2(new_n1008), .ZN(new_n1165));
  INV_X1    g740(.A(G40), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n972), .B2(KEYINPUT45), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1165), .A2(new_n1066), .A3(new_n1167), .A4(G160), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1074), .A2(G301), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT54), .B1(new_n1083), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(G171), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1074), .A2(G301), .A3(new_n1079), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1174), .A2(KEYINPUT54), .A3(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1097), .A2(new_n1176), .A3(new_n1095), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT127), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1080), .A2(G171), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT126), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1080), .A2(new_n1065), .A3(G171), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(new_n1181), .A3(new_n1169), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT54), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1177), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1178), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1107), .B1(new_n1163), .B2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n614), .B(new_n791), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n976), .A2(new_n1190), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n993), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n999), .B1(new_n1189), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g768(.A(new_n461), .B1(new_n888), .B2(new_n892), .ZN(new_n1195));
  NOR2_X1   g769(.A1(G401), .A2(G227), .ZN(new_n1196));
  AND4_X1   g770(.A1(new_n696), .A2(new_n964), .A3(new_n1195), .A4(new_n1196), .ZN(G308));
  NAND4_X1  g771(.A1(new_n964), .A2(new_n1195), .A3(new_n696), .A4(new_n1196), .ZN(G225));
endmodule


