//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT64), .Z(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n209), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT0), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n203), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n207), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NOR4_X1   g0037(.A1(new_n224), .A2(new_n226), .A3(new_n230), .A4(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n234), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n255), .A2(KEYINPUT68), .A3(new_n234), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n207), .A3(G1), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT70), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT70), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n261), .A2(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n258), .A2(new_n264), .A3(new_n266), .A4(new_n259), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n263), .A2(new_n267), .B1(new_n206), .B2(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G50), .ZN(new_n269));
  OAI21_X1  g0069(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n270));
  INV_X1    g0070(.A(G150), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n207), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT8), .ZN(new_n274));
  OR3_X1    g0074(.A1(new_n274), .A2(new_n201), .A3(KEYINPUT69), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n274), .B1(new_n201), .B2(KEYINPUT69), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n207), .A2(G33), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n270), .B1(new_n271), .B2(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n279), .A2(new_n260), .B1(new_n217), .B2(new_n262), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT9), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n272), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G223), .A3(G1698), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G222), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n288), .B1(new_n219), .B2(new_n287), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G1), .A3(G13), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G274), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n297), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT67), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT67), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n294), .A2(new_n302), .A3(new_n297), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n296), .B(new_n299), .C1(new_n218), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n283), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n282), .A2(KEYINPUT9), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT10), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n311), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n306), .A2(new_n308), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(G200), .B2(new_n306), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n313), .A2(new_n314), .A3(new_n316), .A4(new_n283), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n306), .A2(G169), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n306), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n281), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n262), .A2(new_n256), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G1), .B2(new_n207), .ZN(new_n324));
  MUX2_X1   g0124(.A(new_n266), .B(new_n324), .S(G77), .Z(new_n325));
  XOR2_X1   g0125(.A(KEYINPUT8), .B(G58), .Z(new_n326));
  NOR2_X1   g0126(.A1(G20), .A2(G33), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n328), .B1(new_n207), .B2(new_n219), .C1(new_n329), .C2(new_n278), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n256), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n287), .A2(G238), .A3(G1698), .ZN(new_n333));
  INV_X1    g0133(.A(G107), .ZN(new_n334));
  INV_X1    g0134(.A(G232), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n333), .B1(new_n334), .B2(new_n287), .C1(new_n290), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n295), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n299), .C1(new_n220), .C2(new_n305), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(G190), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n332), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n332), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n338), .A2(new_n320), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n338), .A2(G169), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n318), .A2(new_n322), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n277), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(new_n266), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n268), .B2(new_n349), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT74), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G58), .A2(G68), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n207), .B1(new_n203), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G159), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n273), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n353), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(G58), .A2(G68), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G58), .A2(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(G20), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n327), .A2(G159), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(KEYINPUT74), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n285), .A2(new_n207), .A3(new_n286), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n286), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n202), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n352), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT77), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(KEYINPUT77), .B(new_n352), .C1(new_n364), .C2(new_n369), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n256), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n361), .A2(KEYINPUT74), .A3(new_n362), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT74), .B1(new_n361), .B2(new_n362), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n358), .A2(KEYINPUT75), .A3(new_n363), .ZN(new_n379));
  INV_X1    g0179(.A(new_n368), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT73), .ZN(new_n381));
  AND2_X1   g0181(.A1(KEYINPUT3), .A2(G33), .ZN(new_n382));
  NOR2_X1   g0182(.A1(KEYINPUT3), .A2(G33), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n285), .A2(KEYINPUT73), .A3(new_n286), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n207), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n380), .B1(new_n386), .B2(new_n366), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n378), .B(new_n379), .C1(new_n202), .C2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n351), .B1(new_n374), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n299), .B1(new_n300), .B2(new_n335), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n287), .A2(G226), .A3(G1698), .ZN(new_n393));
  INV_X1    g0193(.A(G223), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n393), .B1(new_n272), .B2(new_n211), .C1(new_n290), .C2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n392), .B1(new_n395), .B2(new_n295), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n320), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(G169), .B2(new_n396), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n391), .A2(new_n399), .A3(KEYINPUT18), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT78), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n376), .A2(new_n377), .A3(new_n375), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT75), .B1(new_n358), .B2(new_n363), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n387), .A2(new_n202), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT16), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n255), .A2(new_n234), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n370), .B2(new_n371), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n408), .A3(new_n373), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n398), .B1(new_n409), .B2(new_n351), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT78), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT18), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n391), .A2(new_n399), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n401), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n396), .A2(new_n308), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(G200), .B2(new_n396), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n409), .A2(new_n418), .A3(new_n351), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n348), .B1(KEYINPUT79), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(KEYINPUT79), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n304), .A2(G238), .B1(G274), .B2(new_n298), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n287), .A2(G226), .A3(new_n289), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G97), .ZN(new_n426));
  OAI211_X1 g0226(.A(G232), .B(G1698), .C1(new_n382), .C2(new_n383), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(KEYINPUT71), .A3(new_n295), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT72), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n295), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT71), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n430), .A2(new_n431), .A3(new_n432), .A4(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(new_n424), .A3(new_n432), .A4(new_n429), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT72), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n430), .A2(new_n435), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT13), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(G169), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n436), .A2(new_n438), .B1(new_n440), .B2(KEYINPUT13), .ZN(new_n445));
  INV_X1    g0245(.A(G169), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT14), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n441), .A2(G179), .A3(new_n437), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n265), .A2(G20), .A3(new_n202), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT12), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n327), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n219), .B2(new_n278), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n260), .A2(new_n453), .A3(KEYINPUT11), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n451), .B(new_n454), .C1(new_n202), .C2(new_n324), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT11), .B1(new_n260), .B2(new_n453), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n449), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n441), .A2(G190), .A3(new_n437), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n457), .C1(new_n445), .C2(new_n340), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n423), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n422), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT19), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n465), .A2(new_n207), .A3(G33), .A4(G97), .ZN(new_n466));
  NOR2_X1   g0266(.A1(G87), .A2(G97), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n467), .A2(new_n334), .B1(new_n426), .B2(new_n207), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n468), .B2(new_n465), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n287), .A2(KEYINPUT84), .A3(new_n207), .A4(G68), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n207), .B(G68), .C1(new_n382), .C2(new_n383), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT84), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n474), .A2(new_n256), .B1(new_n329), .B2(new_n262), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n206), .A2(G33), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n258), .A2(new_n266), .A3(new_n259), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n329), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(KEYINPUT85), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT85), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n477), .B2(new_n329), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  OAI21_X1  g0285(.A(G250), .B1(new_n485), .B2(G1), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n487));
  INV_X1    g0287(.A(new_n234), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n293), .ZN(new_n489));
  OAI211_X1 g0289(.A(G238), .B(new_n289), .C1(new_n382), .C2(new_n383), .ZN(new_n490));
  OAI211_X1 g0290(.A(G244), .B(G1698), .C1(new_n382), .C2(new_n383), .ZN(new_n491));
  INV_X1    g0291(.A(G116), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n272), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n489), .B1(new_n495), .B2(new_n295), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(G169), .ZN(new_n497));
  AOI211_X1 g0297(.A(G179), .B(new_n489), .C1(new_n495), .C2(new_n295), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n484), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n496), .A2(new_n320), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(KEYINPUT83), .C1(G169), .C2(new_n496), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n483), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n478), .A2(G87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n495), .A2(new_n295), .ZN(new_n504));
  INV_X1    g0304(.A(new_n489), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(G190), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n496), .A2(G200), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n475), .B(new_n503), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT86), .B1(new_n502), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT86), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n499), .A2(new_n501), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n509), .C1(new_n513), .C2(new_n483), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  AND2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G97), .A2(G107), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n334), .A2(KEYINPUT6), .A3(G97), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n521), .A2(new_n207), .B1(new_n219), .B2(new_n273), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n334), .B1(new_n367), .B2(new_n368), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n256), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT80), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n367), .A2(new_n368), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G107), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n519), .A2(new_n520), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(G20), .B1(G77), .B2(new_n327), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n407), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT80), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n477), .A2(G97), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n266), .A2(new_n213), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G1698), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n287), .A2(G244), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n382), .A2(new_n383), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(new_n220), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n537), .B(new_n540), .C1(new_n542), .C2(KEYINPUT4), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n287), .A2(G250), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n289), .B1(new_n544), .B2(KEYINPUT4), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n295), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT5), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT81), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(G41), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n485), .A2(G1), .ZN(new_n550));
  INV_X1    g0350(.A(G41), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G274), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(G257), .A3(new_n294), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n546), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n533), .A2(new_n536), .B1(new_n446), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n546), .A2(new_n320), .A3(new_n557), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT82), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n546), .A2(new_n562), .A3(new_n320), .A4(new_n557), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n525), .A2(new_n532), .B1(new_n535), .B2(new_n534), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n546), .A2(new_n308), .A3(new_n557), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n553), .A2(new_n294), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n555), .B1(new_n567), .B2(new_n214), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n541), .A2(new_n212), .ZN(new_n569));
  OAI21_X1  g0369(.A(G1698), .B1(new_n569), .B2(new_n538), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n287), .A2(G244), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n538), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n570), .A2(new_n537), .A3(new_n540), .A4(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n568), .B1(new_n573), .B2(new_n295), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n566), .B1(new_n574), .B2(G200), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n559), .A2(new_n564), .B1(new_n565), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(G250), .B(new_n289), .C1(new_n382), .C2(new_n383), .ZN(new_n577));
  OAI211_X1 g0377(.A(G257), .B(G1698), .C1(new_n382), .C2(new_n383), .ZN(new_n578));
  INV_X1    g0378(.A(G294), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n577), .B(new_n578), .C1(new_n272), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n295), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n553), .A2(G264), .A3(new_n294), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT88), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT88), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n553), .A2(new_n584), .A3(G264), .A4(new_n294), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n581), .A2(new_n583), .A3(new_n585), .A4(new_n555), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n340), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n580), .A2(new_n295), .B1(new_n582), .B2(KEYINPUT88), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n588), .A2(new_n308), .A3(new_n585), .A4(new_n555), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n265), .A2(G20), .A3(new_n334), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT25), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n591), .A2(KEYINPUT25), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(new_n593), .C1(new_n477), .C2(new_n334), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT23), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n207), .B2(G107), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n334), .A2(KEYINPUT23), .A3(G20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n493), .A2(new_n207), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n207), .B(G87), .C1(new_n382), .C2(new_n383), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT22), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT22), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n287), .A2(new_n603), .A3(new_n207), .A4(G87), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n605), .A2(KEYINPUT24), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n407), .B1(new_n605), .B2(KEYINPUT24), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n594), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n590), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT89), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT89), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n590), .A2(new_n611), .A3(new_n608), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n407), .A2(new_n266), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n476), .A2(G116), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n614), .A2(new_n615), .B1(G116), .B2(new_n266), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT20), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n207), .A2(new_n492), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n537), .B1(new_n213), .B2(G33), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(new_n207), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n617), .B1(new_n620), .B2(new_n407), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n272), .A2(G97), .ZN(new_n622));
  AOI21_X1  g0422(.A(G20), .B1(new_n622), .B2(new_n537), .ZN(new_n623));
  OAI211_X1 g0423(.A(KEYINPUT20), .B(new_n256), .C1(new_n623), .C2(new_n618), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n616), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(G264), .B(G1698), .C1(new_n382), .C2(new_n383), .ZN(new_n626));
  OAI211_X1 g0426(.A(G257), .B(new_n289), .C1(new_n382), .C2(new_n383), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n285), .A2(G303), .A3(new_n286), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n295), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n553), .A2(G270), .A3(new_n294), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n630), .A2(new_n555), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(G200), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(new_n555), .A3(new_n631), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(G190), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n625), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n621), .A2(new_n624), .ZN(new_n637));
  INV_X1    g0437(.A(new_n615), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n323), .A2(new_n638), .B1(new_n492), .B2(new_n262), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n632), .A2(new_n640), .A3(KEYINPUT87), .A4(G179), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT87), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n630), .A2(G179), .A3(new_n555), .A4(new_n631), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n625), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n640), .A2(KEYINPUT21), .A3(new_n634), .A4(G169), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n640), .A2(G169), .A3(new_n634), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT21), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n636), .A2(new_n645), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n586), .A2(G169), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n588), .A2(G179), .A3(new_n585), .A4(new_n555), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n594), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n605), .A2(KEYINPUT24), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n256), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n605), .A2(KEYINPUT24), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n576), .A2(new_n613), .A3(new_n651), .A4(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n464), .A2(new_n515), .A3(new_n661), .ZN(G372));
  NAND2_X1  g0462(.A1(new_n415), .A2(new_n400), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n449), .A2(new_n458), .B1(new_n346), .B2(new_n461), .ZN(new_n664));
  INV_X1    g0464(.A(new_n420), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n666), .A2(new_n318), .B1(new_n281), .B2(new_n321), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n464), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n497), .A2(new_n498), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n509), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(KEYINPUT90), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n672), .B2(new_n509), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n565), .A2(new_n575), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n660), .A2(new_n645), .A3(new_n646), .A4(new_n649), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n613), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n530), .A2(new_n531), .ZN(new_n681));
  AOI211_X1 g0481(.A(KEYINPUT80), .B(new_n407), .C1(new_n527), .C2(new_n529), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n536), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n558), .A2(new_n446), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n564), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n677), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n564), .A2(new_n683), .A3(new_n684), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n511), .A2(new_n687), .A3(new_n514), .ZN(new_n688));
  XNOR2_X1  g0488(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n686), .A2(KEYINPUT26), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n672), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n668), .B1(new_n669), .B2(new_n691), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT92), .Z(G369));
  INV_X1    g0493(.A(new_n265), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .A3(G20), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT27), .B1(new_n694), .B2(G20), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n660), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n699), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n613), .B1(new_n608), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n702), .B2(new_n660), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n645), .A2(new_n646), .A3(new_n649), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(new_n701), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n700), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n640), .A2(new_n699), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n650), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n704), .B2(new_n707), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n703), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n706), .A2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n227), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n467), .A2(new_n334), .A3(new_n492), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n715), .A2(new_n206), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n233), .B2(new_n715), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT28), .Z(new_n719));
  XNOR2_X1  g0519(.A(new_n673), .B(KEYINPUT90), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT26), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n685), .A2(new_n721), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n688), .A2(new_n689), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n685), .B1(new_n674), .B2(new_n676), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n672), .B1(new_n680), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(KEYINPUT29), .B(new_n701), .C1(new_n723), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n699), .B1(new_n690), .B2(new_n672), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(KEYINPUT29), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n685), .A2(new_n678), .A3(new_n660), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n650), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n511), .A2(new_n514), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n613), .A4(new_n701), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  INV_X1    g0533(.A(new_n643), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n588), .A2(KEYINPUT94), .A3(new_n496), .A4(new_n585), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n574), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n581), .A2(new_n583), .A3(new_n585), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT94), .B1(new_n737), .B2(new_n496), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n733), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n558), .A2(new_n643), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT94), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n588), .A2(new_n585), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(new_n742), .B2(new_n506), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n740), .A2(new_n743), .A3(KEYINPUT30), .A4(new_n735), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n496), .A2(G179), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n558), .A2(new_n586), .A3(new_n634), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n739), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n747), .A2(new_n699), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n747), .B2(new_n699), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n710), .B1(new_n732), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n728), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n719), .B1(new_n755), .B2(G1), .ZN(G364));
  NAND2_X1  g0556(.A1(new_n320), .A2(G200), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT96), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n759), .A2(new_n207), .A3(G190), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n759), .A2(new_n207), .A3(new_n308), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G283), .A2(new_n760), .B1(new_n761), .B2(G303), .ZN(new_n762));
  INV_X1    g0562(.A(G326), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n207), .A2(new_n308), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n320), .A2(new_n340), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT97), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n762), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n207), .A2(G190), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT33), .B(G317), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n320), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n764), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n771), .A2(new_n772), .B1(new_n775), .B2(G322), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n769), .A2(new_n773), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n287), .B1(new_n778), .B2(G311), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n769), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G329), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n780), .A2(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G294), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n776), .A2(new_n779), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n774), .A2(new_n201), .B1(new_n777), .B2(new_n219), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(KEYINPUT95), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n788), .A2(KEYINPUT95), .ZN(new_n790));
  INV_X1    g0590(.A(new_n760), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n789), .B(new_n790), .C1(new_n791), .C2(new_n334), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n761), .A2(G87), .ZN(new_n793));
  OAI21_X1  g0593(.A(KEYINPUT32), .B1(new_n781), .B2(new_n356), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n781), .A2(KEYINPUT32), .A3(new_n356), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G97), .B2(new_n785), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n287), .B1(new_n766), .B2(new_n217), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G68), .B2(new_n771), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n793), .A2(new_n794), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n768), .A2(new_n787), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n234), .B1(G20), .B2(new_n446), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n715), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n261), .A2(G20), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G45), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n803), .A2(G1), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n714), .A2(new_n541), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G355), .B1(new_n492), .B2(new_n714), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n233), .A2(G45), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n250), .B2(G45), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n384), .A2(new_n385), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n714), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n808), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G13), .A2(G33), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(G20), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n801), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n806), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n802), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n709), .B2(new_n817), .ZN(new_n821));
  INV_X1    g0621(.A(new_n806), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n711), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n709), .A2(new_n710), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  AND2_X1   g0626(.A1(new_n344), .A2(new_n345), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n343), .A2(new_n701), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n827), .A2(new_n343), .B1(new_n342), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n346), .A2(new_n701), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n727), .B(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(new_n754), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n754), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(new_n806), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n801), .A2(new_n815), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n806), .B1(new_n219), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  INV_X1    g0639(.A(new_n785), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n541), .B1(new_n781), .B2(new_n839), .C1(new_n840), .C2(new_n213), .ZN(new_n841));
  INV_X1    g0641(.A(G283), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n842), .A2(new_n770), .B1(new_n774), .B2(new_n579), .ZN(new_n843));
  INV_X1    g0643(.A(G303), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n766), .A2(new_n844), .B1(new_n777), .B2(new_n492), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n841), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n760), .A2(G87), .ZN(new_n847));
  INV_X1    g0647(.A(new_n761), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n846), .B(new_n847), .C1(new_n334), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n760), .A2(G68), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n848), .B2(new_n217), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT98), .Z(new_n852));
  NOR2_X1   g0652(.A1(new_n770), .A2(new_n271), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n766), .A2(new_n854), .B1(new_n777), .B2(new_n356), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(G143), .C2(new_n775), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n856), .A2(KEYINPUT34), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(KEYINPUT34), .ZN(new_n858));
  INV_X1    g0658(.A(new_n811), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n840), .A2(new_n201), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n859), .B(new_n860), .C1(G132), .C2(new_n782), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n857), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n849), .B1(new_n852), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT99), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n801), .B1(new_n863), .B2(new_n864), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n838), .B1(new_n865), .B2(new_n866), .C1(new_n832), .C2(new_n816), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n836), .A2(new_n867), .ZN(G384));
  OAI211_X1 g0668(.A(G116), .B(new_n235), .C1(new_n528), .C2(KEYINPUT35), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(KEYINPUT35), .B2(new_n528), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT36), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n232), .A2(new_n219), .A3(new_n359), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n872), .A2(KEYINPUT100), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n872), .A2(KEYINPUT100), .B1(new_n217), .B2(G68), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n206), .B(G13), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n877));
  AND3_X1   g0677(.A1(new_n409), .A2(new_n351), .A3(new_n418), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n410), .ZN(new_n879));
  INV_X1    g0679(.A(new_n697), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n391), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n413), .A2(new_n881), .A3(new_n884), .A4(new_n419), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n881), .B1(new_n420), .B2(new_n663), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n877), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n351), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n372), .A2(new_n256), .A3(new_n373), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n892), .B1(new_n893), .B2(new_n406), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n260), .B1(new_n388), .B2(new_n389), .ZN(new_n895));
  INV_X1    g0695(.A(new_n352), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n404), .B2(new_n405), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n351), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n894), .A2(new_n418), .B1(new_n898), .B2(new_n880), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n399), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n884), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT101), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n879), .A2(new_n902), .A3(new_n884), .A4(new_n881), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n898), .A2(new_n880), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n416), .B2(new_n420), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT104), .B1(new_n891), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n458), .A2(new_n699), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n459), .A2(new_n461), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n461), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n458), .B(new_n699), .C1(new_n449), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n747), .A2(new_n699), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n748), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n732), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT31), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n832), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n916), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n901), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n886), .B2(new_n887), .ZN(new_n926));
  INV_X1    g0726(.A(new_n906), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n421), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n926), .A2(KEYINPUT38), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n877), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n903), .A2(new_n904), .B1(new_n882), .B2(KEYINPUT37), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(new_n931), .B2(new_n889), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT104), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n929), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n910), .A2(KEYINPUT40), .A3(new_n924), .A4(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT103), .B1(new_n916), .B2(new_n923), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT103), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n732), .A2(new_n919), .B1(new_n921), .B2(new_n918), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n915), .A2(new_n937), .A3(new_n832), .A4(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n908), .B1(new_n905), .B2(new_n907), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n936), .A2(new_n939), .B1(new_n929), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n935), .B1(new_n941), .B2(KEYINPUT40), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n669), .A2(new_n938), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n942), .B(new_n943), .Z(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n710), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n459), .A2(new_n699), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n929), .A2(new_n932), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n947), .B1(new_n929), .B2(new_n940), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n688), .A2(new_n689), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n608), .B1(new_n652), .B2(new_n653), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n678), .B1(new_n704), .B2(new_n952), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n590), .A2(new_n611), .A3(new_n608), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n611), .B1(new_n590), .B2(new_n608), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n685), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n720), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n951), .B1(new_n958), .B2(new_n721), .ZN(new_n959));
  INV_X1    g0759(.A(new_n672), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n701), .B(new_n832), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n830), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT38), .B1(new_n926), .B2(new_n928), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n962), .B(new_n915), .C1(new_n909), .C2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n663), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n697), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n950), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n667), .B1(new_n728), .B2(new_n464), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n967), .B(new_n968), .Z(new_n969));
  OAI22_X1  g0769(.A1(new_n945), .A2(new_n969), .B1(new_n206), .B2(new_n804), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n945), .A2(new_n969), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n876), .B1(new_n970), .B2(new_n971), .ZN(G367));
  NAND2_X1  g0772(.A1(new_n475), .A2(new_n503), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n699), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n677), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n960), .B2(new_n974), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT43), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n978), .B1(new_n979), .B2(new_n976), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n703), .A2(new_n705), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n576), .B1(new_n565), .B2(new_n701), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n687), .A2(new_n699), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  OR3_X1    g0785(.A1(new_n981), .A2(new_n985), .A3(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT42), .B1(new_n981), .B2(new_n985), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n660), .B1(new_n565), .B2(new_n575), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n701), .B1(new_n988), .B2(new_n687), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  MUX2_X1   g0790(.A(new_n978), .B(new_n980), .S(new_n990), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n712), .A2(new_n985), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT106), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(KEYINPUT106), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n991), .A2(new_n992), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n715), .B(KEYINPUT41), .Z(new_n998));
  NAND2_X1  g0798(.A1(new_n706), .A2(new_n984), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT45), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n706), .A2(new_n984), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT107), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(KEYINPUT44), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(KEYINPUT44), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT108), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1000), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n712), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1008), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n703), .B(new_n705), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(new_n711), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n755), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1011), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n998), .B1(new_n1017), .B2(new_n755), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n805), .A2(G1), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n994), .B(new_n997), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n976), .A2(new_n817), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n812), .A2(new_n246), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n818), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n714), .B2(new_n479), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n806), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G294), .A2(new_n771), .B1(new_n782), .B2(G317), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n842), .B2(new_n777), .C1(new_n844), .C2(new_n774), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n811), .B(new_n1027), .C1(G107), .C2(new_n785), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n767), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1029), .A2(G311), .B1(G97), .B2(new_n760), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT46), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n848), .B2(new_n492), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n761), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n287), .B1(new_n774), .B2(new_n271), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n840), .A2(new_n202), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n760), .C2(G77), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1029), .A2(G143), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n770), .A2(new_n356), .B1(new_n777), .B2(new_n217), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT109), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n761), .A2(G58), .B1(G137), .B2(new_n782), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT110), .Z(new_n1043));
  OAI21_X1  g0843(.A(new_n1034), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT47), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n801), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1021), .B(new_n1025), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1020), .A2(new_n1048), .ZN(G387));
  NAND2_X1  g0849(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT111), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n807), .A2(new_n716), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(G107), .B2(new_n227), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n243), .A2(G45), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n326), .A2(new_n217), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT50), .Z(new_n1056));
  AOI211_X1 g0856(.A(G45), .B(new_n716), .C1(G68), .C2(G77), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n813), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1053), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n822), .B1(new_n1059), .B2(new_n1023), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n848), .A2(new_n579), .B1(new_n840), .B2(new_n842), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G317), .A2(new_n775), .B1(new_n778), .B2(G303), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n839), .B2(new_n770), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G322), .B2(new_n1029), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1061), .B1(new_n1064), .B2(KEYINPUT48), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT112), .Z(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(KEYINPUT48), .B2(new_n1064), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT49), .Z(new_n1068));
  OAI221_X1 g0868(.A(new_n859), .B1(new_n763), .B2(new_n781), .C1(new_n791), .C2(new_n492), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n479), .A2(new_n785), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n811), .C1(new_n277), .C2(new_n770), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n760), .A2(G97), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n761), .A2(G77), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G68), .A2(new_n778), .B1(new_n782), .B2(G150), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n766), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G159), .A2(new_n1075), .B1(new_n775), .B2(G50), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1068), .A2(new_n1069), .B1(new_n1071), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1060), .B1(new_n1078), .B2(new_n801), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n817), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n703), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n755), .A2(new_n1014), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1015), .A2(new_n715), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1051), .B(new_n1081), .C1(new_n1082), .C2(new_n1083), .ZN(G393));
  INV_X1    g0884(.A(KEYINPUT113), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1010), .B1(new_n1085), .B2(new_n1012), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1012), .A2(new_n1085), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n1087), .A3(new_n1019), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n818), .B1(new_n213), .B2(new_n227), .C1(new_n813), .C2(new_n253), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n822), .ZN(new_n1090));
  INV_X1    g0890(.A(G317), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n766), .A2(new_n1091), .B1(new_n774), .B2(new_n839), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT52), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n760), .A2(G107), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n1093), .B2(new_n1092), .C1(new_n842), .C2(new_n848), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G303), .A2(new_n771), .B1(new_n782), .B2(G322), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n287), .B1(new_n778), .B2(G294), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n492), .C2(new_n840), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n766), .A2(new_n271), .B1(new_n774), .B2(new_n356), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n847), .C1(new_n202), .C2(new_n848), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G50), .A2(new_n771), .B1(new_n778), .B2(new_n326), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n782), .A2(G143), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n785), .A2(G77), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1102), .A2(new_n811), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1095), .A2(new_n1098), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1090), .B1(new_n1106), .B2(new_n801), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n984), .B2(new_n1080), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1016), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1017), .A2(new_n715), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1088), .B(new_n1108), .C1(new_n1109), .C2(new_n1110), .ZN(G390));
  OAI211_X1 g0911(.A(new_n701), .B(new_n829), .C1(new_n723), .C2(new_n725), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n830), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n946), .B1(new_n1113), .B2(new_n915), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n910), .A2(new_n1114), .A3(new_n934), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n946), .B1(new_n962), .B2(new_n915), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT39), .B1(new_n963), .B2(new_n909), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n929), .A2(new_n932), .A3(new_n947), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1115), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n915), .A2(G330), .A3(new_n832), .A4(new_n938), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n710), .B(new_n831), .C1(new_n732), .C2(new_n752), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n915), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1115), .B(new_n1125), .C1(new_n1116), .C2(new_n1119), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n422), .A2(new_n463), .A3(G330), .A4(new_n938), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1127), .B(new_n667), .C1(new_n728), .C2(new_n464), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT114), .B1(new_n1124), .B2(new_n915), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n661), .A2(new_n515), .A3(new_n699), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n917), .A2(new_n921), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n917), .B2(new_n748), .ZN(new_n1132));
  OAI211_X1 g0932(.A(G330), .B(new_n832), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT114), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n912), .A4(new_n914), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1135), .A3(new_n1121), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n962), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n916), .B1(new_n923), .B2(new_n710), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1138), .A2(new_n830), .A3(new_n1112), .A4(new_n1125), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1128), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1123), .A2(new_n1126), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n715), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT115), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT115), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1141), .A2(new_n1144), .A3(new_n715), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT116), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1140), .B(new_n1146), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1143), .B(new_n1145), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n761), .A2(G150), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT53), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n760), .A2(G50), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n287), .B1(new_n770), .B2(new_n854), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G159), .B2(new_n785), .ZN(new_n1154));
  XOR2_X1   g0954(.A(KEYINPUT54), .B(G143), .Z(new_n1155));
  AOI22_X1  g0955(.A1(G132), .A2(new_n775), .B1(new_n778), .B2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1075), .A2(G128), .B1(new_n782), .B2(G125), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1152), .A2(new_n1154), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n770), .A2(new_n334), .B1(new_n777), .B2(new_n213), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT117), .Z(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n793), .A3(new_n850), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1075), .A2(G283), .B1(new_n782), .B2(G294), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n287), .B1(new_n775), .B2(G116), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1104), .A3(new_n1163), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n1151), .A2(new_n1158), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n801), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n806), .B1(new_n277), .B2(new_n837), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n1119), .C2(new_n816), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1148), .B2(new_n1019), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1149), .A2(new_n1170), .ZN(G378));
  OAI211_X1 g0971(.A(G330), .B(new_n935), .C1(new_n941), .C2(KEYINPUT40), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n318), .A2(new_n322), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1175));
  XNOR2_X1  g0975(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n281), .A2(new_n880), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT120), .Z(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1176), .B(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1119), .A2(new_n946), .B1(new_n965), .B2(new_n697), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n964), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n950), .A2(new_n964), .A3(new_n1180), .A4(new_n966), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1173), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1180), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n967), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(new_n1172), .A3(new_n1183), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1019), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n806), .B1(new_n217), .B2(new_n837), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n760), .A2(G58), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n774), .A2(new_n334), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT118), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n811), .A2(G41), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1073), .A2(new_n1192), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n766), .A2(new_n492), .B1(new_n781), .B2(new_n842), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n770), .A2(new_n213), .B1(new_n777), .B2(new_n329), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(new_n1196), .A2(new_n1036), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n761), .A2(new_n1155), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G125), .A2(new_n1075), .B1(new_n775), .B2(G128), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n785), .A2(G150), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G132), .A2(new_n771), .B1(new_n778), .B2(G137), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n760), .A2(G159), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G33), .B(G41), .C1(new_n782), .C2(G124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G50), .B(new_n1195), .C1(new_n272), .C2(new_n551), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1200), .A2(new_n1201), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(KEYINPUT119), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT119), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n801), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1191), .B1(new_n1215), .B2(new_n1217), .C1(new_n1186), .C2(new_n816), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1190), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1128), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1141), .A2(new_n1221), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1187), .A2(new_n1172), .A3(new_n1183), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1172), .B1(new_n1187), .B2(new_n1183), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT57), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT121), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1189), .A2(new_n1228), .A3(KEYINPUT57), .A4(new_n1222), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n715), .A3(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1185), .A2(new_n1188), .B1(new_n1221), .B2(new_n1141), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1228), .B1(new_n1231), .B2(KEYINPUT57), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1220), .B1(new_n1230), .B2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n916), .A2(new_n815), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1075), .A2(G294), .B1(new_n778), .B2(G107), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G283), .A2(new_n775), .B1(new_n782), .B2(G303), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n287), .B1(new_n771), .B2(G116), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1070), .A4(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n219), .A2(new_n791), .B1(new_n848), .B2(new_n213), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n761), .A2(G159), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1075), .A2(G132), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G137), .A2(new_n775), .B1(new_n778), .B2(G150), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1192), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n771), .A2(new_n1155), .B1(new_n782), .B2(G128), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1245), .B(new_n811), .C1(new_n217), .C2(new_n840), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1239), .A2(new_n1240), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1247), .A2(new_n801), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n806), .B(new_n1248), .C1(new_n202), .C2(new_n837), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1234), .A2(new_n1019), .B1(new_n1235), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1137), .A2(new_n1128), .A3(new_n1139), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n998), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1250), .B1(new_n1147), .B2(new_n1253), .ZN(G381));
  OR2_X1    g1054(.A1(G375), .A2(G378), .ZN(new_n1255));
  OR2_X1    g1055(.A1(G387), .A2(G390), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT122), .ZN(new_n1258));
  OR4_X1    g1058(.A1(G381), .A2(new_n1255), .A3(new_n1256), .A4(new_n1258), .ZN(G407));
  OAI211_X1 g1059(.A(G407), .B(G213), .C1(G343), .C2(new_n1255), .ZN(G409));
  XNOR2_X1  g1060(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n698), .A2(G213), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G378), .B(new_n1220), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1225), .A2(new_n998), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1149), .B(new_n1170), .C1(new_n1219), .C2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT123), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1265), .A2(KEYINPUT123), .A3(new_n1267), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1264), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1251), .B(KEYINPUT60), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1140), .A2(new_n803), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT124), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1273), .A2(KEYINPUT124), .A3(new_n1274), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1250), .A3(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(G384), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1262), .B1(new_n1272), .B2(new_n1280), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1265), .A2(KEYINPUT123), .A3(new_n1267), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT123), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1263), .B(new_n1280), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(KEYINPUT125), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1261), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G387), .A2(G390), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(new_n825), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1256), .B(new_n1287), .C1(KEYINPUT127), .C2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(KEYINPUT127), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1289), .B(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1264), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(KEYINPUT63), .A3(new_n1280), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1291), .A2(new_n1292), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1264), .A2(G2897), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1280), .B(new_n1296), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1272), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1286), .A2(new_n1295), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1292), .B1(new_n1297), .B2(new_n1293), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1293), .A2(KEYINPUT62), .A3(new_n1280), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1300), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1299), .B1(new_n1304), .B2(new_n1291), .ZN(G405));
  OR2_X1    g1105(.A1(new_n1291), .A2(new_n1280), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1291), .A2(new_n1280), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  XOR2_X1   g1108(.A(G375), .B(G378), .Z(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1306), .A2(new_n1309), .A3(new_n1307), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(G402));
endmodule


