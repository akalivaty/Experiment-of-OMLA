

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590;

  XOR2_X1 U328 ( .A(n418), .B(n417), .Z(n527) );
  XNOR2_X1 U329 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U330 ( .A(n399), .B(n398), .ZN(n523) );
  AND2_X1 U331 ( .A1(n448), .A2(n447), .ZN(n296) );
  XOR2_X1 U332 ( .A(n389), .B(n388), .Z(n297) );
  XNOR2_X1 U333 ( .A(n423), .B(KEYINPUT96), .ZN(n424) );
  XNOR2_X1 U334 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n464) );
  XNOR2_X1 U335 ( .A(n465), .B(n464), .ZN(n467) );
  INV_X1 U336 ( .A(n449), .ZN(n447) );
  XNOR2_X1 U337 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U338 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U339 ( .A(n390), .B(n297), .ZN(n394) );
  XNOR2_X1 U340 ( .A(n566), .B(n363), .ZN(n588) );
  XNOR2_X1 U341 ( .A(KEYINPUT121), .B(n479), .ZN(n568) );
  XNOR2_X1 U342 ( .A(n362), .B(n361), .ZN(n566) );
  INV_X1 U343 ( .A(G106GAT), .ZN(n456) );
  XOR2_X1 U344 ( .A(KEYINPUT90), .B(n449), .Z(n571) );
  XNOR2_X1 U345 ( .A(G183GAT), .B(KEYINPUT124), .ZN(n480) );
  XNOR2_X1 U346 ( .A(n456), .B(KEYINPUT44), .ZN(n457) );
  XNOR2_X1 U347 ( .A(n481), .B(n480), .ZN(G1350GAT) );
  XOR2_X1 U348 ( .A(G148GAT), .B(KEYINPUT85), .Z(n301) );
  XOR2_X1 U349 ( .A(G50GAT), .B(G218GAT), .Z(n348) );
  XOR2_X1 U350 ( .A(G211GAT), .B(KEYINPUT21), .Z(n299) );
  XNOR2_X1 U351 ( .A(G197GAT), .B(KEYINPUT84), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n392) );
  XNOR2_X1 U353 ( .A(n348), .B(n392), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n306) );
  XNOR2_X1 U355 ( .A(G106GAT), .B(G78GAT), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n302), .B(G204GAT), .ZN(n335) );
  XOR2_X1 U357 ( .A(n335), .B(KEYINPUT83), .Z(n304) );
  NAND2_X1 U358 ( .A1(G228GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U360 ( .A(n306), .B(n305), .Z(n314) );
  XOR2_X1 U361 ( .A(KEYINPUT2), .B(G162GAT), .Z(n308) );
  XNOR2_X1 U362 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U364 ( .A(G141GAT), .B(n309), .Z(n444) );
  XOR2_X1 U365 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n311) );
  XNOR2_X1 U366 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n444), .B(n312), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n314), .B(n313), .ZN(n474) );
  XOR2_X1 U370 ( .A(n474), .B(KEYINPUT28), .Z(n518) );
  XOR2_X1 U371 ( .A(KEYINPUT69), .B(G141GAT), .Z(n316) );
  XNOR2_X1 U372 ( .A(G50GAT), .B(G197GAT), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U374 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n318) );
  XNOR2_X1 U375 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n330) );
  XNOR2_X1 U378 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n321), .B(KEYINPUT7), .ZN(n347) );
  XOR2_X1 U380 ( .A(n347), .B(KEYINPUT70), .Z(n323) );
  NAND2_X1 U381 ( .A1(G229GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U383 ( .A(G169GAT), .B(G8GAT), .Z(n387) );
  XNOR2_X1 U384 ( .A(n324), .B(n387), .ZN(n328) );
  XOR2_X1 U385 ( .A(G36GAT), .B(G29GAT), .Z(n326) );
  XOR2_X1 U386 ( .A(G22GAT), .B(G15GAT), .Z(n367) );
  XOR2_X1 U387 ( .A(G113GAT), .B(G1GAT), .Z(n434) );
  XNOR2_X1 U388 ( .A(n367), .B(n434), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n576) );
  INV_X1 U392 ( .A(n576), .ZN(n549) );
  XNOR2_X1 U393 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n331), .B(KEYINPUT13), .ZN(n370) );
  XOR2_X1 U395 ( .A(KEYINPUT73), .B(G92GAT), .Z(n333) );
  XNOR2_X1 U396 ( .A(G99GAT), .B(G85GAT), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n346) );
  XOR2_X1 U398 ( .A(n370), .B(n346), .Z(n337) );
  XNOR2_X1 U399 ( .A(G120GAT), .B(G148GAT), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n334), .B(G57GAT), .ZN(n432) );
  XNOR2_X1 U401 ( .A(n335), .B(n432), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n344) );
  XOR2_X1 U403 ( .A(G176GAT), .B(G64GAT), .Z(n389) );
  XOR2_X1 U404 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n339) );
  XNOR2_X1 U405 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n338) );
  XNOR2_X1 U406 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U407 ( .A(n389), .B(n340), .Z(n342) );
  NAND2_X1 U408 ( .A1(G230GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U410 ( .A(n344), .B(n343), .Z(n581) );
  XOR2_X1 U411 ( .A(n581), .B(KEYINPUT41), .Z(n563) );
  NAND2_X1 U412 ( .A1(n549), .A2(n563), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n345), .B(KEYINPUT105), .ZN(n509) );
  XNOR2_X1 U414 ( .A(n347), .B(n346), .ZN(n362) );
  XOR2_X1 U415 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n350) );
  XOR2_X1 U416 ( .A(G36GAT), .B(G190GAT), .Z(n391) );
  XNOR2_X1 U417 ( .A(n348), .B(n391), .ZN(n349) );
  XNOR2_X1 U418 ( .A(n350), .B(n349), .ZN(n356) );
  XOR2_X1 U419 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n352) );
  XNOR2_X1 U420 ( .A(G162GAT), .B(G106GAT), .ZN(n351) );
  XNOR2_X1 U421 ( .A(n352), .B(n351), .ZN(n354) );
  AND2_X1 U422 ( .A1(G232GAT), .A2(G233GAT), .ZN(n353) );
  XOR2_X1 U423 ( .A(n357), .B(KEYINPUT64), .Z(n360) );
  XNOR2_X1 U424 ( .A(G29GAT), .B(G134GAT), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n358), .B(KEYINPUT75), .ZN(n428) );
  XNOR2_X1 U426 ( .A(n428), .B(KEYINPUT74), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U428 ( .A(KEYINPUT36), .B(KEYINPUT102), .Z(n363) );
  XOR2_X1 U429 ( .A(G211GAT), .B(G78GAT), .Z(n365) );
  XNOR2_X1 U430 ( .A(G127GAT), .B(G155GAT), .ZN(n364) );
  XNOR2_X1 U431 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U432 ( .A(n366), .B(G64GAT), .Z(n369) );
  XNOR2_X1 U433 ( .A(n367), .B(G183GAT), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n374) );
  XOR2_X1 U435 ( .A(n370), .B(G57GAT), .Z(n372) );
  NAND2_X1 U436 ( .A1(G231GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U438 ( .A(n374), .B(n373), .Z(n382) );
  XOR2_X1 U439 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n376) );
  XNOR2_X1 U440 ( .A(G8GAT), .B(KEYINPUT78), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U442 ( .A(KEYINPUT12), .B(KEYINPUT77), .Z(n378) );
  XNOR2_X1 U443 ( .A(G1GAT), .B(KEYINPUT76), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n584) );
  XOR2_X1 U447 ( .A(G183GAT), .B(KEYINPUT18), .Z(n384) );
  XNOR2_X1 U448 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n384), .B(n383), .ZN(n386) );
  XNOR2_X1 U450 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n416) );
  XNOR2_X1 U452 ( .A(n387), .B(n416), .ZN(n390) );
  XOR2_X1 U453 ( .A(G92GAT), .B(G218GAT), .Z(n388) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U456 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n396) );
  NAND2_X1 U457 ( .A1(G226GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U459 ( .A(G204GAT), .B(n397), .Z(n398) );
  XOR2_X1 U460 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n400) );
  XNOR2_X1 U461 ( .A(n523), .B(n400), .ZN(n450) );
  XOR2_X1 U462 ( .A(KEYINPUT65), .B(G176GAT), .Z(n402) );
  XNOR2_X1 U463 ( .A(G169GAT), .B(G120GAT), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n415) );
  XOR2_X1 U465 ( .A(G99GAT), .B(G190GAT), .Z(n404) );
  XNOR2_X1 U466 ( .A(G43GAT), .B(G134GAT), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U468 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n406) );
  XNOR2_X1 U469 ( .A(G113GAT), .B(G71GAT), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U471 ( .A(n408), .B(n407), .Z(n413) );
  XOR2_X1 U472 ( .A(KEYINPUT0), .B(G127GAT), .Z(n433) );
  XOR2_X1 U473 ( .A(n433), .B(KEYINPUT79), .Z(n410) );
  NAND2_X1 U474 ( .A1(G227GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U476 ( .A(G15GAT), .B(n411), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n418) );
  INV_X1 U479 ( .A(n416), .ZN(n417) );
  NAND2_X1 U480 ( .A1(n474), .A2(n527), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n419), .B(KEYINPUT94), .ZN(n420) );
  XNOR2_X1 U482 ( .A(KEYINPUT26), .B(n420), .ZN(n573) );
  NOR2_X1 U483 ( .A1(n450), .A2(n573), .ZN(n548) );
  NOR2_X1 U484 ( .A1(n527), .A2(n523), .ZN(n421) );
  XOR2_X1 U485 ( .A(KEYINPUT95), .B(n421), .Z(n422) );
  NOR2_X1 U486 ( .A1(n474), .A2(n422), .ZN(n425) );
  INV_X1 U487 ( .A(KEYINPUT25), .ZN(n423) );
  NOR2_X1 U488 ( .A1(n548), .A2(n426), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n427), .B(KEYINPUT97), .ZN(n448) );
  XOR2_X1 U490 ( .A(KEYINPUT89), .B(n428), .Z(n430) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U493 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U496 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n438) );
  XNOR2_X1 U497 ( .A(G85GAT), .B(KEYINPUT6), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n446) );
  XOR2_X1 U500 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n442) );
  XNOR2_X1 U501 ( .A(KEYINPUT86), .B(KEYINPUT4), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n449) );
  NOR2_X1 U505 ( .A1(n571), .A2(n450), .ZN(n451) );
  NAND2_X1 U506 ( .A1(n451), .A2(n518), .ZN(n529) );
  INV_X1 U507 ( .A(n527), .ZN(n530) );
  NOR2_X1 U508 ( .A1(n529), .A2(n530), .ZN(n452) );
  NOR2_X1 U509 ( .A1(n296), .A2(n452), .ZN(n484) );
  NOR2_X1 U510 ( .A1(n584), .A2(n484), .ZN(n453) );
  NAND2_X1 U511 ( .A1(n588), .A2(n453), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT37), .ZN(n497) );
  NAND2_X1 U513 ( .A1(n509), .A2(n497), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n455), .B(KEYINPUT110), .ZN(n526) );
  NOR2_X1 U515 ( .A1(n518), .A2(n526), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(G1339GAT) );
  XNOR2_X1 U517 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n477) );
  INV_X1 U518 ( .A(n563), .ZN(n551) );
  NOR2_X1 U519 ( .A1(n549), .A2(n551), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n459), .B(KEYINPUT46), .ZN(n460) );
  NOR2_X1 U521 ( .A1(n584), .A2(n460), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n461), .A2(n566), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n462), .B(KEYINPUT47), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT112), .ZN(n470) );
  NAND2_X1 U525 ( .A1(n588), .A2(n584), .ZN(n465) );
  INV_X1 U526 ( .A(n581), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n468), .A2(n576), .ZN(n469) );
  NOR2_X1 U529 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U530 ( .A(KEYINPUT48), .B(n471), .ZN(n546) );
  NOR2_X1 U531 ( .A1(n546), .A2(n523), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT54), .ZN(n572) );
  INV_X1 U533 ( .A(n571), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n475) );
  AND2_X1 U535 ( .A1(n572), .A2(n475), .ZN(n476) );
  XOR2_X1 U536 ( .A(n477), .B(n476), .Z(n478) );
  NAND2_X1 U537 ( .A1(n530), .A2(n478), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n568), .A2(n584), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n581), .A2(n549), .ZN(n498) );
  NAND2_X1 U540 ( .A1(n566), .A2(n584), .ZN(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT16), .B(n482), .ZN(n483) );
  NOR2_X1 U542 ( .A1(n484), .A2(n483), .ZN(n508) );
  NAND2_X1 U543 ( .A1(n498), .A2(n508), .ZN(n493) );
  NOR2_X1 U544 ( .A1(n571), .A2(n493), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U547 ( .A(G1GAT), .B(n487), .Z(G1324GAT) );
  NOR2_X1 U548 ( .A1(n523), .A2(n493), .ZN(n488) );
  XOR2_X1 U549 ( .A(G8GAT), .B(n488), .Z(G1325GAT) );
  NOR2_X1 U550 ( .A1(n493), .A2(n527), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n490) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  NOR2_X1 U555 ( .A1(n518), .A2(n493), .ZN(n494) );
  XOR2_X1 U556 ( .A(G22GAT), .B(n494), .Z(G1327GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n496) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n501) );
  NAND2_X1 U560 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(KEYINPUT38), .ZN(n506) );
  NOR2_X1 U562 ( .A1(n571), .A2(n506), .ZN(n500) );
  XOR2_X1 U563 ( .A(n501), .B(n500), .Z(G1328GAT) );
  NOR2_X1 U564 ( .A1(n506), .A2(n523), .ZN(n502) );
  XOR2_X1 U565 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  XNOR2_X1 U566 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n504) );
  NOR2_X1 U567 ( .A1(n527), .A2(n506), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U569 ( .A(G43GAT), .B(n505), .Z(G1330GAT) );
  NOR2_X1 U570 ( .A1(n518), .A2(n506), .ZN(n507) );
  XOR2_X1 U571 ( .A(G50GAT), .B(n507), .Z(G1331GAT) );
  NAND2_X1 U572 ( .A1(n509), .A2(n508), .ZN(n517) );
  NOR2_X1 U573 ( .A1(n571), .A2(n517), .ZN(n511) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U576 ( .A(G57GAT), .B(n512), .Z(G1332GAT) );
  NOR2_X1 U577 ( .A1(n523), .A2(n517), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1333GAT) );
  NOR2_X1 U580 ( .A1(n527), .A2(n517), .ZN(n515) );
  XOR2_X1 U581 ( .A(KEYINPUT108), .B(n515), .Z(n516) );
  XNOR2_X1 U582 ( .A(G71GAT), .B(n516), .ZN(G1334GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n520) );
  XNOR2_X1 U584 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U586 ( .A(G78GAT), .B(n521), .Z(G1335GAT) );
  NOR2_X1 U587 ( .A1(n571), .A2(n526), .ZN(n522) );
  XOR2_X1 U588 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U589 ( .A1(n526), .A2(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1337GAT) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n528), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n546), .A2(n529), .ZN(n531) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n542) );
  NOR2_X1 U596 ( .A1(n549), .A2(n542), .ZN(n532) );
  XOR2_X1 U597 ( .A(KEYINPUT114), .B(n532), .Z(n533) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  NOR2_X1 U599 ( .A1(n542), .A2(n551), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n535) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT116), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n539) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n541) );
  INV_X1 U607 ( .A(n584), .ZN(n555) );
  NOR2_X1 U608 ( .A1(n555), .A2(n542), .ZN(n540) );
  XOR2_X1 U609 ( .A(n541), .B(n540), .Z(G1342GAT) );
  NOR2_X1 U610 ( .A1(n566), .A2(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U613 ( .A(G134GAT), .B(n545), .Z(G1343GAT) );
  NOR2_X1 U614 ( .A1(n571), .A2(n546), .ZN(n547) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n557) );
  NOR2_X1 U616 ( .A1(n549), .A2(n557), .ZN(n550) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n550), .Z(G1344GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n557), .ZN(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n557), .ZN(n556) );
  XOR2_X1 U623 ( .A(G155GAT), .B(n556), .Z(G1346GAT) );
  NOR2_X1 U624 ( .A1(n566), .A2(n557), .ZN(n558) );
  XOR2_X1 U625 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  NAND2_X1 U626 ( .A1(n576), .A2(n568), .ZN(n559) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n560) );
  XNOR2_X1 U630 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U631 ( .A(KEYINPUT122), .B(n562), .Z(n565) );
  NAND2_X1 U632 ( .A1(n568), .A2(n563), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  INV_X1 U635 ( .A(n566), .ZN(n567) );
  NAND2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1351GAT) );
  XNOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n580) );
  XOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT126), .Z(n578) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n574) );
  NOR2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(n575), .Z(n587) );
  NAND2_X1 U643 ( .A1(n587), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U647 ( .A1(n587), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  XOR2_X1 U649 ( .A(G211GAT), .B(KEYINPUT127), .Z(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  NAND2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n589), .B(KEYINPUT62), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

