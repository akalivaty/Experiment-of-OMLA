//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G77), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n234), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G68), .Z(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT68), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT68), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n251), .A2(new_n248), .A3(G13), .A4(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n210), .B1(new_n206), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n257), .B(KEYINPUT69), .Z(new_n258));
  NAND2_X1  g0058(.A1(new_n248), .A2(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  XOR2_X1   g0060(.A(new_n260), .B(KEYINPUT70), .Z(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n254), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n211), .A2(new_n254), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n264), .A2(new_n265), .B1(G150), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n203), .A2(G20), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n256), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n253), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n202), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT9), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G226), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n275), .A2(new_n280), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G222), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n287), .A2(new_n289), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G223), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n292), .B1(new_n220), .B2(new_n293), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n275), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n286), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G200), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n274), .B(new_n302), .C1(new_n303), .C2(new_n301), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT10), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n301), .A2(G179), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n273), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT15), .B(G87), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(new_n265), .B1(new_n219), .B2(G20), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n263), .B2(new_n266), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n255), .ZN(new_n315));
  INV_X1    g0115(.A(new_n257), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(G77), .A3(new_n259), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n271), .A2(new_n220), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n275), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n295), .A2(G238), .B1(G107), .B2(new_n290), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n291), .A2(G232), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n281), .B1(new_n284), .B2(new_n221), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT71), .ZN(new_n326));
  OAI211_X1 g0126(.A(KEYINPUT72), .B(new_n319), .C1(new_n326), .C2(G169), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n319), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT71), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n325), .B(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n333), .B2(new_n307), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(KEYINPUT72), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n319), .B1(new_n326), .B2(G190), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n326), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n281), .B1(new_n284), .B2(new_n218), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n291), .A2(G226), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G97), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n344), .C1(new_n296), .C2(new_n236), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n342), .B1(new_n345), .B2(new_n275), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n341), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n347), .B2(new_n346), .ZN(new_n349));
  OR3_X1    g0149(.A1(new_n346), .A2(KEYINPUT73), .A3(new_n347), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(G169), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT14), .ZN(new_n352));
  OR3_X1    g0152(.A1(new_n346), .A2(KEYINPUT74), .A3(new_n347), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n346), .A2(new_n347), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT74), .B1(new_n346), .B2(new_n347), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n353), .A2(G179), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n349), .A2(new_n357), .A3(G169), .A4(new_n350), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n316), .A2(G68), .A3(new_n259), .ZN(new_n360));
  XOR2_X1   g0160(.A(new_n360), .B(KEYINPUT75), .Z(new_n361));
  AOI22_X1  g0161(.A1(new_n265), .A2(G77), .B1(G20), .B2(new_n217), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n202), .B2(new_n266), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n255), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT11), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n271), .A2(new_n217), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT12), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n361), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n359), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n349), .A2(G200), .A3(new_n350), .ZN(new_n370));
  INV_X1    g0170(.A(new_n368), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n353), .A2(G190), .A3(new_n354), .A4(new_n355), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n310), .A2(new_n340), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n211), .A2(KEYINPUT7), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n254), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n254), .ZN(new_n384));
  NAND2_X1  g0184(.A1(KEYINPUT76), .A2(G33), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT3), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT79), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n385), .ZN(new_n389));
  NOR2_X1   g0189(.A1(KEYINPUT76), .A2(G33), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n387), .B(new_n288), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n378), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT7), .B1(new_n290), .B2(new_n211), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n217), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(G58), .B(G68), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(G20), .B1(new_n267), .B2(G159), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n376), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT80), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n384), .A2(KEYINPUT3), .A3(new_n385), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT77), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n288), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(G33), .A3(new_n379), .ZN(new_n406));
  AOI21_X1  g0206(.A(G20), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT7), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n217), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n403), .A2(new_n406), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT7), .B1(new_n410), .B2(G20), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n412), .B1(new_n409), .B2(new_n411), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT16), .B(new_n398), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n288), .B1(new_n389), .B2(new_n390), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT79), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n391), .A3(new_n382), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n394), .B1(new_n418), .B2(new_n378), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n398), .B1(new_n419), .B2(new_n217), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(KEYINPUT80), .A3(new_n376), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n402), .A2(new_n255), .A3(new_n415), .A4(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n263), .B1(new_n248), .B2(G20), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n258), .A2(new_n423), .B1(new_n271), .B2(new_n263), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n297), .A2(new_n294), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n410), .B(new_n425), .C1(G226), .C2(new_n294), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n320), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n281), .B1(new_n284), .B2(new_n236), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n303), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(G200), .B2(new_n430), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n422), .A2(new_n424), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(KEYINPUT17), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n422), .A2(new_n424), .A3(new_n432), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT83), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT83), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n422), .A2(new_n437), .A3(new_n432), .A4(new_n424), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n434), .B1(new_n439), .B2(KEYINPUT17), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n430), .A2(new_n307), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n428), .A2(new_n328), .A3(new_n429), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT82), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n422), .A2(new_n424), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n422), .A2(KEYINPUT81), .A3(new_n424), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT18), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n445), .A2(new_n448), .A3(new_n452), .A4(new_n449), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n375), .A2(new_n440), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT84), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT84), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n375), .A2(new_n457), .A3(new_n440), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G116), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n271), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n257), .B1(new_n248), .B2(G33), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(new_n461), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  INV_X1    g0266(.A(G97), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n466), .B(new_n211), .C1(G33), .C2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n255), .C1(new_n211), .C2(G116), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n469), .B(KEYINPUT20), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n307), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT5), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n277), .B1(new_n473), .B2(G41), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n248), .B(G45), .C1(new_n278), .C2(KEYINPUT5), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT85), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n473), .A2(G41), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n275), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(G270), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n403), .A2(new_n406), .A3(G264), .A4(G1698), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT87), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n403), .A2(new_n406), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1698), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n486), .A2(G257), .B1(G303), .B2(new_n290), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT88), .B1(new_n488), .B2(new_n275), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT88), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n490), .B(new_n320), .C1(new_n484), .C2(new_n487), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n481), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n472), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT21), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT21), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n472), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n489), .A2(new_n491), .ZN(new_n498));
  INV_X1    g0298(.A(new_n471), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n481), .A2(G179), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n499), .B1(new_n492), .B2(G200), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n303), .B2(new_n492), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n497), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n294), .A2(G257), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n410), .B(new_n505), .C1(G250), .C2(G1698), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n384), .A2(new_n385), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G294), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n320), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n480), .A2(G264), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR4_X1   g0311(.A1(new_n509), .A2(new_n477), .A3(new_n303), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(new_n508), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n513), .B2(new_n275), .ZN(new_n514));
  INV_X1    g0314(.A(new_n477), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n512), .B1(G200), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT22), .ZN(new_n518));
  INV_X1    g0318(.A(G87), .ZN(new_n519));
  NOR4_X1   g0319(.A1(new_n485), .A2(new_n518), .A3(G20), .A4(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n211), .A2(G87), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n518), .B1(new_n290), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n507), .A2(new_n211), .A3(G116), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n525));
  OR3_X1    g0325(.A1(new_n211), .A2(KEYINPUT23), .A3(G107), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n521), .A2(KEYINPUT89), .A3(new_n523), .A4(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT89), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n523), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(new_n520), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n531), .A3(KEYINPUT24), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n532), .B(new_n255), .C1(KEYINPUT24), .C2(new_n531), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT25), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n253), .B2(G107), .ZN(new_n535));
  INV_X1    g0335(.A(G107), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n271), .A2(KEYINPUT25), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n463), .A2(G107), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n517), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n514), .A2(new_n328), .A3(new_n515), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n509), .A2(new_n477), .A3(new_n511), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(G169), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n533), .B2(new_n538), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT90), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n221), .A2(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n410), .B(new_n545), .C1(G238), .C2(G1698), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n507), .A2(G116), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n320), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n279), .A2(G1), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n276), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n320), .B(new_n551), .C1(G250), .C2(new_n550), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT86), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n554), .A3(new_n328), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n410), .A2(new_n211), .A3(G68), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT19), .B1(new_n265), .B2(G97), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n211), .B1(new_n344), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n519), .A2(new_n467), .A3(new_n536), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n255), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n271), .A2(new_n311), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n564), .C1(new_n311), .C2(new_n464), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n307), .B1(new_n548), .B2(new_n553), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n555), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n549), .A2(new_n554), .A3(G190), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n463), .A2(G87), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n563), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(G200), .B1(new_n548), .B2(new_n553), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n393), .A2(new_n395), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G107), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n536), .A2(KEYINPUT6), .A3(G97), .ZN(new_n577));
  XOR2_X1   g0377(.A(G97), .B(G107), .Z(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(KEYINPUT6), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(G20), .B1(G77), .B2(new_n267), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n256), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n271), .A2(new_n467), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n464), .B2(new_n467), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n477), .B1(G257), .B2(new_n480), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n291), .A2(KEYINPUT4), .A3(G244), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n295), .A2(G250), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n466), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n486), .A2(G244), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n586), .B1(new_n592), .B2(new_n320), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n307), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n590), .ZN(new_n595));
  INV_X1    g0395(.A(new_n589), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n320), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n480), .A2(G257), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n515), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n328), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n585), .A2(new_n594), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n593), .A2(G200), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n584), .B(new_n603), .C1(new_n303), .C2(new_n593), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n574), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n533), .A2(new_n538), .ZN(new_n606));
  INV_X1    g0406(.A(new_n542), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT90), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n517), .A2(new_n533), .A3(new_n538), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n544), .A2(new_n605), .A3(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n460), .A2(new_n504), .A3(new_n612), .ZN(G372));
  INV_X1    g0413(.A(new_n309), .ZN(new_n614));
  INV_X1    g0414(.A(new_n336), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n373), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n369), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n440), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n443), .B1(new_n422), .B2(new_n424), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n619), .B(KEYINPUT18), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n614), .B1(new_n621), .B2(new_n305), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n497), .A2(new_n501), .A3(new_n608), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n610), .A2(new_n574), .A3(new_n602), .A4(new_n604), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n601), .A2(new_n594), .ZN(new_n626));
  XNOR2_X1  g0426(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n574), .A2(new_n585), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT26), .B1(new_n602), .B2(new_n573), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n567), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n622), .B1(new_n460), .B2(new_n631), .ZN(G369));
  NAND2_X1  g0432(.A1(new_n497), .A2(new_n501), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n248), .A2(new_n211), .A3(G13), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(G213), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(G343), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n471), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n504), .B2(new_n641), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G330), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n544), .A2(new_n611), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n606), .A2(new_n639), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n608), .B2(new_n640), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n639), .B1(new_n497), .B2(new_n501), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n543), .B2(new_n640), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n650), .A2(new_n653), .ZN(G399));
  INV_X1    g0454(.A(new_n207), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n560), .A2(G116), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G1), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n215), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT28), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n640), .B1(new_n625), .B2(new_n630), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT93), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT29), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT93), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n665), .B(new_n640), .C1(new_n625), .C2(new_n630), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n623), .A2(new_n624), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n574), .A2(new_n669), .A3(new_n626), .A4(new_n585), .ZN(new_n670));
  INV_X1    g0470(.A(new_n627), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n602), .B2(new_n573), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n670), .A2(new_n672), .A3(new_n567), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n639), .B1(new_n668), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT29), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G330), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n548), .A2(new_n553), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n500), .A2(new_n600), .A3(new_n514), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n498), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR4_X1   g0482(.A1(new_n600), .A2(new_n541), .A3(new_n678), .A4(G179), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n492), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT92), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(new_n686), .A3(new_n492), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n679), .A2(KEYINPUT30), .A3(new_n498), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n682), .A2(new_n685), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n639), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n612), .A2(new_n504), .A3(new_n639), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n682), .A2(new_n688), .ZN(new_n694));
  AOI211_X1 g0494(.A(new_n692), .B(new_n640), .C1(new_n694), .C2(new_n684), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n677), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n676), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n661), .B1(new_n698), .B2(G1), .ZN(G364));
  INV_X1    g0499(.A(G13), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G20), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n248), .B1(new_n701), .B2(G45), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n656), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n645), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(G330), .B2(new_n643), .ZN(new_n706));
  INV_X1    g0506(.A(new_n704), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n293), .A2(G355), .A3(new_n207), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n410), .A2(new_n655), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(G45), .B2(new_n215), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n246), .A2(new_n279), .ZN(new_n711));
  OAI221_X1 g0511(.A(new_n708), .B1(G116), .B2(new_n207), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G13), .A2(G33), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n210), .B1(G20), .B2(new_n307), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n707), .B1(new_n712), .B2(new_n717), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT94), .Z(new_n719));
  INV_X1    g0519(.A(new_n716), .ZN(new_n720));
  NAND2_X1  g0520(.A1(G20), .A2(G179), .ZN(new_n721));
  XOR2_X1   g0521(.A(new_n721), .B(KEYINPUT95), .Z(new_n722));
  NOR2_X1   g0522(.A1(new_n303), .A2(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G322), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n303), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n338), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(KEYINPUT33), .B(G317), .Z(new_n730));
  OAI21_X1  g0530(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT98), .Z(new_n732));
  NOR2_X1   g0532(.A1(new_n303), .A2(new_n338), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n211), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n293), .B1(new_n736), .B2(G303), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n303), .A3(new_n338), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G329), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n734), .A2(new_n303), .A3(G200), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n737), .B(new_n740), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n727), .A2(G200), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G311), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT97), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n722), .A2(new_n733), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n723), .A2(new_n328), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n750), .A2(G326), .B1(G294), .B2(new_n752), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n743), .B(new_n747), .C1(new_n748), .C2(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n732), .B(new_n754), .C1(new_n748), .C2(new_n753), .ZN(new_n755));
  INV_X1    g0555(.A(G159), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT32), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n752), .A2(G97), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n759), .B(new_n760), .C1(new_n729), .C2(new_n217), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n219), .B2(new_n744), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n742), .A2(new_n536), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n290), .B(new_n763), .C1(G87), .C2(new_n736), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT96), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n749), .A2(new_n202), .B1(new_n757), .B2(new_n758), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G58), .B2(new_n725), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n762), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n755), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n715), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n719), .B1(new_n720), .B2(new_n769), .C1(new_n643), .C2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n706), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(G396));
  NOR2_X1   g0573(.A1(new_n331), .A2(new_n640), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n339), .B(new_n775), .C1(new_n330), .C2(new_n335), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n336), .B2(new_n775), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n663), .A2(new_n666), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n662), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n777), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n697), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n704), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G137), .A2(new_n750), .B1(new_n725), .B2(G143), .ZN(new_n786));
  INV_X1    g0586(.A(G150), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n786), .B1(new_n745), .B2(new_n756), .C1(new_n787), .C2(new_n729), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT34), .Z(new_n789));
  OAI21_X1  g0589(.A(new_n410), .B1(new_n202), .B2(new_n735), .ZN(new_n790));
  INV_X1    g0590(.A(new_n742), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(G68), .B1(new_n739), .B2(G132), .ZN(new_n792));
  INV_X1    g0592(.A(G58), .ZN(new_n793));
  INV_X1    g0593(.A(new_n752), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n789), .A2(new_n790), .A3(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n461), .A2(new_n745), .B1(new_n729), .B2(new_n741), .ZN(new_n797));
  INV_X1    g0597(.A(G294), .ZN(new_n798));
  INV_X1    g0598(.A(G303), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n798), .A2(new_n724), .B1(new_n749), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n742), .A2(new_n519), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G311), .B2(new_n739), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n293), .B1(new_n736), .B2(G107), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n802), .A2(new_n760), .A3(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n797), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n716), .B1(new_n796), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n716), .A2(new_n713), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n806), .B(new_n704), .C1(G77), .C2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT99), .Z(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n714), .B2(new_n777), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n785), .A2(new_n811), .ZN(G384));
  AOI21_X1  g0612(.A(new_n215), .B1(G58), .B2(G68), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(new_n219), .B1(new_n202), .B2(G68), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n814), .A2(new_n248), .A3(G13), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT101), .Z(new_n816));
  XNOR2_X1  g0616(.A(new_n579), .B(KEYINPUT100), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n461), .B(new_n213), .C1(new_n817), .C2(KEYINPUT35), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(KEYINPUT35), .B2(new_n817), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT36), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  INV_X1    g0622(.A(new_n690), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n497), .A2(new_n501), .A3(new_n503), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n646), .A2(new_n824), .A3(new_n605), .A4(new_n640), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n823), .B1(new_n825), .B2(KEYINPUT31), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n690), .A2(new_n692), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n371), .A2(new_n640), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n369), .A2(new_n373), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT102), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n373), .A2(new_n352), .A3(new_n356), .A4(new_n358), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n829), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n369), .A2(new_n832), .A3(new_n373), .A4(new_n830), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n828), .A2(new_n778), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n440), .A2(new_n451), .A3(new_n453), .ZN(new_n839));
  INV_X1    g0639(.A(new_n424), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n409), .A2(new_n411), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT78), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n399), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(KEYINPUT16), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n256), .B1(new_n844), .B2(KEYINPUT16), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(new_n637), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n839), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n637), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n448), .B(new_n449), .C1(new_n445), .C2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n436), .A2(new_n852), .A3(new_n438), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n847), .B1(new_n443), .B2(new_n637), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n439), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT38), .B1(new_n849), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n849), .A2(KEYINPUT38), .A3(new_n857), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT40), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n838), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n439), .A2(KEYINPUT17), .ZN(new_n865));
  INV_X1    g0665(.A(new_n434), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n620), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n448), .A2(new_n449), .A3(new_n850), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT104), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n433), .B2(new_n619), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n420), .A2(KEYINPUT80), .A3(new_n376), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT80), .B1(new_n420), .B2(new_n376), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n840), .B1(new_n875), .B2(new_n846), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n435), .B(KEYINPUT104), .C1(new_n876), .C2(new_n443), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n872), .A2(new_n868), .A3(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .B1(new_n851), .B2(new_n853), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n870), .B1(new_n879), .B2(KEYINPUT105), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n881), .A2(KEYINPUT105), .A3(new_n854), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n864), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n860), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n838), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n863), .B1(new_n885), .B2(new_n862), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n460), .A2(new_n828), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n677), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n887), .B2(new_n886), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT106), .Z(new_n890));
  NAND3_X1  g0690(.A1(new_n859), .A2(KEYINPUT39), .A3(new_n860), .ZN(new_n891));
  AOI221_X4 g0691(.A(new_n864), .B1(new_n854), .B2(new_n856), .C1(new_n839), .C2(new_n848), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n881), .A2(new_n854), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT105), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n879), .A2(KEYINPUT105), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n896), .A3(new_n870), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n892), .B1(new_n897), .B2(new_n864), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n891), .B1(new_n898), .B2(KEYINPUT39), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n369), .A2(new_n639), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT103), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n620), .A2(new_n850), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n336), .A2(new_n639), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n780), .B2(new_n777), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n837), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n904), .B1(new_n907), .B2(new_n861), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n459), .A2(new_n676), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n622), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n909), .B(new_n911), .Z(new_n912));
  NAND2_X1  g0712(.A1(new_n890), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(G1), .B1(new_n700), .B2(G20), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(KEYINPUT107), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n890), .B2(new_n912), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT107), .B1(new_n913), .B2(new_n914), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n822), .B1(new_n916), .B2(new_n917), .ZN(G367));
  INV_X1    g0718(.A(new_n709), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n234), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n717), .B1(new_n207), .B2(new_n311), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n704), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(G50), .A2(new_n744), .B1(new_n728), .B2(G159), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n293), .B1(new_n735), .B2(new_n793), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(G137), .B2(new_n739), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n219), .A2(new_n791), .B1(new_n752), .B2(G68), .ZN(new_n926));
  AOI22_X1  g0726(.A1(G143), .A2(new_n750), .B1(new_n725), .B2(G150), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n923), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(G317), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n794), .A2(new_n536), .B1(new_n738), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT46), .B1(new_n736), .B2(G116), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n736), .A2(KEYINPUT46), .A3(G116), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n933), .B1(new_n745), .B2(new_n741), .C1(new_n798), .C2(new_n729), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n410), .B1(G97), .B2(new_n791), .ZN(new_n935));
  OAI221_X1 g0735(.A(new_n935), .B1(new_n799), .B2(new_n724), .C1(new_n746), .C2(new_n749), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n928), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT47), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n922), .B1(new_n938), .B2(new_n716), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n570), .A2(new_n640), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n573), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n940), .A2(new_n565), .A3(new_n566), .A4(new_n555), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(new_n715), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n602), .B(new_n604), .C1(new_n584), .C2(new_n640), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n602), .B2(new_n640), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n653), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n653), .A2(new_n947), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT45), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT110), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n949), .A2(new_n650), .A3(new_n952), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n650), .B1(new_n949), .B2(new_n952), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n649), .A2(new_n651), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n652), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n644), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n698), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT111), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(KEYINPUT111), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n953), .A2(new_n954), .A3(new_n650), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n958), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n698), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n656), .B(KEYINPUT41), .Z(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT112), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT112), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n971), .B(new_n968), .C1(new_n966), .C2(new_n698), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n702), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n652), .A2(new_n947), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT42), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT108), .Z(new_n976));
  OR2_X1    g0776(.A1(new_n946), .A2(new_n608), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n639), .B1(new_n977), .B2(new_n602), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n974), .B2(KEYINPUT42), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n941), .A2(new_n942), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT43), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT109), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n983), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n984), .B2(new_n986), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n645), .A2(new_n649), .A3(new_n947), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n988), .B(new_n989), .Z(new_n990));
  AOI21_X1  g0790(.A(new_n945), .B1(new_n973), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(G387));
  OR2_X1    g0792(.A1(new_n649), .A2(new_n770), .ZN(new_n993));
  INV_X1    g0793(.A(new_n658), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(new_n207), .A3(new_n293), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(G107), .B2(new_n207), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT113), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n239), .A2(new_n279), .ZN(new_n998));
  AOI211_X1 g0798(.A(G45), .B(new_n994), .C1(G68), .C2(G77), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n263), .A2(G50), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT50), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n919), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n997), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n717), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n704), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n467), .A2(new_n742), .B1(new_n738), .B2(new_n787), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n485), .B(new_n1006), .C1(new_n219), .C2(new_n736), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT114), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n750), .A2(G159), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n794), .A2(new_n311), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n725), .B2(G50), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G68), .A2(new_n744), .B1(new_n728), .B2(new_n264), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n739), .A2(G326), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n410), .B1(G116), .B2(new_n791), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n794), .A2(new_n741), .B1(new_n735), .B2(new_n798), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G317), .A2(new_n725), .B1(new_n750), .B2(G322), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n745), .B2(new_n799), .C1(new_n746), .C2(new_n729), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT48), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n1019), .B2(new_n1018), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT49), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1014), .B(new_n1015), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1013), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1005), .B1(new_n1025), .B2(new_n716), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n961), .A2(new_n703), .B1(new_n993), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n962), .A2(new_n656), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n961), .A2(new_n698), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(G393));
  NOR2_X1   g0830(.A1(new_n956), .A2(new_n957), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n657), .B1(new_n1032), .B2(new_n962), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1033), .A2(new_n966), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n717), .B1(new_n467), .B2(new_n207), .C1(new_n919), .C2(new_n243), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n704), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n293), .B(new_n763), .C1(G283), .C2(new_n736), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G322), .A2(new_n739), .B1(new_n752), .B2(G116), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n798), .B2(new_n745), .C1(new_n799), .C2(new_n729), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n746), .A2(new_n724), .B1(new_n749), .B2(new_n929), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT52), .Z(new_n1042));
  OAI22_X1  g0842(.A1(new_n787), .A2(new_n749), .B1(new_n724), .B2(new_n756), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT51), .Z(new_n1044));
  INV_X1    g0844(.A(G77), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n794), .A2(new_n1045), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n801), .B(new_n1046), .C1(G143), .C2(new_n739), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n485), .B1(G68), .B2(new_n736), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G50), .A2(new_n728), .B1(new_n744), .B2(new_n264), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1040), .A2(new_n1042), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1036), .B1(new_n1051), .B2(new_n716), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n947), .B2(new_n770), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1032), .B2(new_n702), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1034), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(G390));
  OAI21_X1  g0856(.A(new_n902), .B1(new_n906), .B2(new_n837), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT39), .B1(new_n883), .B2(new_n860), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT39), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n892), .A2(new_n858), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1057), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n835), .A2(new_n777), .A3(new_n836), .ZN(new_n1062));
  OAI211_X1 g0862(.A(G330), .B(new_n1062), .C1(new_n826), .C2(new_n695), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT115), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n905), .B1(new_n674), .B2(new_n777), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n902), .B1(new_n1065), .B2(new_n837), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n898), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1065), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n837), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n901), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT115), .B1(new_n884), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1061), .B(new_n1063), .C1(new_n1067), .C2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1064), .B1(new_n898), .B2(new_n1066), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n884), .A2(new_n1070), .A3(KEYINPUT115), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n899), .A2(new_n1057), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n827), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n677), .B1(new_n693), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n1062), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1072), .B(KEYINPUT116), .C1(new_n1075), .C2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1061), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT116), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1078), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n906), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1069), .B1(new_n697), .B2(new_n777), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1085), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1068), .B1(new_n697), .B2(new_n1062), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT117), .ZN(new_n1089));
  OAI211_X1 g0889(.A(G330), .B(new_n777), .C1(new_n826), .C2(new_n827), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n837), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1089), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1087), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n459), .A2(new_n1077), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n910), .A2(new_n1095), .A3(new_n622), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT118), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n1084), .B2(new_n1098), .ZN(new_n1100));
  AOI211_X1 g0900(.A(KEYINPUT118), .B(new_n1097), .C1(new_n1079), .C2(new_n1083), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n656), .B1(new_n1084), .B2(new_n1098), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n745), .A2(new_n1103), .B1(new_n756), .B2(new_n794), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G137), .B2(new_n728), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT119), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n290), .B1(new_n739), .B2(G125), .ZN(new_n1107));
  INV_X1    g0907(.A(G128), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1107), .B1(new_n749), .B2(new_n1108), .ZN(new_n1109));
  OR3_X1    g0909(.A1(new_n735), .A2(KEYINPUT53), .A3(new_n787), .ZN(new_n1110));
  OAI21_X1  g0910(.A(KEYINPUT53), .B1(new_n735), .B2(new_n787), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n202), .C2(new_n742), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1109), .B(new_n1112), .C1(G132), .C2(new_n725), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n461), .A2(new_n724), .B1(new_n749), .B2(new_n741), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n290), .B1(new_n735), .B2(new_n519), .C1(new_n217), .C2(new_n742), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n738), .A2(new_n798), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1114), .A2(new_n1115), .A3(new_n1046), .A4(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G97), .A2(new_n744), .B1(new_n728), .B2(G107), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1106), .A2(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n704), .B1(new_n264), .B2(new_n808), .C1(new_n1119), .C2(new_n720), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n899), .B2(new_n713), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n1084), .B2(new_n703), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1102), .A2(new_n1122), .ZN(G378));
  OAI21_X1  g0923(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n273), .A2(new_n850), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n310), .B(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n886), .B2(G330), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n886), .A2(G330), .A3(new_n1128), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1130), .A2(new_n1131), .B1(new_n903), .B2(new_n908), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1131), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1133), .A2(new_n909), .A3(new_n1129), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1124), .A2(KEYINPUT57), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n656), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT57), .B1(new_n1124), .B2(new_n1135), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1128), .A2(new_n714), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n704), .B1(new_n808), .B2(G50), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n410), .A2(G41), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n461), .B2(new_n749), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n742), .A2(new_n793), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G283), .B2(new_n739), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n217), .B2(new_n794), .C1(new_n220), .C2(new_n735), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G97), .B2(new_n728), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n311), .B2(new_n745), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1143), .B(new_n1148), .C1(G107), .C2(new_n725), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1149), .A2(KEYINPUT58), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n750), .A2(G125), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n794), .A2(new_n787), .B1(new_n735), .B2(new_n1103), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n725), .B2(G128), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G132), .A2(new_n728), .B1(new_n744), .B2(G137), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1151), .B(new_n1153), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G33), .B(G41), .C1(new_n791), .C2(G159), .ZN(new_n1160));
  INV_X1    g0960(.A(G124), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1160), .B1(new_n1161), .B2(new_n738), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT121), .Z(new_n1163));
  NAND3_X1  g0963(.A1(new_n1158), .A2(new_n1159), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1149), .A2(KEYINPUT58), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1142), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1150), .A2(new_n1164), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1141), .B1(new_n1168), .B2(new_n716), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1140), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n702), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1139), .A2(new_n1173), .ZN(G375));
  OR2_X1    g0974(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n969), .A3(new_n1097), .ZN(new_n1176));
  INV_X1    g0976(.A(G137), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n410), .B1(new_n756), .B2(new_n735), .C1(new_n724), .C2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n738), .A2(new_n1108), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1144), .B(new_n1179), .C1(G50), .C2(new_n752), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n745), .B2(new_n787), .C1(new_n729), .C2(new_n1103), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1178), .B(new_n1181), .C1(G132), .C2(new_n750), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n293), .B(new_n1010), .C1(G97), .C2(new_n736), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n1045), .B2(new_n742), .C1(new_n799), .C2(new_n738), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n741), .A2(new_n724), .B1(new_n749), .B2(new_n798), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n536), .A2(new_n745), .B1(new_n729), .B2(new_n461), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n716), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n707), .B1(new_n217), .B2(new_n807), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n1069), .C2(new_n714), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1094), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1176), .B(new_n1190), .C1(new_n702), .C2(new_n1191), .ZN(G381));
  INV_X1    g0992(.A(G378), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1139), .A2(new_n1193), .A3(new_n1173), .ZN(new_n1194));
  OR2_X1    g0994(.A1(G393), .A2(G396), .ZN(new_n1195));
  OR3_X1    g0995(.A1(G381), .A2(G384), .A3(new_n1195), .ZN(new_n1196));
  OR4_X1    g0996(.A1(G387), .A2(new_n1194), .A3(G390), .A4(new_n1196), .ZN(G407));
  OAI211_X1 g0997(.A(G407), .B(G213), .C1(G343), .C2(new_n1194), .ZN(G409));
  INV_X1    g0998(.A(KEYINPUT122), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1200));
  AOI211_X1 g1000(.A(KEYINPUT116), .B(new_n1078), .C1(new_n1200), .C2(new_n1061), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1081), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1201), .B1(new_n1072), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT118), .B1(new_n1203), .B2(new_n1097), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1084), .A2(new_n1099), .A3(new_n1098), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1171), .B1(new_n1206), .B2(new_n1096), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1172), .B1(new_n1207), .B2(new_n969), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1199), .B1(new_n1208), .B2(G378), .ZN(new_n1209));
  OAI211_X1 g1009(.A(G378), .B(new_n1173), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1124), .A2(new_n969), .A3(new_n1135), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1173), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1193), .A2(new_n1212), .A3(KEYINPUT122), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1209), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n638), .A2(G213), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT123), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1190), .B1(G384), .B2(new_n1216), .C1(new_n1191), .C2(new_n702), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT60), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1175), .B1(new_n1098), .B2(new_n1218), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1094), .A2(new_n1096), .A3(new_n1218), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(new_n657), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1217), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(G384), .A2(new_n1216), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1214), .A2(new_n1215), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT62), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n638), .A2(G213), .A3(G2897), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1224), .B(new_n1228), .Z(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT61), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT62), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1214), .A2(new_n1232), .A3(new_n1215), .A4(new_n1224), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1226), .A2(new_n1230), .A3(new_n1231), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT125), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G387), .A2(G390), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(G393), .B(new_n772), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(KEYINPUT124), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n991), .B2(new_n1055), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(KEYINPUT124), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1236), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1235), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n991), .A2(new_n1055), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n991), .A2(new_n1055), .ZN(new_n1245));
  OAI211_X1 g1045(.A(KEYINPUT124), .B(new_n1237), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1236), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1247), .A3(KEYINPUT125), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1243), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1234), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT61), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1225), .A2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1214), .A2(KEYINPUT63), .A3(new_n1215), .A4(new_n1224), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1250), .A2(new_n1256), .ZN(G405));
  NAND2_X1  g1057(.A1(G375), .A2(new_n1193), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1224), .A2(KEYINPUT126), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1259), .A2(KEYINPUT127), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(KEYINPUT127), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1258), .A2(new_n1210), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1262), .B1(new_n1258), .B2(new_n1210), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1249), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1265), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1267), .A2(new_n1248), .A3(new_n1243), .A4(new_n1263), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(G402));
endmodule


