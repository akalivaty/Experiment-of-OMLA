

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U552 ( .A1(n530), .A2(n529), .ZN(n536) );
  AND2_X1 U553 ( .A1(n531), .A2(n532), .ZN(n530) );
  NAND2_X1 U554 ( .A1(n535), .A2(n534), .ZN(n529) );
  NAND2_X1 U555 ( .A1(n801), .A2(n551), .ZN(n802) );
  NAND2_X1 U556 ( .A1(n540), .A2(n519), .ZN(n537) );
  AND2_X1 U557 ( .A1(n546), .A2(n545), .ZN(n758) );
  NOR2_X1 U558 ( .A1(n723), .A2(n947), .ZN(n725) );
  AND2_X2 U559 ( .A1(n714), .A2(n713), .ZN(n717) );
  NOR2_X1 U560 ( .A1(n997), .A2(n523), .ZN(n719) );
  NOR2_X1 U561 ( .A1(n602), .A2(n601), .ZN(n604) );
  AND2_X2 U562 ( .A1(n526), .A2(n525), .ZN(n524) );
  NOR2_X2 U563 ( .A1(G543), .A2(G651), .ZN(n673) );
  AND2_X2 U564 ( .A1(n712), .A2(G40), .ZN(n713) );
  OR2_X2 U565 ( .A1(G164), .A2(G1384), .ZN(n523) );
  AND2_X4 U566 ( .A1(G2104), .A2(G2105), .ZN(n564) );
  NOR2_X4 U567 ( .A1(G2104), .A2(n559), .ZN(n902) );
  NAND2_X1 U568 ( .A1(n528), .A2(n559), .ZN(n527) );
  XNOR2_X2 U569 ( .A(n784), .B(KEYINPUT98), .ZN(n795) );
  XNOR2_X2 U570 ( .A(n753), .B(KEYINPUT93), .ZN(n735) );
  NOR2_X2 U571 ( .A1(n568), .A2(n567), .ZN(G164) );
  XNOR2_X1 U572 ( .A(n765), .B(KEYINPUT96), .ZN(n777) );
  NAND2_X1 U573 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U574 ( .A(n762), .B(KEYINPUT31), .ZN(n763) );
  AND2_X1 U575 ( .A1(n945), .A2(n787), .ZN(n788) );
  INV_X1 U576 ( .A(n523), .ZN(n716) );
  NAND2_X1 U577 ( .A1(G2105), .A2(KEYINPUT17), .ZN(n525) );
  NAND2_X1 U578 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n526) );
  INV_X1 U579 ( .A(KEYINPUT94), .ZN(n726) );
  NOR2_X1 U580 ( .A1(n975), .A2(n737), .ZN(n738) );
  NOR2_X1 U581 ( .A1(n753), .A2(G2084), .ZN(n755) );
  OR2_X1 U582 ( .A1(n549), .A2(n770), .ZN(n771) );
  AND2_X1 U583 ( .A1(n539), .A2(n520), .ZN(n538) );
  NOR2_X1 U584 ( .A1(n542), .A2(KEYINPUT33), .ZN(n541) );
  INV_X1 U585 ( .A(KEYINPUT13), .ZN(n598) );
  NOR2_X1 U586 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n528) );
  XNOR2_X1 U587 ( .A(n553), .B(KEYINPUT66), .ZN(n554) );
  NAND2_X1 U588 ( .A1(n908), .A2(G137), .ZN(n555) );
  AND2_X1 U589 ( .A1(n543), .A2(KEYINPUT64), .ZN(n519) );
  NAND2_X2 U590 ( .A1(n717), .A2(n716), .ZN(n753) );
  OR2_X1 U591 ( .A1(n541), .A2(n790), .ZN(n520) );
  AND2_X1 U592 ( .A1(n788), .A2(n544), .ZN(n521) );
  AND2_X1 U593 ( .A1(n521), .A2(n543), .ZN(n522) );
  AND2_X2 U594 ( .A1(n793), .A2(n963), .ZN(n552) );
  NOR2_X2 U595 ( .A1(n552), .A2(n802), .ZN(n804) );
  AND2_X1 U596 ( .A1(n717), .A2(n523), .ZN(n847) );
  NAND2_X4 U597 ( .A1(n527), .A2(n524), .ZN(n908) );
  NAND2_X1 U598 ( .A1(n836), .A2(n837), .ZN(n531) );
  AND2_X1 U599 ( .A1(n849), .A2(n533), .ZN(n532) );
  NAND2_X1 U600 ( .A1(n835), .A2(n837), .ZN(n533) );
  NOR2_X1 U601 ( .A1(n835), .A2(n837), .ZN(n534) );
  INV_X1 U602 ( .A(n836), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n791) );
  NAND2_X1 U605 ( .A1(n789), .A2(n522), .ZN(n539) );
  INV_X1 U606 ( .A(n789), .ZN(n540) );
  NOR2_X1 U607 ( .A1(n788), .A2(n544), .ZN(n542) );
  INV_X1 U608 ( .A(n790), .ZN(n543) );
  INV_X1 U609 ( .A(KEYINPUT64), .ZN(n544) );
  INV_X1 U610 ( .A(G168), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n547), .B(n757), .ZN(n546) );
  NAND2_X1 U612 ( .A1(n548), .A2(n775), .ZN(n547) );
  NOR2_X1 U613 ( .A1(n779), .A2(n549), .ZN(n548) );
  INV_X1 U614 ( .A(G8), .ZN(n549) );
  OR2_X1 U615 ( .A1(G301), .A2(n759), .ZN(n550) );
  OR2_X1 U616 ( .A1(n800), .A2(n756), .ZN(n551) );
  INV_X1 U617 ( .A(KEYINPUT30), .ZN(n757) );
  INV_X1 U618 ( .A(KEYINPUT29), .ZN(n746) );
  INV_X1 U619 ( .A(KEYINPUT92), .ZN(n754) );
  INV_X1 U620 ( .A(KEYINPUT32), .ZN(n773) );
  INV_X1 U621 ( .A(KEYINPUT101), .ZN(n803) );
  NAND2_X1 U622 ( .A1(n676), .A2(G56), .ZN(n600) );
  INV_X1 U623 ( .A(KEYINPUT102), .ZN(n837) );
  INV_X1 U624 ( .A(KEYINPUT1), .ZN(n575) );
  XOR2_X1 U625 ( .A(KEYINPUT15), .B(n611), .Z(n955) );
  AND2_X1 U626 ( .A1(n714), .A2(n712), .ZN(G160) );
  NAND2_X1 U627 ( .A1(n604), .A2(n603), .ZN(n947) );
  NOR2_X1 U628 ( .A1(n579), .A2(n578), .ZN(G171) );
  NAND2_X1 U629 ( .A1(n564), .A2(G113), .ZN(n553) );
  NAND2_X1 U630 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U631 ( .A(n556), .B(KEYINPUT67), .ZN(n558) );
  INV_X2 U632 ( .A(G2105), .ZN(n559) );
  NAND2_X1 U633 ( .A1(G125), .A2(n902), .ZN(n557) );
  AND2_X2 U634 ( .A1(n558), .A2(n557), .ZN(n714) );
  AND2_X4 U635 ( .A1(n559), .A2(G2104), .ZN(n910) );
  NAND2_X1 U636 ( .A1(G101), .A2(n910), .ZN(n560) );
  XOR2_X1 U637 ( .A(KEYINPUT23), .B(n560), .Z(n712) );
  NAND2_X1 U638 ( .A1(G138), .A2(n908), .ZN(n563) );
  NAND2_X1 U639 ( .A1(G102), .A2(n910), .ZN(n562) );
  NAND2_X1 U640 ( .A1(n563), .A2(n562), .ZN(n568) );
  NAND2_X1 U641 ( .A1(G126), .A2(n902), .ZN(n566) );
  NAND2_X1 U642 ( .A1(G114), .A2(n564), .ZN(n565) );
  NAND2_X1 U643 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U644 ( .A1(G90), .A2(n673), .ZN(n570) );
  XOR2_X1 U645 ( .A(KEYINPUT0), .B(G543), .Z(n656) );
  INV_X1 U646 ( .A(G651), .ZN(n574) );
  NOR2_X2 U647 ( .A1(n656), .A2(n574), .ZN(n670) );
  NAND2_X1 U648 ( .A1(G77), .A2(n670), .ZN(n569) );
  NAND2_X1 U649 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U650 ( .A(n571), .B(KEYINPUT9), .ZN(n573) );
  NOR2_X2 U651 ( .A1(n656), .A2(G651), .ZN(n672) );
  NAND2_X1 U652 ( .A1(G52), .A2(n672), .ZN(n572) );
  NAND2_X1 U653 ( .A1(n573), .A2(n572), .ZN(n579) );
  NOR2_X1 U654 ( .A1(G543), .A2(n574), .ZN(n576) );
  XNOR2_X2 U655 ( .A(n576), .B(n575), .ZN(n676) );
  NAND2_X1 U656 ( .A1(G64), .A2(n676), .ZN(n577) );
  XNOR2_X1 U657 ( .A(KEYINPUT69), .B(n577), .ZN(n578) );
  XNOR2_X1 U658 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U659 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U660 ( .A(G82), .ZN(G220) );
  INV_X1 U661 ( .A(G120), .ZN(G236) );
  INV_X1 U662 ( .A(G69), .ZN(G235) );
  INV_X1 U663 ( .A(G108), .ZN(G238) );
  NAND2_X1 U664 ( .A1(n673), .A2(G89), .ZN(n580) );
  XNOR2_X1 U665 ( .A(n580), .B(KEYINPUT4), .ZN(n582) );
  NAND2_X1 U666 ( .A1(G76), .A2(n670), .ZN(n581) );
  NAND2_X1 U667 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U668 ( .A(KEYINPUT5), .B(n583), .ZN(n589) );
  NAND2_X1 U669 ( .A1(G63), .A2(n676), .ZN(n585) );
  NAND2_X1 U670 ( .A1(G51), .A2(n672), .ZN(n584) );
  NAND2_X1 U671 ( .A1(n585), .A2(n584), .ZN(n587) );
  XOR2_X1 U672 ( .A(KEYINPUT6), .B(KEYINPUT74), .Z(n586) );
  XNOR2_X1 U673 ( .A(n587), .B(n586), .ZN(n588) );
  NAND2_X1 U674 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U675 ( .A(KEYINPUT7), .B(n590), .ZN(G168) );
  XOR2_X1 U676 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U677 ( .A1(G7), .A2(G661), .ZN(n591) );
  XNOR2_X1 U678 ( .A(n591), .B(KEYINPUT72), .ZN(n592) );
  XNOR2_X1 U679 ( .A(KEYINPUT10), .B(n592), .ZN(G223) );
  INV_X1 U680 ( .A(G223), .ZN(n850) );
  NAND2_X1 U681 ( .A1(n850), .A2(G567), .ZN(n593) );
  XNOR2_X1 U682 ( .A(n593), .B(KEYINPUT73), .ZN(n594) );
  XNOR2_X1 U683 ( .A(KEYINPUT11), .B(n594), .ZN(G234) );
  NAND2_X1 U684 ( .A1(G68), .A2(n670), .ZN(n597) );
  NAND2_X1 U685 ( .A1(n673), .A2(G81), .ZN(n595) );
  XNOR2_X1 U686 ( .A(n595), .B(KEYINPUT12), .ZN(n596) );
  NAND2_X1 U687 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U688 ( .A(n599), .B(n598), .ZN(n602) );
  XOR2_X1 U689 ( .A(KEYINPUT14), .B(n600), .Z(n601) );
  NAND2_X1 U690 ( .A1(n672), .A2(G43), .ZN(n603) );
  INV_X1 U691 ( .A(G860), .ZN(n624) );
  OR2_X1 U692 ( .A1(n947), .A2(n624), .ZN(G153) );
  INV_X1 U693 ( .A(G171), .ZN(G301) );
  NAND2_X1 U694 ( .A1(G868), .A2(G301), .ZN(n613) );
  NAND2_X1 U695 ( .A1(G66), .A2(n676), .ZN(n606) );
  NAND2_X1 U696 ( .A1(G92), .A2(n673), .ZN(n605) );
  NAND2_X1 U697 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U698 ( .A1(G54), .A2(n672), .ZN(n608) );
  NAND2_X1 U699 ( .A1(G79), .A2(n670), .ZN(n607) );
  NAND2_X1 U700 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U701 ( .A1(n610), .A2(n609), .ZN(n611) );
  OR2_X1 U702 ( .A1(n955), .A2(G868), .ZN(n612) );
  NAND2_X1 U703 ( .A1(n613), .A2(n612), .ZN(G284) );
  NAND2_X1 U704 ( .A1(G91), .A2(n673), .ZN(n615) );
  NAND2_X1 U705 ( .A1(G78), .A2(n670), .ZN(n614) );
  NAND2_X1 U706 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n672), .A2(G53), .ZN(n616) );
  XOR2_X1 U708 ( .A(KEYINPUT70), .B(n616), .Z(n617) );
  NOR2_X1 U709 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U710 ( .A1(n676), .A2(G65), .ZN(n619) );
  NAND2_X1 U711 ( .A1(n620), .A2(n619), .ZN(G299) );
  XNOR2_X1 U712 ( .A(KEYINPUT75), .B(G868), .ZN(n621) );
  NOR2_X1 U713 ( .A1(G286), .A2(n621), .ZN(n623) );
  NOR2_X1 U714 ( .A1(G868), .A2(G299), .ZN(n622) );
  NOR2_X1 U715 ( .A1(n623), .A2(n622), .ZN(G297) );
  NAND2_X1 U716 ( .A1(n624), .A2(G559), .ZN(n625) );
  NAND2_X1 U717 ( .A1(n625), .A2(n955), .ZN(n626) );
  XNOR2_X1 U718 ( .A(n626), .B(KEYINPUT16), .ZN(n627) );
  XNOR2_X1 U719 ( .A(KEYINPUT76), .B(n627), .ZN(G148) );
  NOR2_X1 U720 ( .A1(G868), .A2(n947), .ZN(n630) );
  NAND2_X1 U721 ( .A1(n955), .A2(G868), .ZN(n628) );
  NOR2_X1 U722 ( .A1(G559), .A2(n628), .ZN(n629) );
  NOR2_X1 U723 ( .A1(n630), .A2(n629), .ZN(G282) );
  NAND2_X1 U724 ( .A1(G123), .A2(n902), .ZN(n631) );
  XOR2_X1 U725 ( .A(KEYINPUT77), .B(n631), .Z(n632) );
  XNOR2_X1 U726 ( .A(n632), .B(KEYINPUT18), .ZN(n634) );
  NAND2_X1 U727 ( .A1(G111), .A2(n564), .ZN(n633) );
  NAND2_X1 U728 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U729 ( .A1(G135), .A2(n908), .ZN(n636) );
  NAND2_X1 U730 ( .A1(G99), .A2(n910), .ZN(n635) );
  NAND2_X1 U731 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U732 ( .A1(n638), .A2(n637), .ZN(n1027) );
  XNOR2_X1 U733 ( .A(n1027), .B(G2096), .ZN(n640) );
  INV_X1 U734 ( .A(G2100), .ZN(n639) );
  NAND2_X1 U735 ( .A1(n640), .A2(n639), .ZN(G156) );
  NAND2_X1 U736 ( .A1(n955), .A2(G559), .ZN(n690) );
  XNOR2_X1 U737 ( .A(n947), .B(n690), .ZN(n641) );
  NOR2_X1 U738 ( .A1(n641), .A2(G860), .ZN(n648) );
  NAND2_X1 U739 ( .A1(G67), .A2(n676), .ZN(n643) );
  NAND2_X1 U740 ( .A1(G93), .A2(n673), .ZN(n642) );
  NAND2_X1 U741 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U742 ( .A1(G55), .A2(n672), .ZN(n645) );
  NAND2_X1 U743 ( .A1(G80), .A2(n670), .ZN(n644) );
  NAND2_X1 U744 ( .A1(n645), .A2(n644), .ZN(n646) );
  OR2_X1 U745 ( .A1(n647), .A2(n646), .ZN(n693) );
  XOR2_X1 U746 ( .A(n648), .B(n693), .Z(G145) );
  NAND2_X1 U747 ( .A1(G60), .A2(n676), .ZN(n650) );
  NAND2_X1 U748 ( .A1(G47), .A2(n672), .ZN(n649) );
  NAND2_X1 U749 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U750 ( .A(KEYINPUT68), .B(n651), .Z(n655) );
  NAND2_X1 U751 ( .A1(G85), .A2(n673), .ZN(n653) );
  NAND2_X1 U752 ( .A1(G72), .A2(n670), .ZN(n652) );
  AND2_X1 U753 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U754 ( .A1(n655), .A2(n654), .ZN(G290) );
  NAND2_X1 U755 ( .A1(G49), .A2(n672), .ZN(n658) );
  NAND2_X1 U756 ( .A1(G87), .A2(n656), .ZN(n657) );
  NAND2_X1 U757 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U758 ( .A1(n676), .A2(n659), .ZN(n661) );
  NAND2_X1 U759 ( .A1(G651), .A2(G74), .ZN(n660) );
  NAND2_X1 U760 ( .A1(n661), .A2(n660), .ZN(G288) );
  NAND2_X1 U761 ( .A1(G86), .A2(n673), .ZN(n668) );
  NAND2_X1 U762 ( .A1(G61), .A2(n676), .ZN(n663) );
  NAND2_X1 U763 ( .A1(G48), .A2(n672), .ZN(n662) );
  NAND2_X1 U764 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U765 ( .A1(n670), .A2(G73), .ZN(n664) );
  XOR2_X1 U766 ( .A(KEYINPUT2), .B(n664), .Z(n665) );
  NOR2_X1 U767 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U768 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U769 ( .A(n669), .B(KEYINPUT78), .ZN(G305) );
  NAND2_X1 U770 ( .A1(G75), .A2(n670), .ZN(n671) );
  XNOR2_X1 U771 ( .A(n671), .B(KEYINPUT80), .ZN(n681) );
  NAND2_X1 U772 ( .A1(G50), .A2(n672), .ZN(n675) );
  NAND2_X1 U773 ( .A1(G88), .A2(n673), .ZN(n674) );
  NAND2_X1 U774 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U775 ( .A1(G62), .A2(n676), .ZN(n677) );
  XNOR2_X1 U776 ( .A(KEYINPUT79), .B(n677), .ZN(n678) );
  NOR2_X1 U777 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U778 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U779 ( .A(KEYINPUT81), .B(n682), .ZN(G166) );
  XNOR2_X1 U780 ( .A(KEYINPUT19), .B(G290), .ZN(n683) );
  XNOR2_X1 U781 ( .A(n683), .B(G288), .ZN(n684) );
  XNOR2_X1 U782 ( .A(KEYINPUT82), .B(n684), .ZN(n686) );
  XNOR2_X1 U783 ( .A(n947), .B(G305), .ZN(n685) );
  XNOR2_X1 U784 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U785 ( .A(n687), .B(n693), .ZN(n689) );
  INV_X1 U786 ( .A(G299), .ZN(n944) );
  XNOR2_X1 U787 ( .A(G166), .B(n944), .ZN(n688) );
  XNOR2_X1 U788 ( .A(n689), .B(n688), .ZN(n922) );
  XNOR2_X1 U789 ( .A(KEYINPUT83), .B(n690), .ZN(n691) );
  XNOR2_X1 U790 ( .A(n922), .B(n691), .ZN(n692) );
  NAND2_X1 U791 ( .A1(n692), .A2(G868), .ZN(n696) );
  INV_X1 U792 ( .A(G868), .ZN(n694) );
  NAND2_X1 U793 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U794 ( .A1(n696), .A2(n695), .ZN(G295) );
  NAND2_X1 U795 ( .A1(G2078), .A2(G2084), .ZN(n697) );
  XOR2_X1 U796 ( .A(KEYINPUT20), .B(n697), .Z(n698) );
  NAND2_X1 U797 ( .A1(G2090), .A2(n698), .ZN(n699) );
  XNOR2_X1 U798 ( .A(KEYINPUT21), .B(n699), .ZN(n700) );
  NAND2_X1 U799 ( .A1(n700), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U800 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U801 ( .A1(G235), .A2(G236), .ZN(n701) );
  XOR2_X1 U802 ( .A(KEYINPUT84), .B(n701), .Z(n702) );
  NOR2_X1 U803 ( .A1(G238), .A2(n702), .ZN(n703) );
  NAND2_X1 U804 ( .A1(G57), .A2(n703), .ZN(n854) );
  NAND2_X1 U805 ( .A1(G567), .A2(n854), .ZN(n704) );
  XNOR2_X1 U806 ( .A(n704), .B(KEYINPUT85), .ZN(n709) );
  NOR2_X1 U807 ( .A1(G220), .A2(G219), .ZN(n705) );
  XNOR2_X1 U808 ( .A(KEYINPUT22), .B(n705), .ZN(n706) );
  NAND2_X1 U809 ( .A1(n706), .A2(G96), .ZN(n707) );
  OR2_X1 U810 ( .A1(G218), .A2(n707), .ZN(n855) );
  AND2_X1 U811 ( .A1(G2106), .A2(n855), .ZN(n708) );
  NOR2_X1 U812 ( .A1(n709), .A2(n708), .ZN(G319) );
  INV_X1 U813 ( .A(G319), .ZN(n711) );
  NAND2_X1 U814 ( .A1(G483), .A2(G661), .ZN(n710) );
  NOR2_X1 U815 ( .A1(n711), .A2(n710), .ZN(n853) );
  NAND2_X1 U816 ( .A1(n853), .A2(G36), .ZN(G176) );
  INV_X1 U817 ( .A(G166), .ZN(G303) );
  NAND2_X1 U818 ( .A1(n753), .A2(G8), .ZN(n756) );
  INV_X1 U819 ( .A(n756), .ZN(n787) );
  NOR2_X1 U820 ( .A1(G1976), .A2(G288), .ZN(n948) );
  NAND2_X1 U821 ( .A1(n787), .A2(n948), .ZN(n718) );
  AND2_X1 U822 ( .A1(KEYINPUT33), .A2(n718), .ZN(n790) );
  INV_X1 U823 ( .A(G1996), .ZN(n997) );
  NAND2_X1 U824 ( .A1(n717), .A2(n719), .ZN(n720) );
  XNOR2_X1 U825 ( .A(n720), .B(KEYINPUT26), .ZN(n722) );
  NAND2_X1 U826 ( .A1(n753), .A2(G1341), .ZN(n721) );
  NAND2_X1 U827 ( .A1(n722), .A2(n721), .ZN(n723) );
  INV_X1 U828 ( .A(KEYINPUT65), .ZN(n724) );
  XNOR2_X1 U829 ( .A(n725), .B(n724), .ZN(n728) );
  NOR2_X1 U830 ( .A1(n728), .A2(n955), .ZN(n727) );
  XNOR2_X1 U831 ( .A(n727), .B(n726), .ZN(n734) );
  NAND2_X1 U832 ( .A1(n728), .A2(n955), .ZN(n732) );
  NAND2_X1 U833 ( .A1(G1348), .A2(n753), .ZN(n730) );
  BUF_X2 U834 ( .A(n735), .Z(n737) );
  NAND2_X1 U835 ( .A1(G2067), .A2(n737), .ZN(n729) );
  NAND2_X1 U836 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U837 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U838 ( .A1(n734), .A2(n733), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n735), .A2(G2072), .ZN(n736) );
  XNOR2_X1 U840 ( .A(n736), .B(KEYINPUT27), .ZN(n739) );
  INV_X1 U841 ( .A(G1956), .ZN(n975) );
  NOR2_X1 U842 ( .A1(n739), .A2(n738), .ZN(n742) );
  NAND2_X1 U843 ( .A1(n944), .A2(n742), .ZN(n740) );
  NAND2_X1 U844 ( .A1(n741), .A2(n740), .ZN(n745) );
  NOR2_X1 U845 ( .A1(n944), .A2(n742), .ZN(n743) );
  XOR2_X1 U846 ( .A(n743), .B(KEYINPUT28), .Z(n744) );
  NAND2_X1 U847 ( .A1(n745), .A2(n744), .ZN(n747) );
  XNOR2_X1 U848 ( .A(n747), .B(n746), .ZN(n752) );
  XOR2_X1 U849 ( .A(G2078), .B(KEYINPUT25), .Z(n1002) );
  INV_X1 U850 ( .A(n737), .ZN(n748) );
  NOR2_X1 U851 ( .A1(n1002), .A2(n748), .ZN(n751) );
  INV_X1 U852 ( .A(n753), .ZN(n749) );
  NOR2_X1 U853 ( .A1(n749), .A2(G1961), .ZN(n750) );
  NOR2_X1 U854 ( .A1(n751), .A2(n750), .ZN(n759) );
  NAND2_X1 U855 ( .A1(n752), .A2(n550), .ZN(n764) );
  XNOR2_X1 U856 ( .A(n755), .B(n754), .ZN(n775) );
  NOR2_X1 U857 ( .A1(G1966), .A2(n756), .ZN(n779) );
  XNOR2_X1 U858 ( .A(n758), .B(KEYINPUT95), .ZN(n761) );
  NAND2_X1 U859 ( .A1(n759), .A2(G301), .ZN(n760) );
  NAND2_X1 U860 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U861 ( .A1(n777), .A2(G286), .ZN(n772) );
  NOR2_X1 U862 ( .A1(G2090), .A2(n753), .ZN(n766) );
  XNOR2_X1 U863 ( .A(KEYINPUT97), .B(n766), .ZN(n769) );
  NOR2_X1 U864 ( .A1(G1971), .A2(n756), .ZN(n767) );
  NOR2_X1 U865 ( .A1(G166), .A2(n767), .ZN(n768) );
  NAND2_X1 U866 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U867 ( .A1(n772), .A2(n771), .ZN(n774) );
  XNOR2_X1 U868 ( .A(n774), .B(n773), .ZN(n783) );
  INV_X1 U869 ( .A(n775), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n776), .A2(G8), .ZN(n781) );
  INV_X1 U871 ( .A(n777), .ZN(n778) );
  NOR2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U875 ( .A1(G1971), .A2(G303), .ZN(n785) );
  NOR2_X1 U876 ( .A1(n785), .A2(n948), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n795), .A2(n786), .ZN(n789) );
  NAND2_X1 U878 ( .A1(G1976), .A2(G288), .ZN(n945) );
  XNOR2_X1 U879 ( .A(n791), .B(KEYINPUT99), .ZN(n793) );
  XOR2_X1 U880 ( .A(G1981), .B(G305), .Z(n792) );
  XNOR2_X1 U881 ( .A(KEYINPUT100), .B(n792), .ZN(n963) );
  NOR2_X1 U882 ( .A1(G2090), .A2(G303), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G8), .A2(n794), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n797), .A2(n756), .ZN(n801) );
  NOR2_X1 U886 ( .A1(G1981), .A2(G305), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n798), .B(KEYINPUT91), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n799), .B(KEYINPUT24), .ZN(n800) );
  XNOR2_X1 U889 ( .A(n804), .B(n803), .ZN(n836) );
  NAND2_X1 U890 ( .A1(G105), .A2(n910), .ZN(n805) );
  XNOR2_X1 U891 ( .A(n805), .B(KEYINPUT38), .ZN(n812) );
  NAND2_X1 U892 ( .A1(G129), .A2(n902), .ZN(n807) );
  NAND2_X1 U893 ( .A1(G117), .A2(n564), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U895 ( .A1(G141), .A2(n908), .ZN(n808) );
  XNOR2_X1 U896 ( .A(KEYINPUT89), .B(n808), .ZN(n809) );
  NOR2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U898 ( .A1(n812), .A2(n811), .ZN(n899) );
  NAND2_X1 U899 ( .A1(G1996), .A2(n899), .ZN(n813) );
  XNOR2_X1 U900 ( .A(n813), .B(KEYINPUT90), .ZN(n823) );
  XNOR2_X1 U901 ( .A(KEYINPUT88), .B(G1991), .ZN(n1001) );
  NAND2_X1 U902 ( .A1(n902), .A2(G119), .ZN(n820) );
  NAND2_X1 U903 ( .A1(G95), .A2(n910), .ZN(n815) );
  NAND2_X1 U904 ( .A1(G107), .A2(n564), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n815), .A2(n814), .ZN(n818) );
  NAND2_X1 U906 ( .A1(n908), .A2(G131), .ZN(n816) );
  XOR2_X1 U907 ( .A(KEYINPUT86), .B(n816), .Z(n817) );
  NOR2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U910 ( .A(KEYINPUT87), .B(n821), .Z(n918) );
  NAND2_X1 U911 ( .A1(n1001), .A2(n918), .ZN(n822) );
  NAND2_X1 U912 ( .A1(n823), .A2(n822), .ZN(n840) );
  INV_X1 U913 ( .A(n840), .ZN(n1021) );
  XOR2_X1 U914 ( .A(G1986), .B(G290), .Z(n954) );
  NAND2_X1 U915 ( .A1(n1021), .A2(n954), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n824), .A2(n847), .ZN(n834) );
  XNOR2_X1 U917 ( .A(KEYINPUT37), .B(G2067), .ZN(n845) );
  NAND2_X1 U918 ( .A1(G140), .A2(n908), .ZN(n826) );
  NAND2_X1 U919 ( .A1(G104), .A2(n910), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U921 ( .A(KEYINPUT34), .B(n827), .ZN(n832) );
  NAND2_X1 U922 ( .A1(G128), .A2(n902), .ZN(n829) );
  NAND2_X1 U923 ( .A1(G116), .A2(n564), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U925 ( .A(KEYINPUT35), .B(n830), .Z(n831) );
  NOR2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U927 ( .A(KEYINPUT36), .B(n833), .ZN(n915) );
  NOR2_X1 U928 ( .A1(n845), .A2(n915), .ZN(n1023) );
  NAND2_X1 U929 ( .A1(n847), .A2(n1023), .ZN(n843) );
  NAND2_X1 U930 ( .A1(n834), .A2(n843), .ZN(n835) );
  NOR2_X1 U931 ( .A1(G1996), .A2(n899), .ZN(n1032) );
  NOR2_X1 U932 ( .A1(n1001), .A2(n918), .ZN(n1022) );
  NOR2_X1 U933 ( .A1(G1986), .A2(G290), .ZN(n838) );
  NOR2_X1 U934 ( .A1(n1022), .A2(n838), .ZN(n839) );
  NOR2_X1 U935 ( .A1(n840), .A2(n839), .ZN(n841) );
  NOR2_X1 U936 ( .A1(n1032), .A2(n841), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n842), .B(KEYINPUT39), .ZN(n844) );
  NAND2_X1 U938 ( .A1(n844), .A2(n843), .ZN(n846) );
  NAND2_X1 U939 ( .A1(n845), .A2(n915), .ZN(n1020) );
  NAND2_X1 U940 ( .A1(n846), .A2(n1020), .ZN(n848) );
  NAND2_X1 U941 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n850), .ZN(G217) );
  AND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U944 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U945 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U946 ( .A1(n853), .A2(n852), .ZN(G188) );
  INV_X1 U948 ( .A(G96), .ZN(G221) );
  NOR2_X1 U949 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U950 ( .A(KEYINPUT104), .B(n856), .ZN(G325) );
  INV_X1 U951 ( .A(G325), .ZN(G261) );
  XOR2_X1 U952 ( .A(KEYINPUT105), .B(G2678), .Z(n858) );
  XNOR2_X1 U953 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U955 ( .A(KEYINPUT42), .B(G2072), .Z(n860) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2090), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U958 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U959 ( .A(G2096), .B(G2100), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(n866) );
  XOR2_X1 U961 ( .A(G2078), .B(G2084), .Z(n865) );
  XNOR2_X1 U962 ( .A(n866), .B(n865), .ZN(G227) );
  XOR2_X1 U963 ( .A(G1976), .B(G1971), .Z(n868) );
  XNOR2_X1 U964 ( .A(G1986), .B(G1961), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U966 ( .A(n869), .B(G2474), .Z(n871) );
  XNOR2_X1 U967 ( .A(G1996), .B(G1991), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U969 ( .A(KEYINPUT41), .B(G1981), .Z(n873) );
  XNOR2_X1 U970 ( .A(G1966), .B(G1956), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(G229) );
  NAND2_X1 U973 ( .A1(G124), .A2(n902), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n876), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G136), .A2(n908), .ZN(n877) );
  XOR2_X1 U976 ( .A(KEYINPUT107), .B(n877), .Z(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U978 ( .A1(G100), .A2(n910), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G112), .A2(n564), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U981 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U982 ( .A1(G130), .A2(n902), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G118), .A2(n564), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n891) );
  NAND2_X1 U985 ( .A1(G142), .A2(n908), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G106), .A2(n910), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U988 ( .A(KEYINPUT45), .B(n888), .Z(n889) );
  XNOR2_X1 U989 ( .A(KEYINPUT108), .B(n889), .ZN(n890) );
  NOR2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n901) );
  XOR2_X1 U991 ( .A(KEYINPUT113), .B(KEYINPUT109), .Z(n893) );
  XNOR2_X1 U992 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U994 ( .A(n894), .B(KEYINPUT114), .Z(n896) );
  XNOR2_X1 U995 ( .A(G164), .B(G162), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U997 ( .A(n1027), .B(n897), .Z(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n917) );
  XNOR2_X1 U1000 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n902), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(G115), .A2(n564), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n905), .B(KEYINPUT47), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n914) );
  NAND2_X1 U1006 ( .A1(n908), .A2(G139), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n909), .B(KEYINPUT110), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(G103), .A2(n910), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n1037) );
  XNOR2_X1 U1011 ( .A(n915), .B(n1037), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n920) );
  XOR2_X1 U1013 ( .A(G160), .B(n918), .Z(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n921), .ZN(G395) );
  XOR2_X1 U1016 ( .A(KEYINPUT115), .B(n922), .Z(n924) );
  XNOR2_X1 U1017 ( .A(n955), .B(G286), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(n924), .B(n923), .ZN(n925) );
  XNOR2_X1 U1019 ( .A(G171), .B(n925), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(G37), .A2(n926), .ZN(G397) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n928), .B(n927), .ZN(n940) );
  XOR2_X1 U1024 ( .A(KEYINPUT103), .B(G2451), .Z(n930) );
  XNOR2_X1 U1025 ( .A(G2446), .B(G2427), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n930), .B(n929), .ZN(n937) );
  XOR2_X1 U1027 ( .A(G2438), .B(G2435), .Z(n932) );
  XNOR2_X1 U1028 ( .A(G2443), .B(G2430), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n932), .B(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(n933), .B(G2454), .Z(n935) );
  XNOR2_X1 U1031 ( .A(G1348), .B(G1341), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(n935), .B(n934), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(n937), .B(n936), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n938), .A2(G14), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(G319), .A2(n943), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(G395), .A2(G397), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(G225) );
  INV_X1 U1039 ( .A(G225), .ZN(G308) );
  INV_X1 U1040 ( .A(G57), .ZN(G237) );
  INV_X1 U1041 ( .A(n943), .ZN(G401) );
  XNOR2_X1 U1042 ( .A(KEYINPUT56), .B(G16), .ZN(n969) );
  XNOR2_X1 U1043 ( .A(n944), .B(G1956), .ZN(n946) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n952) );
  XOR2_X1 U1045 ( .A(n947), .B(G1341), .Z(n950) );
  XNOR2_X1 U1046 ( .A(n948), .B(KEYINPUT123), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n962) );
  XOR2_X1 U1050 ( .A(G1348), .B(n955), .Z(n957) );
  XOR2_X1 U1051 ( .A(G171), .B(G1961), .Z(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(KEYINPUT122), .B(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G166), .B(G1971), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G168), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n965), .B(KEYINPUT57), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n1050) );
  XOR2_X1 U1062 ( .A(G16), .B(KEYINPUT124), .Z(n995) );
  XNOR2_X1 U1063 ( .A(G1348), .B(KEYINPUT59), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(n970), .B(G4), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(G1341), .B(G19), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G1981), .B(G6), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n978) );
  XOR2_X1 U1069 ( .A(KEYINPUT126), .B(n975), .Z(n976) );
  XNOR2_X1 U1070 ( .A(G20), .B(n976), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(KEYINPUT60), .B(n979), .ZN(n989) );
  XOR2_X1 U1073 ( .A(G1966), .B(KEYINPUT127), .Z(n980) );
  XNOR2_X1 U1074 ( .A(G21), .B(n980), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(G1986), .B(G24), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(G1971), .B(G22), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n984) );
  XOR2_X1 U1078 ( .A(G1976), .B(G23), .Z(n983) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT58), .B(n985), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n992) );
  XOR2_X1 U1083 ( .A(KEYINPUT125), .B(G1961), .Z(n990) );
  XNOR2_X1 U1084 ( .A(G5), .B(n990), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n993), .B(KEYINPUT61), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(G11), .A2(n996), .ZN(n1048) );
  XNOR2_X1 U1089 ( .A(G32), .B(n997), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n998), .A2(G28), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(G2067), .B(G26), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(G33), .B(G2072), .ZN(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(n1001), .B(G25), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(G27), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT53), .B(n1009), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT119), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(G2090), .B(G35), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n1011) );
  XNOR2_X1 U1103 ( .A(n1011), .B(G34), .ZN(n1012) );
  XNOR2_X1 U1104 ( .A(n1012), .B(G2084), .ZN(n1013) );
  NOR2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(KEYINPUT121), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(G29), .A2(n1018), .ZN(n1019) );
  XNOR2_X1 U1109 ( .A(n1019), .B(KEYINPUT55), .ZN(n1046) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1030) );
  XNOR2_X1 U1111 ( .A(G160), .B(G2084), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(KEYINPUT117), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1036) );
  XOR2_X1 U1117 ( .A(G2090), .B(G162), .Z(n1031) );
  XNOR2_X1 U1118 ( .A(KEYINPUT118), .B(n1031), .ZN(n1033) );
  NOR2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1120 ( .A(KEYINPUT51), .B(n1034), .Z(n1035) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1042) );
  XOR2_X1 U1122 ( .A(G2072), .B(n1037), .Z(n1039) );
  XOR2_X1 U1123 ( .A(G164), .B(G2078), .Z(n1038) );
  NOR2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XOR2_X1 U1125 ( .A(KEYINPUT50), .B(n1040), .Z(n1041) );
  NOR2_X1 U1126 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XOR2_X1 U1127 ( .A(KEYINPUT52), .B(n1043), .Z(n1044) );
  NAND2_X1 U1128 ( .A1(G29), .A2(n1044), .ZN(n1045) );
  NAND2_X1 U1129 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NOR2_X1 U1130 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NAND2_X1 U1131 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  XOR2_X1 U1132 ( .A(KEYINPUT62), .B(n1051), .Z(G311) );
  INV_X1 U1133 ( .A(G311), .ZN(G150) );
endmodule

