//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n621, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n454), .A2(new_n458), .B1(new_n449), .B2(new_n455), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(KEYINPUT67), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n461), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  AOI21_X1  g049(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n461), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(G136), .B2(new_n467), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(G162));
  NOR2_X1   g056(.A1(new_n461), .A2(G114), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n475), .B2(G126), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n467), .A2(new_n487), .A3(G138), .ZN(new_n488));
  INV_X1    g063(.A(new_n466), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n461), .C1(new_n489), .C2(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT70), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n471), .A2(new_n493), .A3(G138), .A4(new_n461), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n486), .B1(new_n492), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(KEYINPUT5), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(new_n497), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n496), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n511), .B1(new_n509), .B2(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .A3(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n497), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n514), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n510), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  AOI22_X1  g098(.A1(new_n500), .A2(new_n506), .B1(new_n512), .B2(new_n514), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(G89), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(KEYINPUT75), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(KEYINPUT75), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n515), .A2(G51), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n507), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n507), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR3_X1   g108(.A1(new_n526), .A2(new_n527), .A3(new_n533), .ZN(G168));
  NAND3_X1  g109(.A1(new_n507), .A2(G90), .A3(new_n517), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n515), .A2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n540), .B1(new_n507), .B2(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n538), .B1(new_n541), .B2(new_n509), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n500), .B2(new_n506), .ZN(new_n544));
  OAI211_X1 g119(.A(KEYINPUT76), .B(G651), .C1(new_n544), .C2(new_n540), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n537), .B1(new_n542), .B2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n509), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT77), .B(G43), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n524), .A2(G81), .B1(new_n515), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n500), .B2(new_n506), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT78), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n564), .B(G651), .C1(new_n559), .C2(new_n561), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n515), .A2(G53), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n515), .A2(new_n569), .A3(G53), .ZN(new_n570));
  AOI22_X1  g145(.A1(G91), .A2(new_n524), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n566), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n542), .A2(new_n545), .ZN(new_n574));
  INV_X1    g149(.A(new_n537), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI211_X1 g151(.A(KEYINPUT79), .B(new_n537), .C1(new_n542), .C2(new_n545), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(G301));
  OR2_X1    g153(.A1(new_n525), .A2(KEYINPUT75), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n525), .A2(KEYINPUT75), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n531), .A2(new_n532), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n528), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT80), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n524), .A2(G87), .B1(G49), .B2(new_n515), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G288));
  AND2_X1   g162(.A1(new_n507), .A2(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT81), .Z(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n524), .A2(G86), .B1(G48), .B2(new_n515), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n524), .A2(G85), .B1(G47), .B2(new_n515), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n509), .B2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  NOR3_X1   g175(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n497), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT73), .B1(new_n501), .B2(G543), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n505), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n600), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(G54), .B2(new_n515), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n518), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  AOI21_X1  g189(.A(KEYINPUT82), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n599), .B1(new_n597), .B2(new_n615), .ZN(G284));
  AOI21_X1  g191(.A(new_n599), .B1(new_n597), .B2(new_n615), .ZN(G321));
  NOR2_X1   g192(.A1(G168), .A2(new_n614), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(KEYINPUT83), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n619), .A2(KEYINPUT83), .ZN(new_n621));
  NAND2_X1  g196(.A1(G299), .A2(new_n614), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(G297));
  AOI21_X1  g198(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(G280));
  INV_X1    g199(.A(new_n613), .ZN(new_n625));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n551), .A2(new_n614), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n613), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n467), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n461), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  AND3_X1   g209(.A1(new_n475), .A2(KEYINPUT84), .A3(G123), .ZN(new_n635));
  AOI21_X1  g210(.A(KEYINPUT84), .B1(new_n475), .B2(G123), .ZN(new_n636));
  OAI221_X1 g211(.A(new_n632), .B1(new_n633), .B2(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND3_X1  g213(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n638), .A2(new_n642), .ZN(G156));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AND2_X1   g234(.A1(new_n659), .A2(KEYINPUT86), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(KEYINPUT86), .B2(new_n659), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n661), .C2(new_n662), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n659), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT88), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n681), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n682), .A2(KEYINPUT89), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(KEYINPUT89), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n690), .A2(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(KEYINPUT20), .ZN(new_n692));
  OAI221_X1 g267(.A(new_n687), .B1(new_n686), .B2(new_n681), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT90), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n695), .A2(G1986), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n699), .B1(new_n696), .B2(new_n700), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n677), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n703), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n705), .A2(new_n676), .A3(new_n701), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G4), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n625), .B2(new_n709), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT96), .B(G1348), .Z(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G26), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT97), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n467), .A2(G140), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n475), .A2(G128), .ZN(new_n719));
  OR2_X1    g294(.A1(G104), .A2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n720), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n717), .B1(new_n723), .B2(new_n714), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2067), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT92), .B(G16), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(G19), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n552), .B2(new_n726), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1341), .ZN(new_n729));
  NOR3_X1   g304(.A1(new_n713), .A2(new_n725), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT98), .ZN(new_n731));
  NOR2_X1   g306(.A1(G168), .A2(new_n709), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n709), .B2(G21), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G1961), .ZN(new_n736));
  NOR2_X1   g311(.A1(G171), .A2(new_n709), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G5), .B2(new_n709), .ZN(new_n738));
  OAI22_X1  g313(.A1(new_n733), .A2(new_n734), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n735), .B(new_n739), .C1(new_n736), .C2(new_n738), .ZN(new_n740));
  INV_X1    g315(.A(G20), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n726), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT23), .Z(new_n743));
  AND2_X1   g318(.A1(new_n566), .A2(new_n571), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n709), .ZN(new_n745));
  INV_X1    g320(.A(G1956), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G35), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G162), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT29), .B(G2090), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n714), .A2(G33), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT25), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n471), .A2(G127), .ZN(new_n755));
  NAND2_X1  g330(.A1(G115), .A2(G2104), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n461), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n754), .B(new_n757), .C1(G139), .C2(new_n467), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(new_n714), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G2072), .Z(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT31), .B(G11), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n762), .A2(G28), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n714), .B1(new_n762), .B2(G28), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n761), .B1(new_n763), .B2(new_n764), .C1(new_n637), .C2(new_n714), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n714), .A2(G32), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n467), .A2(G141), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n475), .A2(G129), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT26), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  INV_X1    g347(.A(G2104), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G2105), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n771), .A2(new_n772), .B1(G105), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n767), .A2(new_n768), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n766), .B1(new_n777), .B2(new_n714), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT27), .B(G1996), .Z(new_n779));
  AOI21_X1  g354(.A(new_n765), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  INV_X1    g356(.A(G34), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n782), .A2(KEYINPUT24), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(KEYINPUT24), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n714), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G160), .B2(new_n714), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT99), .B(G2084), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n760), .A2(new_n780), .A3(new_n781), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G27), .A2(G29), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G164), .B2(G29), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2078), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n751), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n731), .A2(new_n740), .A3(new_n747), .A4(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n795));
  MUX2_X1   g370(.A(G6), .B(G305), .S(G16), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1981), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n726), .A2(G22), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G166), .B2(new_n726), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(G1971), .Z(new_n801));
  AND2_X1   g376(.A1(new_n709), .A2(G23), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G288), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT33), .B(G1976), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n801), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT34), .B1(new_n798), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT95), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n798), .A2(KEYINPUT34), .A3(new_n807), .ZN(new_n810));
  XNOR2_X1  g385(.A(G290), .B(KEYINPUT93), .ZN(new_n811));
  MUX2_X1   g386(.A(G24), .B(new_n811), .S(new_n726), .Z(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT94), .B(G1986), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n467), .A2(G131), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT91), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(G107), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G2105), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n475), .B2(G119), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  MUX2_X1   g396(.A(G25), .B(new_n821), .S(G29), .Z(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XOR2_X1   g398(.A(new_n822), .B(new_n823), .Z(new_n824));
  AND2_X1   g399(.A1(new_n812), .A2(new_n813), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n810), .A2(new_n814), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n795), .B1(new_n809), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n809), .A2(new_n826), .A3(new_n795), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n794), .B1(new_n828), .B2(new_n829), .ZN(G311));
  INV_X1    g405(.A(new_n794), .ZN(new_n831));
  INV_X1    g406(.A(new_n829), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n827), .ZN(G150));
  XOR2_X1   g408(.A(KEYINPUT102), .B(G860), .Z(new_n834));
  AOI22_X1  g409(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(new_n509), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n524), .A2(G93), .B1(G55), .B2(new_n515), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n613), .A2(new_n626), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n836), .A2(new_n837), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n551), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n548), .A2(new_n836), .A3(new_n550), .A4(new_n837), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n843), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT101), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n834), .B1(new_n848), .B2(new_n849), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n840), .B1(new_n851), .B2(new_n852), .ZN(G145));
  XNOR2_X1  g428(.A(new_n821), .B(new_n640), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n758), .B(new_n777), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(G164), .B(new_n723), .ZN(new_n857));
  AOI22_X1  g432(.A1(G130), .A2(new_n475), .B1(new_n467), .B2(G142), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n860));
  INV_X1    g435(.A(G118), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n859), .A2(new_n860), .B1(new_n861), .B2(G2105), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n860), .B2(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n857), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n856), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G160), .ZN(new_n867));
  XNOR2_X1  g442(.A(G162), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n637), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n866), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT105), .B(G37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(KEYINPUT106), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n870), .B2(new_n871), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(G395));
  NAND2_X1  g453(.A1(new_n844), .A2(new_n614), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n847), .B(new_n629), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n566), .A2(new_n571), .A3(new_n607), .A4(new_n612), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n566), .A2(new_n571), .B1(new_n607), .B2(new_n612), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT107), .Z(new_n886));
  XNOR2_X1  g461(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n882), .B2(new_n883), .ZN(new_n889));
  NAND2_X1  g464(.A1(G299), .A2(new_n613), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n891), .A3(new_n881), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n880), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G288), .B(G305), .ZN(new_n895));
  XOR2_X1   g470(.A(G166), .B(G290), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT42), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n894), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n879), .B1(new_n899), .B2(new_n614), .ZN(G295));
  OAI21_X1  g475(.A(new_n879), .B1(new_n899), .B2(new_n614), .ZN(G331));
  OAI21_X1  g476(.A(G168), .B1(new_n576), .B2(new_n577), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n845), .A2(new_n846), .ZN(new_n903));
  OAI21_X1  g478(.A(G64), .B1(new_n601), .B2(new_n603), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n539), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT76), .B1(new_n905), .B2(G651), .ZN(new_n906));
  INV_X1    g481(.A(new_n545), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n575), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(G286), .A2(new_n908), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n902), .A2(new_n903), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n903), .B1(new_n902), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n884), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(KEYINPUT79), .ZN(new_n913));
  NAND2_X1  g488(.A1(G171), .A2(new_n573), .ZN(new_n914));
  AOI21_X1  g489(.A(G286), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n909), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n847), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n889), .A2(new_n892), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n902), .A2(new_n903), .A3(new_n909), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n912), .A2(new_n897), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n897), .B1(new_n912), .B2(new_n920), .ZN(new_n924));
  OR3_X1    g499(.A1(new_n923), .A2(KEYINPUT43), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n897), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n890), .A2(new_n881), .A3(new_n887), .ZN(new_n927));
  OAI211_X1 g502(.A(KEYINPUT110), .B(new_n927), .C1(new_n884), .C2(new_n891), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n884), .A2(new_n929), .A3(new_n887), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n928), .A2(new_n917), .A3(new_n919), .A4(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n884), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n917), .B2(new_n919), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n912), .A2(KEYINPUT111), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n926), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n921), .A2(new_n871), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  OAI211_X1 g515(.A(KEYINPUT44), .B(new_n925), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT43), .B1(new_n923), .B2(new_n924), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT109), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n944), .B(KEYINPUT43), .C1(new_n923), .C2(new_n924), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n940), .A3(new_n938), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n948), .B1(new_n947), .B2(new_n949), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n941), .B1(new_n950), .B2(new_n951), .ZN(G397));
  NAND2_X1  g527(.A1(new_n492), .A2(new_n494), .ZN(new_n953));
  AOI21_X1  g528(.A(G1384), .B1(new_n953), .B2(new_n485), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n955));
  AND2_X1   g530(.A1(G160), .A2(G40), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G164), .B2(G1384), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(G2078), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n960), .A2(KEYINPUT53), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n956), .A3(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n960), .A2(KEYINPUT53), .B1(new_n736), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(new_n966), .A3(G301), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n961), .A2(new_n966), .ZN(new_n968));
  OAI211_X1 g543(.A(KEYINPUT54), .B(new_n967), .C1(new_n968), .C2(new_n908), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT54), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n961), .A2(new_n966), .A3(G301), .ZN(new_n971));
  AOI21_X1  g546(.A(G301), .B1(new_n961), .B2(new_n966), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT126), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(KEYINPUT51), .ZN(new_n975));
  INV_X1    g550(.A(G8), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n964), .A2(new_n956), .ZN(new_n977));
  INV_X1    g552(.A(G2084), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n978), .A3(new_n963), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n959), .A2(new_n734), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI22_X1  g556(.A1(G286), .A2(G8), .B1(new_n974), .B2(KEYINPUT51), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n975), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n975), .ZN(new_n985));
  INV_X1    g560(.A(new_n965), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n986), .A2(new_n978), .B1(new_n959), .B2(new_n734), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n982), .B(new_n985), .C1(new_n987), .C2(new_n976), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n979), .A2(new_n980), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(G8), .A3(G286), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n984), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n969), .A2(new_n973), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n585), .A2(G1976), .A3(new_n586), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n956), .A2(new_n954), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G8), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT116), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n998), .A3(G8), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n994), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(G288), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(G305), .A2(G1981), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n591), .A2(new_n694), .A3(new_n592), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1003), .A2(new_n1007), .A3(new_n1004), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n997), .A2(new_n999), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1000), .A2(new_n1002), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT117), .B1(new_n1000), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G303), .A2(G8), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT115), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OR4_X1    g591(.A1(KEYINPUT115), .A2(G166), .A3(new_n1015), .A4(new_n976), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G2090), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n977), .A2(new_n1020), .A3(new_n963), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT114), .B(G1971), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n959), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n976), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n999), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n998), .B1(new_n995), .B2(G8), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n993), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(KEYINPUT52), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1011), .A2(new_n1013), .A3(new_n1025), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1019), .ZN(new_n1033));
  AOI21_X1  g608(.A(G2090), .B1(new_n965), .B2(KEYINPUT118), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n977), .A2(new_n1035), .A3(new_n963), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1023), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(KEYINPUT119), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1034), .A2(new_n1036), .B1(new_n959), .B2(new_n1022), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1033), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1032), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n992), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n995), .ZN(new_n1046));
  INV_X1    g621(.A(G2067), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n965), .A2(new_n712), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT60), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n625), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1048), .B(new_n625), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n1049), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n965), .A2(new_n746), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n568), .A2(new_n570), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT122), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n524), .B2(G91), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1054), .A2(KEYINPUT122), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI22_X1  g634(.A1(G299), .A2(KEYINPUT57), .B1(new_n1059), .B2(new_n566), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n955), .A2(new_n958), .A3(new_n956), .A4(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1053), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT61), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1060), .B1(new_n1053), .B2(new_n1062), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1059), .A2(new_n566), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(new_n744), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1956), .B1(new_n977), .B2(new_n963), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1062), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT61), .B1(new_n1073), .B2(new_n1063), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1067), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n1076));
  INV_X1    g651(.A(G1996), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n955), .A2(new_n958), .A3(new_n1077), .A4(new_n956), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(G1341), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n995), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n551), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1076), .B1(new_n1082), .B2(KEYINPUT124), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(KEYINPUT124), .B2(new_n1082), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1082), .A2(KEYINPUT124), .A3(KEYINPUT59), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1075), .A2(KEYINPUT125), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1065), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1073), .A2(KEYINPUT61), .A3(new_n1063), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1084), .A2(new_n1087), .A3(new_n1085), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1052), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1048), .A2(new_n613), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1073), .B1(new_n1093), .B2(new_n1064), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1045), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n984), .A2(new_n988), .A3(new_n1097), .A4(new_n990), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n972), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT127), .B1(new_n1099), .B2(new_n1044), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1098), .A2(new_n972), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1038), .A2(KEYINPUT119), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(G8), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1031), .B1(new_n1104), .B2(new_n1033), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT127), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1101), .A2(new_n1105), .A3(new_n1106), .A4(new_n1096), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g683(.A(G1976), .B(G288), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1004), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1010), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1011), .A2(new_n1030), .A3(new_n1013), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n1025), .B2(new_n1112), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n987), .A2(new_n976), .A3(G286), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1032), .A2(new_n1043), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1011), .A2(new_n1030), .A3(new_n1013), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1019), .B1(new_n1024), .B2(KEYINPUT120), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(KEYINPUT120), .B2(new_n1024), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1024), .A2(KEYINPUT120), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1124), .B(new_n976), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1123), .A2(new_n1125), .A3(new_n1019), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT121), .B1(new_n1126), .B2(new_n1112), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1114), .A2(KEYINPUT63), .A3(new_n1025), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1122), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1113), .B1(new_n1117), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1095), .A2(new_n1108), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(G160), .A2(G40), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n954), .A2(KEYINPUT45), .A3(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n722), .B(new_n1047), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT113), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1133), .B1(new_n1136), .B2(new_n776), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1077), .B2(new_n1135), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1133), .A2(new_n1077), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1138), .B1(new_n777), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1133), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n821), .B(new_n823), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(G290), .B(G1986), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1133), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1131), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1141), .A2(new_n823), .A3(new_n816), .A4(new_n820), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n723), .A2(new_n1047), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1142), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1139), .B(KEYINPUT46), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1137), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT47), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1142), .A2(G1986), .A3(G290), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT48), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1144), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1147), .A2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  XNOR2_X1  g733(.A(new_n872), .B(KEYINPUT106), .ZN(new_n1160));
  NOR3_X1   g734(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1161));
  NAND4_X1  g735(.A1(new_n1160), .A2(new_n707), .A3(new_n947), .A4(new_n1161), .ZN(G225));
  INV_X1    g736(.A(G225), .ZN(G308));
endmodule


