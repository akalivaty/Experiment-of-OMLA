//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n204));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT2), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT81), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT81), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(new_n205), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n211), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n212), .A2(new_n213), .ZN(new_n221));
  AND2_X1   g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n221), .A2(new_n224), .A3(new_n218), .A4(new_n206), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n220), .A2(new_n225), .A3(KEYINPUT3), .ZN(new_n226));
  XNOR2_X1  g025(.A(G211gat), .B(G218gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G197gat), .B(G204gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT78), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n230), .A2(KEYINPUT78), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n228), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n233), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n235), .A2(new_n227), .A3(new_n231), .A4(new_n229), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT79), .B(KEYINPUT29), .Z(new_n238));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n225), .A3(new_n238), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n204), .B(new_n226), .C1(new_n237), .C2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n236), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n220), .A2(new_n225), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(new_n238), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n204), .B1(new_n244), .B2(new_n226), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT3), .B1(new_n220), .B2(new_n225), .ZN(new_n247));
  INV_X1    g046(.A(new_n238), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT87), .B1(new_n249), .B2(new_n242), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n220), .A2(new_n225), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n238), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT87), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n255), .A3(new_n237), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n203), .B1(new_n246), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n252), .B1(new_n237), .B2(KEYINPUT29), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n202), .B1(new_n259), .B2(new_n243), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT88), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n249), .A2(KEYINPUT88), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n237), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(G22gat), .B1(new_n258), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n226), .B1(new_n237), .B2(new_n239), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT86), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n269), .A2(new_n256), .A3(new_n250), .A4(new_n240), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n270), .A2(new_n202), .B1(new_n264), .B2(new_n260), .ZN(new_n271));
  INV_X1    g070(.A(G22gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT89), .ZN(new_n274));
  XOR2_X1   g073(.A(G78gat), .B(G106gat), .Z(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT85), .B(G50gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n267), .A2(new_n273), .A3(new_n274), .A4(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT89), .B1(new_n271), .B2(new_n272), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n282), .A2(new_n279), .B1(new_n267), .B2(new_n273), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT77), .B(KEYINPUT34), .Z(new_n285));
  INV_X1    g084(.A(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G113gat), .ZN(new_n287));
  INV_X1    g086(.A(G113gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G120gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(KEYINPUT74), .A2(KEYINPUT1), .ZN(new_n291));
  NOR2_X1   g090(.A1(KEYINPUT74), .A2(KEYINPUT1), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G127gat), .B(G134gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G127gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G134gat), .ZN(new_n297));
  INV_X1    g096(.A(G134gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G127gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n296), .A2(KEYINPUT73), .A3(G134gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT1), .B1(new_n287), .B2(new_n289), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n295), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n308));
  XNOR2_X1  g107(.A(G113gat), .B(G120gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n301), .B(new_n302), .C1(KEYINPUT1), .C2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(KEYINPUT75), .A3(new_n295), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n313));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT26), .ZN(new_n315));
  INV_X1    g114(.A(G169gat), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  AND4_X1   g116(.A1(KEYINPUT71), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT71), .B1(new_n319), .B2(new_n315), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n322), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n314), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT70), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT27), .B(G183gat), .ZN(new_n331));
  INV_X1    g130(.A(G190gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G183gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT27), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G183gat), .ZN(new_n337));
  AND4_X1   g136(.A1(new_n332), .A2(new_n335), .A3(new_n337), .A4(new_n330), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n313), .B1(new_n328), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n337), .A3(new_n332), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(KEYINPUT70), .A3(new_n329), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n331), .A2(new_n332), .A3(new_n330), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n323), .A2(G169gat), .A3(G176gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n347), .B(new_n322), .C1(new_n318), .C2(new_n320), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n344), .A2(KEYINPUT72), .A3(new_n314), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n340), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n314), .ZN(new_n352));
  NAND3_X1  g151(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(G176gat), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n357), .B2(new_n316), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  OAI22_X1  g158(.A1(KEYINPUT67), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI22_X1  g161(.A1(new_n324), .A2(new_n326), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT69), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n360), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n365), .A2(new_n361), .B1(new_n345), .B2(new_n346), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT69), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n354), .A4(new_n358), .ZN(new_n368));
  AND2_X1   g167(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(KEYINPUT65), .A3(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n352), .A3(new_n372), .ZN(new_n373));
  OR2_X1    g172(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n366), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n378));
  AOI22_X1  g177(.A1(new_n364), .A2(new_n368), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n312), .B1(new_n350), .B2(new_n379), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n307), .A2(new_n308), .A3(new_n311), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n308), .B1(new_n307), .B2(new_n311), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n376), .B(new_n347), .C1(new_n362), .C2(new_n360), .ZN(new_n384));
  INV_X1    g183(.A(new_n373), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n378), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n314), .A2(new_n351), .B1(new_n369), .B2(G190gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT23), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT25), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n367), .B1(new_n390), .B2(new_n366), .ZN(new_n391));
  NOR4_X1   g190(.A1(new_n363), .A2(new_n387), .A3(KEYINPUT69), .A4(new_n389), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n386), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n340), .A3(new_n349), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n380), .B1(new_n383), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G227gat), .ZN(new_n396));
  INV_X1    g195(.A(G233gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT33), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G15gat), .B(G43gat), .Z(new_n400));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n285), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n285), .ZN(new_n405));
  INV_X1    g204(.A(new_n398), .ZN(new_n406));
  INV_X1    g205(.A(new_n350), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n407), .B(new_n393), .C1(new_n382), .C2(new_n381), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n408), .B2(new_n380), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n405), .B(new_n402), .C1(new_n409), .C2(KEYINPUT33), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n398), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(new_n406), .A3(new_n380), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT32), .ZN(new_n414));
  OR3_X1    g213(.A1(new_n395), .A2(KEYINPUT32), .A3(new_n398), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n404), .A2(new_n410), .A3(new_n415), .A4(new_n414), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  XOR2_X1   g219(.A(G1gat), .B(G29gat), .Z(new_n421));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT5), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n243), .A2(new_n305), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n251), .A2(new_n310), .A3(new_n295), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n426), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n243), .A2(KEYINPUT4), .A3(new_n305), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n307), .A2(new_n251), .A3(new_n311), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(KEYINPUT4), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n226), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n220), .A2(new_n225), .A3(KEYINPUT82), .A4(KEYINPUT3), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n437), .A2(new_n253), .A3(new_n438), .A4(new_n305), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n430), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n432), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n243), .A2(new_n442), .A3(new_n305), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n442), .B2(new_n434), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n444), .A2(new_n426), .A3(new_n430), .A4(new_n439), .ZN(new_n445));
  AOI211_X1 g244(.A(new_n420), .B(new_n425), .C1(new_n441), .C2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(new_n445), .A3(new_n425), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n447), .A2(new_n420), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n445), .ZN(new_n449));
  INV_X1    g248(.A(new_n425), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n446), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G226gat), .A2(G233gat), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n248), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n350), .B2(new_n379), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n328), .A2(new_n339), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n393), .A2(new_n459), .A3(new_n455), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n457), .A2(new_n237), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n393), .A2(new_n455), .A3(new_n340), .A4(new_n349), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n455), .A2(KEYINPUT29), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n379), .B2(new_n458), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n237), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT80), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n464), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n242), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n457), .A2(new_n237), .A3(new_n460), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G8gat), .B(G36gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G64gat), .B(G92gat), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n472), .B(new_n473), .Z(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n466), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n468), .A2(new_n469), .A3(new_n474), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n379), .A2(new_n458), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n394), .A2(new_n456), .B1(new_n480), .B2(new_n455), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n465), .B1(new_n237), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(KEYINPUT30), .A3(new_n474), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n476), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n284), .A2(new_n419), .A3(new_n453), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n270), .A2(new_n202), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n272), .B1(new_n487), .B2(new_n265), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n279), .B1(new_n488), .B2(new_n274), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n267), .A2(new_n273), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n280), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(new_n418), .B2(new_n417), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT90), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n425), .B(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n441), .B2(new_n445), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n446), .B1(new_n448), .B2(new_n497), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n484), .A2(new_n498), .A3(KEYINPUT35), .ZN(new_n499));
  AOI22_X1  g298(.A1(KEYINPUT35), .A2(new_n486), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  INV_X1    g300(.A(new_n418), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n404), .A2(new_n410), .B1(new_n415), .B2(new_n414), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI22_X1  g303(.A1(new_n281), .A2(new_n283), .B1(new_n484), .B2(new_n452), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n417), .A2(KEYINPUT36), .A3(new_n418), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT39), .B1(new_n429), .B2(new_n431), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n434), .A2(new_n442), .ZN(new_n509));
  INV_X1    g308(.A(new_n443), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n439), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n508), .B1(new_n511), .B2(new_n431), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT39), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n514), .A3(new_n431), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n513), .A2(KEYINPUT40), .A3(new_n495), .A4(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT40), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n495), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n512), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n484), .A2(new_n497), .A3(new_n516), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n449), .A2(KEYINPUT6), .A3(new_n450), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n447), .A2(new_n420), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n521), .B(new_n477), .C1(new_n522), .C2(new_n496), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n237), .B1(new_n457), .B2(new_n460), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n526));
  OAI22_X1  g325(.A1(new_n525), .A2(new_n526), .B1(new_n467), .B2(new_n242), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n481), .A2(KEYINPUT91), .A3(new_n237), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT37), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT38), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n474), .B1(new_n482), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n466), .A2(KEYINPUT37), .A3(new_n471), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n530), .B1(new_n534), .B2(new_n532), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n524), .B(new_n533), .C1(new_n535), .C2(KEYINPUT92), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  AOI211_X1 g336(.A(new_n537), .B(new_n530), .C1(new_n534), .C2(new_n532), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n284), .B(new_n520), .C1(new_n536), .C2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n507), .B1(new_n539), .B2(KEYINPUT93), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n534), .A2(new_n532), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT38), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n537), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n535), .A2(KEYINPUT92), .ZN(new_n544));
  AOI211_X1 g343(.A(KEYINPUT38), .B(new_n474), .C1(new_n482), .C2(new_n531), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n523), .B1(new_n529), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n519), .A2(new_n516), .A3(new_n497), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n477), .B(KEYINPUT30), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n476), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(new_n492), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n500), .B1(new_n540), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G43gat), .B(G50gat), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(G29gat), .B2(G36gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(G29gat), .A2(G36gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT14), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n557), .B(new_n560), .C1(KEYINPUT15), .C2(new_n555), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(KEYINPUT95), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n563));
  INV_X1    g362(.A(G29gat), .ZN(new_n564));
  INV_X1    g363(.A(G36gat), .ZN(new_n565));
  OAI22_X1  g364(.A1(new_n559), .A2(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n556), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT17), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G1gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT16), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n572), .A3(G1gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G8gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n571), .A2(G1gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(KEYINPUT97), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n579), .B(new_n582), .Z(new_n583));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n569), .A2(new_n583), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT18), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592));
  INV_X1    g391(.A(G197gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT11), .B(G169gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT12), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n586), .A2(KEYINPUT18), .A3(new_n587), .A4(new_n588), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n569), .B(new_n583), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n587), .B(KEYINPUT13), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n591), .A2(new_n597), .A3(new_n598), .A4(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n589), .A2(new_n590), .B1(new_n599), .B2(new_n600), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n605), .A2(KEYINPUT98), .A3(new_n597), .A4(new_n598), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n598), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n597), .B(KEYINPUT94), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G57gat), .B(G64gat), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g414(.A1(KEYINPUT99), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(G71gat), .B2(G78gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n615), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n618), .A2(new_n619), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT21), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G127gat), .ZN(new_n628));
  XOR2_X1   g427(.A(G183gat), .B(G211gat), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n628), .A2(new_n630), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n583), .B1(new_n623), .B2(new_n624), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(new_n215), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n635), .B(new_n637), .Z(new_n638));
  OR3_X1    g437(.A1(new_n631), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n631), .B2(new_n632), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G85gat), .A2(G92gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT7), .ZN(new_n643));
  NAND2_X1  g442(.A1(G99gat), .A2(G106gat), .ZN(new_n644));
  INV_X1    g443(.A(G85gat), .ZN(new_n645));
  INV_X1    g444(.A(G92gat), .ZN(new_n646));
  AOI22_X1  g445(.A1(KEYINPUT8), .A2(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G99gat), .B(G106gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(G232gat), .A2(G233gat), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n568), .A2(new_n651), .B1(KEYINPUT41), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n585), .A2(new_n650), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n568), .A2(new_n584), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G190gat), .B(G218gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT104), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n652), .A2(KEYINPUT41), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT103), .ZN(new_n662));
  XNOR2_X1  g461(.A(G134gat), .B(G162gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n658), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n666), .B(new_n653), .C1(new_n654), .C2(new_n655), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n660), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n664), .B1(new_n659), .B2(new_n667), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT10), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n650), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n672), .B1(new_n623), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n615), .B(new_n617), .Z(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT100), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n620), .A3(new_n650), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n649), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n648), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n677), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n679), .A2(new_n673), .A3(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n674), .B(KEYINPUT106), .C1(new_n621), .C2(new_n622), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n676), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(G230gat), .A2(G233gat), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(G120gat), .B(G148gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(G176gat), .B(G204gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(new_n691));
  NAND2_X1  g490(.A1(new_n679), .A2(new_n683), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693));
  INV_X1    g492(.A(new_n687), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT107), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n688), .A2(new_n691), .A3(new_n695), .A4(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n698), .B2(new_n699), .ZN(new_n703));
  INV_X1    g502(.A(new_n691), .ZN(new_n704));
  INV_X1    g503(.A(new_n688), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n697), .A2(new_n695), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n702), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n707), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n698), .A2(new_n699), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT109), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(new_n701), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n641), .A2(new_n671), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n554), .A2(new_n612), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n452), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n484), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT110), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n715), .A2(new_n720), .A3(new_n484), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT16), .B(G8gat), .Z(new_n723));
  AOI21_X1  g522(.A(KEYINPUT42), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n719), .A2(G8gat), .A3(new_n721), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n715), .A2(KEYINPUT42), .A3(new_n484), .A4(new_n723), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n724), .A2(new_n727), .A3(KEYINPUT111), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT111), .B1(new_n724), .B2(new_n727), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1325gat));
  INV_X1    g529(.A(new_n715), .ZN(new_n731));
  INV_X1    g530(.A(new_n504), .ZN(new_n732));
  INV_X1    g531(.A(new_n506), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G15gat), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n554), .A2(new_n612), .ZN(new_n736));
  INV_X1    g535(.A(new_n419), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n714), .A2(G15gat), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(G1326gat));
  NAND2_X1  g539(.A1(new_n715), .A2(new_n492), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT43), .B(G22gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1327gat));
  INV_X1    g542(.A(new_n641), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n713), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n671), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n736), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n747), .A2(G29gat), .A3(new_n453), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n745), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n611), .ZN(new_n752));
  INV_X1    g551(.A(new_n671), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n548), .B1(new_n547), .B2(new_n552), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n754), .A2(new_n755), .A3(new_n507), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n753), .B1(new_n756), .B2(new_n500), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(KEYINPUT113), .A3(KEYINPUT44), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n539), .A2(KEYINPUT93), .ZN(new_n760));
  INV_X1    g559(.A(new_n507), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(new_n553), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n500), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n671), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n759), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n756), .B2(new_n500), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n554), .A2(KEYINPUT114), .ZN(new_n770));
  INV_X1    g569(.A(new_n669), .ZN(new_n771));
  INV_X1    g570(.A(new_n670), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(KEYINPUT115), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n669), .B2(new_n670), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n769), .A2(new_n770), .A3(new_n765), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n752), .B1(new_n767), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(new_n452), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n750), .B1(new_n779), .B2(new_n564), .ZN(G1328gat));
  NOR3_X1   g579(.A1(new_n747), .A2(G36gat), .A3(new_n485), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT46), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n778), .A2(new_n484), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n565), .ZN(G1329gat));
  NOR3_X1   g583(.A1(new_n747), .A2(G43gat), .A3(new_n737), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n734), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n778), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(G43gat), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT47), .B(new_n786), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n778), .B2(new_n787), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n785), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(G1330gat));
  INV_X1    g593(.A(KEYINPUT48), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT113), .B1(new_n757), .B2(KEYINPUT44), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n764), .A2(new_n759), .A3(new_n765), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n777), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n798), .A2(new_n492), .A3(new_n611), .A4(new_n751), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G50gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n747), .A2(G50gat), .A3(new_n284), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n795), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  AOI211_X1 g602(.A(KEYINPUT48), .B(new_n801), .C1(new_n799), .C2(G50gat), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(G1331gat));
  AND2_X1   g604(.A1(new_n769), .A2(new_n770), .ZN(new_n806));
  NOR4_X1   g605(.A1(new_n744), .A2(new_n611), .A3(new_n753), .A4(new_n713), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n452), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g609(.A(new_n485), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT116), .ZN(new_n813));
  NOR2_X1   g612(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n808), .A2(new_n815), .A3(new_n811), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n814), .B1(new_n813), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(G1333gat));
  NAND2_X1  g618(.A1(new_n806), .A2(new_n807), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n419), .B(KEYINPUT117), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n787), .A2(G71gat), .ZN(new_n824));
  OAI22_X1  g623(.A1(new_n823), .A2(G71gat), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g625(.A1(new_n820), .A2(new_n284), .ZN(new_n827));
  XOR2_X1   g626(.A(KEYINPUT118), .B(G78gat), .Z(new_n828));
  XNOR2_X1  g627(.A(new_n827), .B(new_n828), .ZN(G1335gat));
  INV_X1    g628(.A(new_n713), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n639), .A2(new_n640), .A3(new_n612), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT51), .B1(new_n764), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n834));
  NOR4_X1   g633(.A1(new_n554), .A2(new_n834), .A3(new_n671), .A4(new_n831), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n830), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n645), .A3(new_n452), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n831), .A2(new_n713), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n767), .B2(new_n777), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n452), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n838), .B1(new_n842), .B2(new_n645), .ZN(G1336gat));
  NOR3_X1   g642(.A1(new_n836), .A2(G92gat), .A3(new_n485), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n841), .A2(new_n484), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n845), .B(new_n846), .C1(new_n847), .C2(new_n646), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n646), .B1(new_n841), .B2(new_n484), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT52), .B1(new_n849), .B2(new_n844), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1337gat));
  INV_X1    g650(.A(G99gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n852), .A3(new_n419), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n841), .A2(new_n787), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n852), .ZN(G1338gat));
  INV_X1    g654(.A(G106gat), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n841), .B2(new_n492), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n833), .A2(new_n835), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n713), .A2(G106gat), .A3(new_n284), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT119), .Z(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT53), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n798), .A2(new_n492), .A3(new_n839), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G106gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n859), .B1(new_n833), .B2(new_n835), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT120), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870));
  AOI211_X1 g669(.A(new_n870), .B(new_n867), .C1(new_n863), .C2(G106gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n862), .B1(new_n869), .B2(new_n871), .ZN(G1339gat));
  NAND4_X1  g671(.A1(new_n641), .A2(new_n612), .A3(new_n671), .A4(new_n713), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n688), .A2(KEYINPUT54), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n676), .A2(new_n684), .A3(new_n694), .A4(new_n685), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n688), .A2(KEYINPUT54), .A3(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n874), .A2(KEYINPUT55), .A3(new_n704), .A4(new_n876), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n698), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n586), .A2(new_n588), .ZN(new_n879));
  OAI22_X1  g678(.A1(new_n879), .A2(new_n587), .B1(new_n599), .B2(new_n600), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n604), .A2(new_n606), .B1(new_n596), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n874), .A2(new_n704), .A3(new_n876), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND4_X1   g683(.A1(new_n776), .A2(new_n878), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n708), .B2(new_n712), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n611), .A2(new_n884), .A3(new_n878), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n776), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n873), .B1(new_n890), .B2(new_n641), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n453), .A2(new_n484), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n891), .A2(new_n284), .A3(new_n419), .A4(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(new_n288), .A3(new_n612), .ZN(new_n894));
  INV_X1    g693(.A(new_n891), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n453), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n493), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n485), .A3(new_n611), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n894), .B1(new_n899), .B2(new_n288), .ZN(G1340gat));
  NOR3_X1   g699(.A1(new_n893), .A2(new_n286), .A3(new_n713), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n485), .A3(new_n830), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n286), .ZN(G1341gat));
  OAI21_X1  g702(.A(G127gat), .B1(new_n893), .B2(new_n744), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n898), .A2(new_n485), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n641), .A2(new_n296), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(G1342gat));
  NAND2_X1  g706(.A1(new_n753), .A2(new_n485), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(G134gat), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  OR3_X1    g709(.A1(new_n897), .A2(KEYINPUT56), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G134gat), .B1(new_n893), .B2(new_n671), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT56), .B1(new_n897), .B2(new_n910), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(G1343gat));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n734), .A2(new_n892), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT57), .B1(new_n891), .B2(new_n492), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT57), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n284), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n753), .B1(new_n886), .B2(new_n887), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n744), .B1(new_n921), .B2(new_n885), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n922), .B2(new_n873), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n611), .B(new_n916), .C1(new_n917), .C2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n915), .B1(new_n924), .B2(G141gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n787), .A2(new_n284), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n891), .A2(new_n452), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n611), .A2(new_n207), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n927), .A2(new_n484), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n929), .B1(new_n924), .B2(G141gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n925), .A2(new_n930), .A3(KEYINPUT58), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT58), .ZN(new_n932));
  AOI221_X4 g731(.A(new_n929), .B1(new_n915), .B2(new_n932), .C1(G141gat), .C2(new_n924), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n931), .A2(new_n933), .ZN(G1344gat));
  NAND2_X1  g733(.A1(new_n888), .A2(new_n671), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n878), .A2(new_n881), .A3(new_n753), .A4(new_n884), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n641), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n873), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n492), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n918), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n891), .A2(new_n919), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n830), .A3(new_n916), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n927), .A2(new_n484), .A3(new_n713), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n208), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n917), .A2(new_n923), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n948), .A2(new_n946), .A3(new_n830), .A4(new_n916), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n944), .A2(new_n947), .A3(new_n949), .ZN(G1345gat));
  AND2_X1   g749(.A1(new_n948), .A2(new_n916), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n641), .A2(G155gat), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT122), .ZN(new_n953));
  OR3_X1    g752(.A1(new_n927), .A2(new_n484), .A3(new_n744), .ZN(new_n954));
  AOI22_X1  g753(.A1(new_n951), .A2(new_n953), .B1(new_n215), .B2(new_n954), .ZN(G1346gat));
  OR3_X1    g754(.A1(new_n927), .A2(G162gat), .A3(new_n908), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n951), .A2(new_n776), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n216), .ZN(G1347gat));
  NOR2_X1   g757(.A1(new_n485), .A2(new_n452), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n822), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n891), .A2(new_n284), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(G169gat), .B1(new_n962), .B2(new_n612), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n895), .A2(new_n452), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n737), .A2(new_n485), .A3(new_n492), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n611), .A2(new_n374), .A3(new_n375), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(G1348gat));
  INV_X1    g767(.A(new_n966), .ZN(new_n969));
  AOI21_X1  g768(.A(G176gat), .B1(new_n969), .B2(new_n830), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n962), .A2(new_n317), .A3(new_n713), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(KEYINPUT123), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(KEYINPUT123), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(G1349gat));
  NAND4_X1  g773(.A1(new_n964), .A2(new_n331), .A3(new_n641), .A4(new_n965), .ZN(new_n975));
  OAI21_X1  g774(.A(G183gat), .B1(new_n962), .B2(new_n744), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT60), .ZN(new_n977));
  AOI22_X1  g776(.A1(new_n975), .A2(new_n976), .B1(KEYINPUT124), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n978), .B(new_n979), .ZN(G1350gat));
  OAI21_X1  g779(.A(G190gat), .B1(new_n962), .B2(new_n671), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT61), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n969), .A2(new_n332), .A3(new_n776), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1351gat));
  NAND2_X1  g783(.A1(new_n926), .A2(new_n484), .ZN(new_n985));
  XOR2_X1   g784(.A(new_n985), .B(KEYINPUT125), .Z(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(new_n964), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(G197gat), .B1(new_n988), .B2(new_n611), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n787), .A2(new_n960), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n991), .B1(new_n940), .B2(new_n941), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n612), .A2(new_n593), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(G1352gat));
  NOR2_X1   g793(.A1(new_n713), .A2(G204gat), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n986), .A2(new_n964), .A3(new_n995), .ZN(new_n996));
  XOR2_X1   g795(.A(new_n996), .B(KEYINPUT62), .Z(new_n997));
  NAND2_X1  g796(.A1(new_n992), .A2(new_n830), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT126), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(G204gat), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n998), .A2(new_n999), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n997), .B1(new_n1001), .B2(new_n1002), .ZN(G1353gat));
  OR3_X1    g802(.A1(new_n987), .A2(G211gat), .A3(new_n744), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n992), .A2(new_n641), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  AOI21_X1  g807(.A(G218gat), .B1(new_n988), .B2(new_n776), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n753), .A2(G218gat), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1010), .B(KEYINPUT127), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n1009), .B1(new_n992), .B2(new_n1011), .ZN(G1355gat));
endmodule


