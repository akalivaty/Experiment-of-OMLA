//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203));
  AND2_X1   g002(.A1(G113gat), .A2(G120gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G113gat), .A2(G120gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G127gat), .ZN(new_n210));
  INV_X1    g009(.A(G127gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G134gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n208), .A2(new_n210), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G113gat), .B(G120gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT73), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(KEYINPUT72), .B(KEYINPUT1), .Z(new_n217));
  INV_X1    g016(.A(KEYINPUT73), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n217), .A2(new_n218), .A3(new_n202), .A4(new_n206), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n207), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT26), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n222), .A2(new_n227), .B1(G183gat), .B2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT28), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT27), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G183gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT27), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT71), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT71), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n233), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n231), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT27), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n232), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(new_n230), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT68), .A4(new_n230), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n240), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n246), .A2(KEYINPUT70), .A3(new_n247), .A4(new_n248), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n229), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n230), .A2(G183gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n234), .A2(G190gat), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT24), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OR3_X1    g055(.A1(new_n234), .A2(new_n230), .A3(KEYINPUT24), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n221), .B2(KEYINPUT23), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT64), .B1(new_n221), .B2(KEYINPUT23), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT23), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n262), .B(new_n263), .C1(G169gat), .C2(G176gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n225), .A2(new_n266), .A3(new_n226), .ZN(new_n267));
  INV_X1    g066(.A(new_n226), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT66), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n265), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n225), .A2(new_n226), .B1(KEYINPUT23), .B2(new_n221), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n265), .A2(new_n272), .A3(new_n256), .A4(new_n257), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n260), .A2(new_n271), .B1(new_n273), .B2(new_n258), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n220), .B1(new_n253), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n244), .A2(new_n245), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n248), .A2(new_n247), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n250), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n240), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n252), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n228), .ZN(new_n281));
  INV_X1    g080(.A(new_n220), .ZN(new_n282));
  INV_X1    g081(.A(new_n274), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G227gat), .ZN(new_n285));
  INV_X1    g084(.A(G233gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n275), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT32), .ZN(new_n289));
  XNOR2_X1  g088(.A(G15gat), .B(G43gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT74), .ZN(new_n291));
  INV_X1    g090(.A(G71gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(G99gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n288), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT34), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n275), .A2(new_n284), .ZN(new_n298));
  INV_X1    g097(.A(new_n287), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI211_X1 g099(.A(KEYINPUT34), .B(new_n287), .C1(new_n275), .C2(new_n284), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n296), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n296), .A2(new_n300), .A3(new_n301), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n289), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT35), .ZN(new_n306));
  XNOR2_X1  g105(.A(G78gat), .B(G106gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(G22gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT22), .ZN(new_n311));
  INV_X1    g110(.A(G211gat), .ZN(new_n312));
  INV_X1    g111(.A(G218gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G211gat), .B(G218gat), .Z(new_n316));
  AND3_X1   g115(.A1(new_n315), .A2(KEYINPUT77), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(KEYINPUT77), .B2(new_n316), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT81), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT81), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n323), .A3(KEYINPUT2), .ZN(new_n324));
  AND2_X1   g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n322), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  AND3_X1   g127(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n321), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G155gat), .B(G162gat), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n328), .A2(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT78), .B(KEYINPUT29), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n319), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n317), .B2(new_n318), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n337), .B1(new_n344), .B2(new_n338), .ZN(new_n345));
  OAI211_X1 g144(.A(G228gat), .B(G233gat), .C1(new_n342), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n339), .A2(new_n341), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n317), .A2(new_n318), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G228gat), .A2(G233gat), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n310), .A2(new_n314), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(new_n316), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(new_n340), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n316), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT3), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n349), .B(new_n350), .C1(new_n337), .C2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT31), .B(G50gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n346), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n346), .B2(new_n356), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n309), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n361), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(new_n308), .A3(new_n359), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n298), .A2(new_n299), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT34), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n298), .A2(new_n297), .A3(new_n299), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n288), .A2(new_n295), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n368), .C1(new_n369), .C2(new_n294), .ZN(new_n370));
  INV_X1    g169(.A(new_n289), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n371), .A3(new_n302), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n305), .A2(new_n306), .A3(new_n365), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n374));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n253), .B2(new_n274), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n341), .B1(new_n253), .B2(new_n274), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n374), .A2(new_n377), .B1(new_n378), .B2(new_n375), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n274), .B1(new_n280), .B2(new_n228), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n374), .B(new_n375), .C1(new_n380), .C2(new_n340), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n348), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n375), .B1(new_n380), .B2(KEYINPUT29), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n384), .A2(new_n319), .A3(new_n377), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(G1gat), .B(G29gat), .Z(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n337), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT3), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n399), .A2(new_n282), .A3(new_n339), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n400), .A2(KEYINPUT5), .A3(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n337), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT4), .B1(new_n220), .B2(new_n337), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT83), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n216), .A2(new_n219), .ZN(new_n407));
  INV_X1    g206(.A(new_n207), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n337), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n337), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n406), .A2(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n403), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n220), .B(new_n337), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(new_n402), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n399), .A2(new_n282), .A3(new_n339), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(new_n411), .A3(new_n413), .A4(new_n401), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT6), .B(new_n397), .C1(new_n416), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n403), .A2(new_n415), .B1(new_n419), .B2(new_n421), .ZN(new_n426));
  INV_X1    g225(.A(new_n397), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n403), .A2(new_n415), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n429), .A2(new_n422), .A3(new_n427), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n424), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n389), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n375), .B1(new_n380), .B2(new_n340), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n374), .B1(new_n380), .B2(new_n375), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n319), .B1(new_n435), .B2(new_n381), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n432), .B1(new_n436), .B2(new_n385), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n383), .A2(KEYINPUT30), .A3(new_n386), .A4(new_n389), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n392), .A2(new_n431), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n373), .B1(KEYINPUT86), .B2(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n438), .A2(new_n437), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n392), .A4(new_n431), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n370), .A2(new_n371), .A3(new_n302), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n371), .B1(new_n370), .B2(new_n302), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(new_n428), .B2(new_n430), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n397), .B1(new_n416), .B2(new_n423), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n426), .A2(new_n427), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n450), .A4(new_n425), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n451), .A3(new_n424), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n438), .A2(new_n437), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n381), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n385), .B1(new_n454), .B2(new_n348), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT30), .B1(new_n455), .B2(new_n389), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n446), .A2(new_n452), .A3(new_n457), .A4(new_n365), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n440), .A2(new_n443), .B1(new_n458), .B2(KEYINPUT35), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n365), .B1(new_n457), .B2(new_n452), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n362), .A2(new_n364), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n400), .B1(new_n406), .B2(new_n414), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(new_n401), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT39), .B1(new_n418), .B2(new_n402), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n462), .A2(KEYINPUT39), .A3(new_n401), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT85), .B1(new_n466), .B2(new_n397), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT83), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n412), .B1(new_n411), .B2(new_n413), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n420), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT39), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n402), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n427), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n465), .B1(new_n467), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n449), .B1(new_n475), .B2(KEYINPUT40), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  AOI211_X1 g276(.A(new_n477), .B(new_n465), .C1(new_n467), .C2(new_n474), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n392), .A2(new_n437), .A3(new_n438), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n461), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n348), .B1(new_n435), .B2(new_n381), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n384), .A2(new_n348), .A3(new_n377), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT37), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n389), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n485), .B1(new_n437), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n383), .A2(new_n386), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n487), .B1(new_n490), .B2(new_n432), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT38), .B1(new_n455), .B2(new_n486), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n489), .A2(KEYINPUT38), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n431), .B1(new_n455), .B2(new_n389), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n460), .B1(new_n481), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n305), .A2(new_n372), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT75), .B1(new_n497), .B2(KEYINPUT76), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT36), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n497), .B2(KEYINPUT75), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n459), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G43gat), .A2(G50gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(KEYINPUT15), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT90), .B(G43gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(G50gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(G43gat), .A2(G50gat), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT15), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT89), .B(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G29gat), .ZN(new_n512));
  NOR3_X1   g311(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n508), .A2(new_n510), .A3(new_n512), .A4(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n515), .B(KEYINPUT87), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n514), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT88), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n515), .A2(KEYINPUT87), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n515), .A2(KEYINPUT87), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT88), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n521), .A2(new_n526), .A3(new_n512), .ZN(new_n527));
  INV_X1    g326(.A(new_n510), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n518), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT91), .ZN(new_n531));
  INV_X1    g330(.A(G1gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT16), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n530), .A2(new_n535), .B1(new_n536), .B2(G8gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n536), .A2(G8gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT93), .B1(new_n529), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n526), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n512), .B1(new_n524), .B2(new_n525), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n528), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n517), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546));
  INV_X1    g345(.A(new_n539), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n538), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n541), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n529), .A2(new_n540), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT13), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n545), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n529), .A2(KEYINPUT17), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n540), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n550), .A2(new_n559), .A3(KEYINPUT18), .A4(new_n553), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n550), .A2(new_n559), .A3(new_n553), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G197gat), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT11), .B(G169gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT12), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n561), .B(new_n564), .C1(KEYINPUT94), .C2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n560), .A3(KEYINPUT94), .ZN(new_n572));
  INV_X1    g371(.A(new_n564), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n560), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n572), .B(new_n569), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n503), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT102), .B(G85gat), .Z(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT103), .B(G92gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT100), .B1(G85gat), .B2(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(KEYINPUT8), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT101), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(G85gat), .A3(G92gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n583), .A2(new_n586), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G99gat), .B(G106gat), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n590), .B1(new_n592), .B2(new_n588), .ZN(new_n597));
  INV_X1    g396(.A(new_n595), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n583), .A4(new_n586), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n599), .A3(KEYINPUT104), .ZN(new_n600));
  OR3_X1    g399(.A1(new_n594), .A2(KEYINPUT104), .A3(new_n595), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n557), .A2(new_n558), .A3(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n545), .B2(new_n602), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G190gat), .B(G218gat), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n608), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n610), .A3(new_n606), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  AND2_X1   g413(.A1(new_n614), .A2(KEYINPUT105), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(KEYINPUT105), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n609), .A2(new_n611), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n607), .B(new_n610), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n619), .B1(new_n620), .B2(new_n615), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n623), .A2(KEYINPUT96), .ZN(new_n624));
  XOR2_X1   g423(.A(G57gat), .B(G64gat), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(KEYINPUT96), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G71gat), .B(G78gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(new_n624), .A3(new_n626), .A4(new_n625), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n548), .B1(KEYINPUT21), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G127gat), .B(G155gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT99), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT98), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n639), .B(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n633), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n632), .B1(new_n599), .B2(new_n596), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n602), .B2(new_n632), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n650), .B2(KEYINPUT10), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(G120gat), .B(G148gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT106), .ZN(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n653), .A2(new_n655), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n622), .A2(new_n647), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT107), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n580), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n452), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT108), .B(G1gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1324gat));
  NAND3_X1  g470(.A1(new_n580), .A2(new_n480), .A3(new_n667), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT16), .B(G8gat), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT109), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(KEYINPUT42), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(G8gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(KEYINPUT42), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(G1325gat));
  OAI21_X1  g477(.A(G15gat), .B1(new_n668), .B2(new_n502), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n497), .A2(G15gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n668), .B2(new_n680), .ZN(G1326gat));
  NOR2_X1   g480(.A1(new_n668), .A2(new_n365), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT43), .B(G22gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  INV_X1    g483(.A(KEYINPUT113), .ZN(new_n685));
  INV_X1    g484(.A(G29gat), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT112), .ZN(new_n687));
  INV_X1    g486(.A(new_n576), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n664), .A2(new_n647), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT44), .B1(new_n503), .B2(new_n622), .ZN(new_n693));
  INV_X1    g492(.A(new_n465), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n466), .A2(KEYINPUT85), .A3(new_n397), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n473), .B1(new_n472), .B2(new_n427), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n477), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n475), .A2(KEYINPUT40), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n480), .A2(new_n698), .A3(new_n449), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n495), .A2(new_n365), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n460), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT75), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT76), .B1(new_n444), .B2(new_n445), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT75), .B1(new_n444), .B2(new_n445), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n703), .A2(new_n704), .B1(new_n705), .B2(KEYINPUT36), .ZN(new_n706));
  AOI211_X1 g505(.A(KEYINPUT75), .B(new_n500), .C1(new_n497), .C2(KEYINPUT76), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n701), .B(new_n702), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n439), .A2(KEYINPUT86), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n444), .A2(new_n445), .A3(new_n461), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n709), .A2(new_n710), .A3(new_n443), .A4(new_n306), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n457), .A2(new_n452), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n305), .A2(new_n372), .A3(new_n365), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT35), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n711), .A2(new_n714), .A3(KEYINPUT111), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT111), .B1(new_n711), .B2(new_n714), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n708), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n622), .A2(KEYINPUT44), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n687), .B(new_n692), .C1(new_n693), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n711), .A2(new_n714), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n711), .A2(new_n714), .A3(KEYINPUT111), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n723), .A2(new_n724), .B1(new_n496), .B2(new_n502), .ZN(new_n725));
  INV_X1    g524(.A(new_n718), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n622), .B1(new_n708), .B2(new_n721), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  OAI22_X1  g527(.A1(new_n725), .A2(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT112), .B1(new_n729), .B2(new_n691), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n720), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n452), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n686), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n690), .A2(new_n622), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n580), .A2(new_n686), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n685), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n737), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n720), .A2(new_n730), .A3(new_n452), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n739), .B(KEYINPUT113), .C1(new_n740), .C2(new_n686), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(G1328gat));
  AND2_X1   g541(.A1(new_n580), .A2(new_n734), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n511), .B1(new_n744), .B2(KEYINPUT46), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n480), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n691), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n687), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n729), .A2(KEYINPUT112), .A3(new_n691), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(new_n480), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n511), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n748), .B1(new_n755), .B2(new_n756), .ZN(G1329gat));
  NAND2_X1  g556(.A1(new_n580), .A2(new_n734), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n758), .A2(new_n497), .A3(new_n507), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n507), .B1(new_n749), .B2(new_n502), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n502), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n731), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n759), .B1(new_n765), .B2(new_n507), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n763), .B1(new_n766), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g566(.A(G50gat), .B1(new_n749), .B2(new_n365), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n758), .A2(KEYINPUT116), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n365), .A2(G50gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n758), .B2(KEYINPUT116), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n768), .B(KEYINPUT48), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n769), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n731), .A2(new_n461), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(G50gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n772), .B1(new_n775), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g575(.A(new_n647), .ZN(new_n777));
  NOR4_X1   g576(.A1(new_n725), .A2(new_n576), .A3(new_n777), .A4(new_n621), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n664), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n452), .B(KEYINPUT117), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n785));
  INV_X1    g584(.A(G64gat), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n780), .B(new_n480), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1333gat));
  OAI21_X1  g588(.A(G71gat), .B1(new_n779), .B2(new_n502), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n497), .A2(new_n665), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n778), .A2(new_n292), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n461), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g596(.A1(new_n576), .A2(new_n647), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n717), .A2(new_n621), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT51), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(KEYINPUT118), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n732), .A2(new_n581), .A3(new_n664), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n729), .A2(new_n664), .A3(new_n798), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n452), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n805), .A2(new_n806), .B1(new_n581), .B2(new_n808), .ZN(G1336gat));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  INV_X1    g609(.A(new_n582), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n807), .B2(new_n457), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n457), .A2(G92gat), .A3(new_n665), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n810), .B(new_n812), .C1(new_n805), .C2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n800), .B2(new_n813), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT52), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1337gat));
  OAI21_X1  g616(.A(G99gat), .B1(new_n807), .B2(new_n502), .ZN(new_n818));
  INV_X1    g617(.A(G99gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n791), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n805), .B2(new_n820), .ZN(G1338gat));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  OAI21_X1  g621(.A(G106gat), .B1(new_n807), .B2(new_n365), .ZN(new_n823));
  OR3_X1    g622(.A1(new_n665), .A2(G106gat), .A3(new_n365), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n822), .B(new_n823), .C1(new_n805), .C2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n800), .B2(new_n824), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1339gat));
  NOR2_X1   g627(.A1(new_n666), .A2(new_n576), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT119), .Z(new_n830));
  NOR2_X1   g629(.A1(new_n653), .A2(KEYINPUT54), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n662), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n651), .B2(new_n652), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n654), .B(new_n648), .C1(new_n650), .C2(KEYINPUT10), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n835), .B1(new_n834), .B2(new_n836), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n832), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n653), .A2(KEYINPUT54), .A3(new_n836), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT120), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n837), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n842), .A2(new_n576), .A3(new_n663), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n561), .A2(new_n564), .A3(new_n570), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n552), .A2(new_n554), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n553), .B1(new_n550), .B2(new_n559), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n568), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n664), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n621), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n846), .A2(new_n663), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT55), .B1(new_n845), .B2(new_n832), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n621), .A2(new_n848), .A3(new_n851), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT121), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n777), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n854), .A2(KEYINPUT121), .A3(new_n858), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n830), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n781), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n713), .A2(new_n480), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(G113gat), .B1(new_n867), .B2(new_n576), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n452), .A2(new_n480), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n710), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n862), .A2(KEYINPUT122), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT122), .B1(new_n862), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n578), .A2(G113gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n868), .B1(new_n874), .B2(new_n875), .ZN(G1340gat));
  AOI21_X1  g675(.A(G120gat), .B1(new_n867), .B2(new_n664), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n664), .A2(G120gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n874), .B2(new_n878), .ZN(G1341gat));
  NOR3_X1   g678(.A1(new_n872), .A2(new_n873), .A3(new_n777), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n211), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n647), .A2(new_n211), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT123), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885));
  OAI221_X1 g684(.A(new_n885), .B1(new_n866), .B2(new_n882), .C1(new_n880), .C2(new_n211), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1342gat));
  NAND2_X1  g686(.A1(new_n621), .A2(new_n209), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n866), .A2(KEYINPUT56), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT56), .B1(new_n866), .B2(new_n888), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n872), .A2(new_n873), .A3(new_n622), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n889), .B(new_n890), .C1(new_n209), .C2(new_n891), .ZN(G1343gat));
  AND2_X1   g691(.A1(new_n502), .A2(new_n869), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT57), .B1(new_n862), .B2(new_n461), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n365), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n858), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n855), .A2(new_n856), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n578), .A2(new_n899), .B1(new_n664), .B2(new_n852), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n900), .B2(new_n621), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n777), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n897), .B1(new_n902), .B2(new_n830), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n893), .B1(new_n894), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G141gat), .B1(new_n904), .B2(new_n579), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n862), .A2(new_n782), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n502), .A2(new_n461), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n906), .A2(new_n480), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n579), .A2(G141gat), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT58), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n576), .B(new_n893), .C1(new_n894), .C2(new_n903), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n912), .A2(G141gat), .B1(new_n908), .B2(new_n909), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1344gat));
  OR2_X1    g714(.A1(new_n893), .A2(KEYINPUT124), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n893), .A2(KEYINPUT124), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n664), .A3(new_n917), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n901), .A2(new_n777), .B1(new_n667), .B2(new_n579), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n895), .B1(new_n919), .B2(new_n365), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n862), .A2(new_n896), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(G148gat), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT59), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(KEYINPUT59), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n904), .B2(new_n665), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n908), .A2(new_n923), .A3(new_n664), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1345gat));
  OAI211_X1 g728(.A(new_n647), .B(new_n893), .C1(new_n894), .C2(new_n903), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G155gat), .ZN(new_n931));
  INV_X1    g730(.A(G155gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n908), .A2(new_n932), .A3(new_n647), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n931), .A2(KEYINPUT125), .A3(new_n933), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1346gat));
  INV_X1    g737(.A(G162gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n904), .A2(new_n939), .A3(new_n622), .ZN(new_n940));
  AOI21_X1  g739(.A(G162gat), .B1(new_n908), .B2(new_n621), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(G1347gat));
  NOR2_X1   g741(.A1(new_n863), .A2(new_n732), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n713), .A2(new_n457), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(G169gat), .B1(new_n945), .B2(new_n576), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n782), .A2(new_n457), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n365), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n863), .A2(new_n497), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n578), .A2(G169gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(G1348gat));
  AOI21_X1  g750(.A(G176gat), .B1(new_n945), .B2(new_n664), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n863), .A2(new_n948), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n791), .A2(G176gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(G1349gat));
  INV_X1    g754(.A(new_n948), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n862), .A2(new_n446), .A3(new_n647), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G183gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n777), .B1(new_n239), .B2(new_n237), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n862), .A2(new_n452), .A3(new_n944), .A4(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n958), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n945), .A2(new_n230), .A3(new_n621), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n949), .A2(new_n621), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(G190gat), .ZN(new_n969));
  AOI211_X1 g768(.A(KEYINPUT61), .B(new_n230), .C1(new_n949), .C2(new_n621), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  NOR2_X1   g770(.A1(new_n907), .A2(new_n457), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n943), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n576), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n920), .A2(new_n921), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n947), .A2(new_n502), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n578), .A2(G197gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  NOR2_X1   g778(.A1(new_n665), .A2(G204gat), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n943), .A2(new_n972), .A3(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n975), .A2(new_n664), .A3(new_n976), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G204gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n981), .A2(new_n982), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(G1353gat));
  NAND3_X1  g786(.A1(new_n973), .A2(new_n312), .A3(new_n647), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n975), .A2(new_n647), .A3(new_n976), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n989), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT63), .B1(new_n989), .B2(G211gat), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(G1354gat));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n621), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(G218gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n973), .A2(new_n313), .A3(new_n621), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(G1355gat));
endmodule


