//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n809, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  AND2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT73), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT73), .ZN(new_n210));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n206), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n219), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT75), .A3(new_n217), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT75), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(new_n218), .B2(new_n219), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n204), .A2(new_n205), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n217), .A2(KEYINPUT2), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n223), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT76), .ZN(new_n230));
  INV_X1    g029(.A(G134gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G127gat), .ZN(new_n232));
  INV_X1    g031(.A(G127gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G134gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G120gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(KEYINPUT1), .ZN(new_n237));
  INV_X1    g036(.A(G120gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G113gat), .ZN(new_n239));
  INV_X1    g038(.A(G113gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G120gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n237), .A2(new_n245), .A3(KEYINPUT77), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT77), .B1(new_n237), .B2(new_n245), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT76), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n221), .A2(new_n249), .A3(new_n228), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n230), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n251), .A2(KEYINPUT79), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT79), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n230), .A2(new_n248), .A3(new_n253), .A4(new_n250), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n221), .A2(new_n228), .A3(new_n245), .A4(new_n237), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n203), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n230), .A2(KEYINPUT3), .A3(new_n250), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n221), .A2(new_n259), .A3(new_n228), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n237), .A2(new_n245), .A3(KEYINPUT77), .ZN(new_n261));
  INV_X1    g060(.A(new_n247), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n203), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n255), .A2(KEYINPUT4), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n242), .A2(new_n244), .B1(new_n232), .B2(new_n234), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n237), .A2(new_n245), .A3(KEYINPUT69), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n273), .A2(new_n223), .B1(new_n216), .B2(new_n220), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n266), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT78), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n265), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n229), .B1(new_n271), .B2(new_n270), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n278), .A2(KEYINPUT78), .A3(new_n266), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n264), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n257), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n264), .A2(new_n281), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n272), .A2(new_n266), .A3(new_n274), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT82), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n255), .A2(KEYINPUT4), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT82), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n288), .A3(new_n266), .A4(new_n274), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G1gat), .B(G29gat), .Z(new_n293));
  XNOR2_X1  g092(.A(G57gat), .B(G85gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(KEYINPUT6), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G226gat), .ZN(new_n299));
  INV_X1    g098(.A(G233gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(KEYINPUT29), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT23), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n305), .A2(KEYINPUT25), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  AND2_X1   g109(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n313), .A2(KEYINPUT65), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT65), .B1(new_n313), .B2(new_n314), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n309), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n312), .B(KEYINPUT66), .C1(new_n315), .C2(new_n316), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT64), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n308), .B1(new_n304), .B2(KEYINPUT23), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n306), .A2(G169gat), .A3(G176gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n313), .A2(new_n314), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n312), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n305), .A2(KEYINPUT64), .A3(new_n307), .A4(new_n308), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n321), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT27), .B(G183gat), .ZN(new_n335));
  INV_X1    g134(.A(G190gat), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G183gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT27), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G183gat), .ZN(new_n341));
  AND4_X1   g140(.A1(new_n334), .A2(new_n339), .A3(new_n341), .A4(new_n336), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n333), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n341), .A3(new_n336), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT67), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n335), .A2(new_n334), .A3(new_n336), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(KEYINPUT28), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n304), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT26), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n308), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n304), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT68), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT68), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n348), .B(new_n353), .C1(new_n304), .C2(new_n350), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n343), .A2(new_n347), .A3(new_n352), .A4(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n303), .B1(new_n332), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT71), .ZN(new_n357));
  AND4_X1   g156(.A1(new_n343), .A2(new_n347), .A3(new_n352), .A4(new_n354), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n319), .A2(new_n320), .B1(new_n329), .B2(new_n330), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n332), .A2(KEYINPUT71), .A3(new_n355), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n356), .B1(new_n362), .B2(new_n301), .ZN(new_n363));
  OR2_X1    g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT22), .ZN(new_n366));
  NAND2_X1  g165(.A1(G211gat), .A2(G218gat), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n364), .A2(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT70), .ZN(new_n370));
  INV_X1    g169(.A(G211gat), .ZN(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n373), .B2(new_n367), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n370), .A3(new_n367), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n369), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n376), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n368), .B1(new_n378), .B2(new_n374), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT72), .B1(new_n363), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n332), .A2(new_n355), .A3(new_n301), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n383), .B(new_n381), .C1(new_n362), .C2(new_n303), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT72), .ZN(new_n385));
  INV_X1    g184(.A(new_n301), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n360), .B2(new_n361), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n385), .B(new_n380), .C1(new_n387), .C2(new_n356), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  NAND4_X1  g190(.A1(new_n382), .A2(new_n384), .A3(new_n388), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n297), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n283), .A2(new_n393), .A3(new_n291), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n283), .B2(new_n291), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n298), .B(new_n392), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n391), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n384), .A3(new_n388), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n401), .B2(KEYINPUT37), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT37), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n384), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n405), .B2(new_n382), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT38), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n363), .A2(new_n381), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT90), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT90), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n363), .A2(new_n410), .A3(new_n381), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n383), .B1(new_n362), .B2(new_n303), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n380), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT38), .B1(new_n414), .B2(KEYINPUT37), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n362), .A2(new_n301), .ZN(new_n416));
  INV_X1    g215(.A(new_n356), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n385), .B1(new_n418), .B2(new_n380), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n400), .B1(new_n419), .B2(new_n404), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n400), .A2(KEYINPUT37), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n415), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n407), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G78gat), .B(G106gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT31), .B(G50gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n380), .B1(new_n260), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G228gat), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n430), .A2(new_n431), .A3(new_n300), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT29), .B1(new_n377), .B2(new_n379), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n259), .B1(new_n433), .B2(KEYINPUT85), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n380), .A2(KEYINPUT85), .A3(new_n429), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n230), .A2(new_n250), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n377), .A2(new_n379), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n369), .A2(new_n375), .A3(KEYINPUT84), .A4(new_n376), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n429), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n274), .B1(new_n442), .B2(new_n259), .ZN(new_n443));
  OAI22_X1  g242(.A1(new_n443), .A2(new_n430), .B1(new_n431), .B2(new_n300), .ZN(new_n444));
  INV_X1    g243(.A(G22gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n438), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n445), .B1(new_n438), .B2(new_n444), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n428), .B(new_n446), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n447), .A2(new_n448), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n447), .A2(KEYINPUT86), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n446), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n438), .A2(new_n444), .A3(KEYINPUT86), .A4(new_n445), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n427), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n450), .A2(new_n452), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n258), .A2(new_n263), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n288), .B1(new_n278), .B2(new_n266), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n289), .A2(new_n287), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n203), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n251), .A2(KEYINPUT79), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(new_n202), .A3(new_n255), .A4(new_n254), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n254), .A2(new_n255), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n468), .A2(KEYINPUT89), .A3(new_n202), .A4(new_n464), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n463), .A2(new_n467), .A3(KEYINPUT39), .A4(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n202), .B1(new_n290), .B2(new_n459), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT39), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n297), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n470), .A2(KEYINPUT40), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT40), .B1(new_n470), .B2(new_n473), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n474), .A2(new_n475), .A3(new_n397), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n392), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n400), .A2(new_n477), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n405), .A2(new_n382), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n420), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n458), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n424), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  XOR2_X1   g283(.A(G15gat), .B(G43gat), .Z(new_n485));
  XNOR2_X1  g284(.A(G71gat), .B(G99gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n332), .A2(new_n271), .A3(new_n270), .A4(new_n355), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n272), .B1(new_n358), .B2(new_n359), .ZN(new_n490));
  INV_X1    g289(.A(G227gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(new_n300), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n489), .A2(new_n490), .ZN(new_n497));
  INV_X1    g296(.A(new_n492), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI211_X1 g298(.A(KEYINPUT34), .B(new_n492), .C1(new_n489), .C2(new_n490), .ZN(new_n500));
  OR3_X1    g299(.A1(new_n495), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n493), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT32), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n501), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n484), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n505), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n495), .A2(new_n499), .A3(new_n500), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n509), .A2(new_n510), .B1(new_n503), .B2(new_n502), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT36), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT83), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT78), .B1(new_n278), .B2(new_n266), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n275), .A2(new_n276), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n265), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n281), .B1(new_n518), .B2(new_n264), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n519), .A2(new_n257), .B1(new_n290), .B2(new_n284), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n515), .B1(new_n520), .B2(new_n393), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT6), .B1(new_n520), .B2(new_n393), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n397), .A2(KEYINPUT83), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n481), .B1(new_n298), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n446), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n526), .A2(new_n447), .A3(KEYINPUT86), .ZN(new_n527));
  OAI22_X1  g326(.A1(new_n527), .A2(new_n456), .B1(new_n449), .B2(new_n451), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI221_X1 g329(.A(KEYINPUT88), .B1(new_n449), .B2(new_n451), .C1(new_n527), .C2(new_n456), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n514), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n512), .A3(new_n511), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n534), .B1(new_n525), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n298), .B1(new_n396), .B2(new_n397), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n534), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n535), .A2(new_n539), .A3(new_n481), .ZN(new_n540));
  OAI22_X1  g339(.A1(new_n483), .A2(new_n533), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n298), .ZN(new_n544));
  INV_X1    g343(.A(new_n481), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT35), .B1(new_n546), .B2(new_n535), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n536), .A2(new_n534), .A3(new_n538), .A4(new_n545), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n530), .A2(new_n531), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n546), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n424), .A2(new_n482), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n514), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n553), .A3(KEYINPUT91), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n555));
  XNOR2_X1  g354(.A(G15gat), .B(G22gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT16), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(G1gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(G1gat), .B2(new_n556), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(G8gat), .Z(new_n560));
  NOR2_X1   g359(.A1(G29gat), .A2(G36gat), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n561), .A2(KEYINPUT14), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(KEYINPUT14), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT92), .B(G36gat), .Z(new_n564));
  INV_X1    g363(.A(G29gat), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G43gat), .B(G50gat), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n567), .A2(KEYINPUT15), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n566), .A2(KEYINPUT93), .A3(new_n568), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n567), .B(KEYINPUT15), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT94), .B1(new_n574), .B2(new_n566), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n567), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n578));
  INV_X1    g377(.A(new_n564), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G29gat), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n562), .A2(new_n563), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n577), .A2(new_n578), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n573), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT95), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n571), .A2(new_n572), .B1(new_n575), .B2(new_n582), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(KEYINPUT17), .ZN(new_n589));
  AND4_X1   g388(.A1(new_n587), .A2(new_n573), .A3(new_n583), .A4(KEYINPUT17), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n560), .B(new_n586), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n560), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n584), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT96), .B1(new_n588), .B2(new_n560), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT18), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G113gat), .B(G141gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G197gat), .ZN(new_n602));
  XOR2_X1   g401(.A(KEYINPUT11), .B(G169gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT12), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n591), .A2(KEYINPUT18), .A3(new_n592), .A4(new_n597), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n597), .B1(new_n584), .B2(new_n593), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n592), .B(KEYINPUT13), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n600), .A2(new_n606), .A3(new_n607), .A4(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n598), .A2(new_n599), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n606), .B1(new_n613), .B2(new_n607), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n555), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n607), .A3(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n605), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(KEYINPUT97), .A3(new_n611), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n543), .A2(new_n554), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(G71gat), .A2(G78gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(G71gat), .A2(G78gat), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(KEYINPUT9), .B2(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(KEYINPUT98), .B(G57gat), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(G64gat), .ZN(new_n626));
  INV_X1    g425(.A(G64gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(G57gat), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n624), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G57gat), .B(G64gat), .Z(new_n630));
  AOI211_X1 g429(.A(new_n622), .B(new_n623), .C1(new_n630), .C2(KEYINPUT9), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT21), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G127gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G183gat), .B(G211gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n636), .A2(new_n233), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n636), .A2(new_n233), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n641), .A2(new_n642), .A3(new_n638), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n560), .B1(new_n633), .B2(new_n632), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n645), .B(KEYINPUT99), .Z(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n647));
  INV_X1    g446(.A(G155gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n646), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n649), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n646), .B(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n643), .B2(new_n640), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G232gat), .A2(G233gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(KEYINPUT41), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT100), .ZN(new_n659));
  XNOR2_X1  g458(.A(G134gat), .B(G162gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT8), .ZN(new_n663));
  NAND2_X1  g462(.A1(G99gat), .A2(G106gat), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(KEYINPUT102), .A2(G99gat), .A3(G106gat), .ZN(new_n667));
  INV_X1    g466(.A(G85gat), .ZN(new_n668));
  INV_X1    g467(.A(G92gat), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n666), .A2(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT103), .ZN(new_n671));
  AOI211_X1 g470(.A(new_n668), .B(new_n669), .C1(KEYINPUT101), .C2(KEYINPUT7), .ZN(new_n672));
  NOR2_X1   g471(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(G99gat), .B(G106gat), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n676), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n671), .A2(new_n678), .A3(new_n674), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n586), .B(new_n680), .C1(new_n589), .C2(new_n590), .ZN(new_n681));
  INV_X1    g480(.A(new_n680), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n682), .A2(new_n584), .B1(KEYINPUT41), .B2(new_n657), .ZN(new_n683));
  XNOR2_X1  g482(.A(G190gat), .B(G218gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT104), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n681), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(new_n681), .B2(new_n683), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n662), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n681), .A2(new_n683), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n685), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n661), .A3(new_n687), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n655), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n632), .B1(new_n679), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n677), .B(new_n679), .C1(new_n696), .C2(new_n632), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT10), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT10), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n680), .A2(new_n701), .A3(new_n632), .ZN(new_n702));
  INV_X1    g501(.A(G230gat), .ZN(new_n703));
  OAI22_X1  g502(.A1(new_n700), .A2(new_n702), .B1(new_n703), .B2(new_n300), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n300), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n698), .A2(new_n699), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(G120gat), .B(G148gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(G176gat), .B(G204gat), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n707), .B(new_n708), .Z(new_n709));
  AND3_X1   g508(.A1(new_n704), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n704), .B2(new_n706), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n695), .A2(KEYINPUT106), .A3(new_n712), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n621), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n544), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(G1gat), .Z(G1324gat));
  XOR2_X1   g520(.A(KEYINPUT16), .B(G8gat), .Z(new_n722));
  NAND4_X1  g521(.A1(new_n621), .A2(new_n481), .A3(new_n718), .A4(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G8gat), .B1(new_n719), .B2(new_n545), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n723), .ZN(new_n725));
  MUX2_X1   g524(.A(new_n723), .B(new_n725), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g525(.A(G15gat), .B1(new_n719), .B2(new_n514), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n506), .A2(new_n507), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n729), .A2(G15gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n719), .B2(new_n730), .ZN(G1326gat));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n719), .B2(new_n532), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n621), .A2(KEYINPUT107), .A3(new_n550), .A4(new_n718), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT43), .B(G22gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1327gat));
  NAND2_X1  g536(.A1(new_n617), .A2(new_n611), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n655), .A2(new_n738), .A3(new_n712), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n543), .A2(new_n554), .A3(new_n694), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT44), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n690), .A2(new_n693), .A3(KEYINPUT109), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT109), .B1(new_n690), .B2(new_n693), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n551), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n550), .A2(new_n546), .A3(KEYINPUT108), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n748), .A2(new_n552), .A3(new_n514), .A4(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n746), .B1(new_n750), .B2(new_n549), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n739), .B1(new_n741), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G29gat), .B1(new_n754), .B2(new_n544), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n756));
  INV_X1    g555(.A(new_n655), .ZN(new_n757));
  INV_X1    g556(.A(new_n694), .ZN(new_n758));
  INV_X1    g557(.A(new_n712), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n543), .A2(new_n554), .A3(new_n620), .A4(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n544), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n565), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n756), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n761), .A2(new_n756), .A3(new_n763), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n755), .A2(new_n764), .A3(new_n765), .ZN(G1328gat));
  OAI21_X1  g565(.A(new_n579), .B1(new_n754), .B2(new_n545), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n481), .A2(new_n564), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT46), .B1(new_n761), .B2(new_n768), .ZN(new_n769));
  OR3_X1    g568(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n768), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(G1329gat));
  AOI21_X1  g570(.A(new_n751), .B1(new_n740), .B2(KEYINPUT44), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n772), .A2(new_n514), .A3(new_n739), .ZN(new_n773));
  INV_X1    g572(.A(G43gat), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT110), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n621), .A2(new_n774), .A3(new_n728), .A4(new_n760), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI221_X1 g578(.A(new_n776), .B1(KEYINPUT110), .B2(KEYINPUT47), .C1(new_n773), .C2(new_n774), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(G1330gat));
  INV_X1    g580(.A(KEYINPUT48), .ZN(new_n782));
  INV_X1    g581(.A(G50gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n550), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n761), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT111), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n783), .B1(new_n753), .B2(new_n550), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n782), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n753), .B2(new_n458), .ZN(new_n790));
  NOR4_X1   g589(.A1(new_n772), .A2(KEYINPUT112), .A3(new_n528), .A4(new_n739), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n790), .A2(new_n791), .A3(new_n783), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT48), .B1(new_n761), .B2(new_n784), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n788), .B1(new_n792), .B2(new_n793), .ZN(G1331gat));
  NAND2_X1  g593(.A1(new_n750), .A2(new_n549), .ZN(new_n795));
  NOR4_X1   g594(.A1(new_n655), .A2(new_n738), .A3(new_n694), .A4(new_n712), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n544), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(new_n625), .ZN(G1332gat));
  NOR2_X1   g598(.A1(new_n797), .A2(new_n545), .ZN(new_n800));
  NOR2_X1   g599(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n801));
  AND2_X1   g600(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n800), .B2(new_n801), .ZN(G1333gat));
  OR3_X1    g603(.A1(new_n797), .A2(G71gat), .A3(new_n729), .ZN(new_n805));
  OAI21_X1  g604(.A(G71gat), .B1(new_n797), .B2(new_n514), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n807), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g607(.A1(new_n797), .A2(new_n532), .ZN(new_n809));
  XOR2_X1   g608(.A(KEYINPUT113), .B(G78gat), .Z(new_n810));
  XNOR2_X1  g609(.A(new_n809), .B(new_n810), .ZN(G1335gat));
  NOR3_X1   g610(.A1(new_n757), .A2(new_n738), .A3(new_n758), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT51), .B1(new_n795), .B2(new_n812), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n759), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n668), .A3(new_n762), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n757), .A2(new_n738), .A3(new_n712), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT114), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n772), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G85gat), .B1(new_n822), .B2(new_n544), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1336gat));
  OAI21_X1  g623(.A(G92gat), .B1(new_n822), .B2(new_n545), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n545), .A2(G92gat), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n759), .B(new_n827), .C1(new_n815), .C2(new_n816), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n772), .A2(new_n821), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n669), .B1(new_n830), .B2(new_n481), .ZN(new_n831));
  INV_X1    g630(.A(new_n828), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT52), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n829), .A2(new_n833), .ZN(G1337gat));
  INV_X1    g633(.A(G99gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n818), .A2(new_n835), .A3(new_n728), .ZN(new_n836));
  OAI21_X1  g635(.A(G99gat), .B1(new_n822), .B2(new_n514), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1338gat));
  OAI21_X1  g637(.A(G106gat), .B1(new_n822), .B2(new_n528), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n712), .A2(new_n528), .A3(G106gat), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT53), .B1(new_n817), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n830), .A2(new_n550), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n840), .B(KEYINPUT115), .Z(new_n844));
  AOI22_X1  g643(.A1(new_n843), .A2(G106gat), .B1(new_n817), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(G1339gat));
  NOR2_X1   g646(.A1(new_n713), .A2(new_n738), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n698), .A2(new_n699), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n701), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n632), .A2(new_n701), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n682), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n705), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n705), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT54), .B1(new_n855), .B2(new_n700), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n709), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n704), .B2(KEYINPUT54), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n849), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n853), .A2(new_n705), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n851), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n849), .B1(new_n863), .B2(new_n704), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n709), .B1(new_n854), .B2(new_n861), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n704), .A2(new_n706), .A3(new_n709), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n860), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n608), .A2(new_n609), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n592), .B1(new_n591), .B2(new_n597), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n604), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n611), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(new_n744), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n712), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n868), .B2(new_n738), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n876), .B2(new_n744), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n848), .B1(new_n877), .B2(new_n655), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n550), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n544), .A2(new_n481), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n728), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(new_n240), .A3(new_n619), .ZN(new_n882));
  INV_X1    g681(.A(new_n875), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n710), .B1(new_n864), .B2(new_n865), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n738), .A2(new_n884), .A3(new_n860), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n744), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n742), .A2(new_n743), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n873), .A2(new_n884), .A3(new_n860), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n655), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n713), .A2(new_n738), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n762), .A3(new_n536), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT116), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n545), .A3(new_n738), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n882), .B1(new_n895), .B2(new_n240), .ZN(G1340gat));
  NOR3_X1   g695(.A1(new_n881), .A2(new_n238), .A3(new_n712), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n545), .A3(new_n759), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n238), .ZN(G1341gat));
  OAI21_X1  g698(.A(G127gat), .B1(new_n881), .B2(new_n655), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n894), .A2(new_n545), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n757), .A2(new_n233), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(G1342gat));
  NOR3_X1   g702(.A1(new_n758), .A2(new_n481), .A3(G134gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n894), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n906));
  OAI21_X1  g705(.A(G134gat), .B1(new_n881), .B2(new_n758), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G1343gat));
  AOI21_X1  g708(.A(new_n528), .B1(new_n508), .B2(new_n513), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n762), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n481), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n207), .A3(new_n620), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n880), .A2(new_n514), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT57), .B1(new_n892), .B2(new_n458), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n550), .A2(KEYINPUT57), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(new_n857), .B2(new_n859), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n863), .A2(new_n704), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n865), .A2(new_n923), .A3(KEYINPUT117), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n922), .A2(new_n924), .A3(new_n849), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n925), .A2(new_n615), .A3(new_n618), .A4(new_n884), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n694), .B1(new_n926), .B2(new_n883), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n655), .B1(new_n927), .B2(new_n889), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n920), .B1(new_n928), .B2(new_n891), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n918), .B1(new_n919), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n916), .B1(new_n930), .B2(new_n619), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G141gat), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n930), .A2(new_n916), .A3(new_n619), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n915), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n738), .B(new_n918), .C1(new_n919), .C2(new_n929), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G141gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n913), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT118), .B1(new_n937), .B2(KEYINPUT58), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n939));
  AOI211_X1 g738(.A(new_n939), .B(new_n914), .C1(new_n936), .C2(new_n913), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n934), .B1(new_n938), .B2(new_n940), .ZN(G1344gat));
  NAND3_X1  g740(.A1(new_n912), .A2(new_n208), .A3(new_n759), .ZN(new_n942));
  INV_X1    g741(.A(new_n930), .ZN(new_n943));
  AOI211_X1 g742(.A(KEYINPUT59), .B(new_n208), .C1(new_n943), .C2(new_n759), .ZN(new_n944));
  XNOR2_X1  g743(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n532), .A2(KEYINPUT57), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n926), .A2(new_n883), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n758), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n868), .A2(new_n694), .A3(new_n873), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n757), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n715), .A2(new_n619), .A3(new_n716), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n946), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT57), .B1(new_n878), .B2(new_n528), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n953), .A2(new_n954), .A3(new_n759), .A4(new_n918), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n945), .B1(new_n955), .B2(G148gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n942), .B1(new_n944), .B2(new_n956), .ZN(G1345gat));
  OAI21_X1  g756(.A(G155gat), .B1(new_n930), .B2(new_n655), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n912), .A2(new_n648), .A3(new_n757), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1346gat));
  OAI21_X1  g759(.A(G162gat), .B1(new_n930), .B2(new_n887), .ZN(new_n961));
  OR3_X1    g760(.A1(new_n758), .A2(new_n481), .A3(G162gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n911), .B2(new_n962), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n762), .A2(new_n545), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n892), .A2(new_n536), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(G169gat), .B1(new_n965), .B2(new_n738), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n728), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT121), .Z(new_n968));
  NAND2_X1  g767(.A1(new_n879), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n620), .A2(G169gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT122), .ZN(G1348gat));
  NAND4_X1  g772(.A1(new_n879), .A2(G176gat), .A3(new_n759), .A4(new_n968), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n974), .A2(KEYINPUT123), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n965), .A2(new_n759), .ZN(new_n976));
  INV_X1    g775(.A(G176gat), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n974), .A2(KEYINPUT123), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT124), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n975), .A2(new_n982), .A3(new_n978), .A4(new_n979), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1349gat));
  OAI21_X1  g783(.A(G183gat), .B1(new_n969), .B2(new_n655), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n965), .A2(new_n335), .A3(new_n757), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g786(.A(new_n987), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g787(.A1(new_n965), .A2(new_n336), .A3(new_n744), .ZN(new_n989));
  OAI21_X1  g788(.A(G190gat), .B1(new_n969), .B2(new_n758), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n990), .A2(KEYINPUT61), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n990), .A2(KEYINPUT61), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1351gat));
  AND3_X1   g792(.A1(new_n892), .A2(new_n910), .A3(new_n964), .ZN(new_n994));
  AOI21_X1  g793(.A(G197gat), .B1(new_n994), .B2(new_n738), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n964), .A2(new_n514), .ZN(new_n996));
  XOR2_X1   g795(.A(new_n996), .B(KEYINPUT125), .Z(new_n997));
  NAND3_X1  g796(.A1(new_n953), .A2(new_n954), .A3(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(new_n998), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n620), .A2(G197gat), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n995), .B1(new_n999), .B2(new_n1000), .ZN(G1352gat));
  NOR2_X1   g800(.A1(new_n712), .A2(G204gat), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n892), .A2(new_n910), .A3(new_n964), .A4(new_n1002), .ZN(new_n1003));
  XOR2_X1   g802(.A(new_n1003), .B(KEYINPUT62), .Z(new_n1004));
  OAI21_X1  g803(.A(G204gat), .B1(new_n998), .B2(new_n712), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1006), .B(new_n1007), .ZN(G1353gat));
  NAND3_X1  g807(.A1(new_n994), .A2(new_n371), .A3(new_n757), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n996), .A2(new_n655), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n953), .A2(new_n954), .A3(new_n1010), .ZN(new_n1011));
  AND3_X1   g810(.A1(new_n1011), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1012));
  AOI21_X1  g811(.A(KEYINPUT63), .B1(new_n1011), .B2(G211gat), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1009), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g815(.A(KEYINPUT127), .B(new_n1009), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1016), .A2(new_n1017), .ZN(G1354gat));
  OAI21_X1  g817(.A(G218gat), .B1(new_n998), .B2(new_n758), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n994), .A2(new_n372), .A3(new_n744), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1019), .A2(new_n1020), .ZN(G1355gat));
endmodule


