//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(KEYINPUT64), .A3(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(new_n190), .B2(G146), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n192), .A2(KEYINPUT66), .A3(new_n194), .A4(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n194), .A2(new_n189), .A3(new_n196), .A4(new_n191), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n190), .C2(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(G128), .A3(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n197), .A2(new_n200), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  OR2_X1    g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n190), .A2(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n188), .A2(G143), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n211), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n194), .A2(new_n189), .A3(new_n191), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n210), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G224), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT7), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n210), .A2(KEYINPUT7), .A3(new_n222), .A4(new_n219), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(new_n228), .B2(KEYINPUT81), .ZN(new_n229));
  INV_X1    g043(.A(G101), .ZN(new_n230));
  INV_X1    g044(.A(G104), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G107), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n227), .A4(G104), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n229), .A2(new_n230), .A3(new_n232), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT82), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n235), .A2(new_n232), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT82), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n238), .A2(new_n239), .A3(new_n230), .A4(new_n229), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n238), .A2(new_n229), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(G101), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n230), .B1(new_n238), .B2(new_n229), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G119), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT68), .B(G116), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G119), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT2), .B(G113), .Z(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(KEYINPUT68), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G116), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n253), .A2(new_n255), .A3(G119), .ZN(new_n256));
  INV_X1    g070(.A(new_n248), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n251), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n242), .A2(new_n246), .B1(new_n252), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n245), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G110), .B(G122), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n230), .B1(new_n228), .B2(new_n232), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(new_n237), .B2(new_n240), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n266));
  INV_X1    g080(.A(G113), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n267), .B1(new_n248), .B2(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n266), .A2(new_n269), .B1(new_n250), .B2(new_n251), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n262), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT86), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n245), .A2(new_n261), .B1(new_n265), .B2(new_n270), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(new_n263), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n226), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n263), .B(KEYINPUT8), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n265), .A2(new_n270), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n279), .A2(KEYINPUT88), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n269), .B(KEYINPUT87), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n266), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n265), .A2(new_n282), .A3(new_n252), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n279), .B2(KEYINPUT88), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n278), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(G902), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT89), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n274), .A2(new_n263), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT6), .ZN(new_n291));
  INV_X1    g105(.A(new_n290), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n272), .A2(KEYINPUT86), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n275), .B1(new_n274), .B2(new_n263), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n291), .B1(new_n295), .B2(KEYINPUT6), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n220), .B(new_n222), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n286), .B(new_n289), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n291), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n290), .B1(new_n273), .B2(new_n276), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT6), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n297), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n289), .B1(new_n305), .B2(new_n286), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n187), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(G237), .A2(G953), .ZN(new_n308));
  AOI21_X1  g122(.A(G143), .B1(new_n308), .B2(G214), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(G143), .A3(G214), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT18), .ZN(new_n312));
  INV_X1    g126(.A(G131), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n310), .B(new_n311), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n311), .ZN(new_n315));
  OAI211_X1 g129(.A(KEYINPUT18), .B(G131), .C1(new_n315), .C2(new_n309), .ZN(new_n316));
  INV_X1    g130(.A(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n209), .A2(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G146), .ZN(new_n321));
  XNOR2_X1  g135(.A(G125), .B(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n188), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n314), .A2(new_n316), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT91), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT90), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT19), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n322), .A2(new_n327), .A3(KEYINPUT19), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n326), .B1(new_n332), .B2(new_n188), .ZN(new_n333));
  AOI211_X1 g147(.A(KEYINPUT91), .B(G146), .C1(new_n330), .C2(new_n331), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G131), .B1(new_n315), .B2(new_n309), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n310), .A2(new_n313), .A3(new_n311), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT16), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n317), .A3(G125), .ZN(new_n340));
  OAI211_X1 g154(.A(G146), .B(new_n340), .C1(new_n320), .C2(new_n339), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n325), .B1(new_n335), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT92), .ZN(new_n344));
  INV_X1    g158(.A(G122), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G113), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n267), .A2(G122), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n347), .A3(new_n344), .ZN(new_n350));
  AOI21_X1  g164(.A(G104), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n350), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n352), .A2(new_n348), .A3(new_n231), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT17), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n336), .A2(new_n337), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n340), .B1(new_n320), .B2(new_n339), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n188), .ZN(new_n360));
  OAI211_X1 g174(.A(KEYINPUT17), .B(G131), .C1(new_n315), .C2(new_n309), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(new_n341), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n354), .B(new_n325), .C1(new_n358), .C2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT93), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n357), .A2(new_n360), .A3(new_n341), .A4(new_n361), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n366), .A2(KEYINPUT93), .A3(new_n325), .A4(new_n354), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n343), .A2(new_n355), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(G475), .A2(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT20), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n367), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n332), .A2(new_n188), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT91), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n332), .A2(new_n326), .A3(new_n188), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n342), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n325), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n355), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT20), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n369), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n366), .A2(new_n325), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n355), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n372), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G902), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g200(.A(KEYINPUT94), .B(G475), .Z(new_n387));
  AOI22_X1  g201(.A1(new_n371), .A2(new_n381), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(G234), .A2(G237), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n389), .A2(G952), .A3(new_n221), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(G902), .A3(G953), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n391), .B(KEYINPUT96), .Z(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT21), .B(G898), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT9), .B(G234), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n396), .A2(new_n397), .A3(G953), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n249), .A2(G122), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n345), .A2(G116), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G107), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n227), .A3(new_n400), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n190), .A2(G128), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n195), .A2(G143), .ZN(new_n406));
  INV_X1    g220(.A(G134), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT13), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n406), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT95), .ZN(new_n411));
  INV_X1    g225(.A(new_n405), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(KEYINPUT13), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n405), .A2(KEYINPUT95), .A3(new_n409), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n404), .B(new_n408), .C1(new_n407), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n405), .A2(new_n406), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G134), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n408), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n399), .A2(new_n420), .A3(new_n400), .ZN(new_n421));
  OAI21_X1  g235(.A(G107), .B1(new_n399), .B2(new_n420), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n403), .B(new_n419), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n398), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n402), .A2(new_n403), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n408), .B1(new_n415), .B2(new_n407), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n423), .B(new_n398), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n385), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G478), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(KEYINPUT15), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OAI221_X1 g246(.A(new_n385), .B1(KEYINPUT15), .B2(new_n430), .C1(new_n424), .C2(new_n428), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n388), .A2(new_n395), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n307), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT26), .B(G101), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n308), .A2(G210), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n252), .A2(new_n260), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT69), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n218), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n215), .A2(KEYINPUT69), .A3(new_n217), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT11), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n407), .B2(G137), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n407), .A2(G137), .ZN(new_n451));
  INV_X1    g265(.A(G137), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT11), .A3(G134), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G131), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n450), .A2(new_n453), .A3(new_n313), .A4(new_n451), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT65), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT65), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n454), .A2(new_n458), .A3(G131), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n451), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n407), .A2(G137), .ZN(new_n462));
  OAI21_X1  g276(.A(G131), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n456), .ZN(new_n464));
  OAI22_X1  g278(.A1(new_n448), .A2(new_n460), .B1(new_n208), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n444), .B1(new_n465), .B2(KEYINPUT72), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n456), .A2(KEYINPUT65), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n455), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n215), .A2(KEYINPUT69), .A3(new_n217), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT69), .B1(new_n215), .B2(new_n217), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n205), .A2(new_n207), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n198), .A2(new_n199), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n198), .A2(new_n199), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n464), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n468), .A2(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT72), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n466), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT28), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n475), .A2(new_n476), .ZN(new_n483));
  INV_X1    g297(.A(new_n444), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n446), .A2(new_n457), .A3(new_n447), .A4(new_n459), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n218), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n457), .A2(new_n488), .A3(new_n459), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n484), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT28), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n443), .B1(new_n482), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n443), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n465), .A2(KEYINPUT30), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT30), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n489), .B(new_n496), .C1(new_n208), .C2(new_n464), .ZN(new_n497));
  AOI211_X1 g311(.A(KEYINPUT70), .B(new_n484), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT70), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n477), .B2(new_n496), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(new_n444), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n494), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT31), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n497), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n496), .B1(new_n483), .B2(new_n485), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n444), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n500), .A2(new_n499), .A3(new_n444), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT31), .A3(new_n494), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n492), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(G472), .A2(G902), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT73), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT32), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT75), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n515), .B1(new_n512), .B2(new_n514), .ZN(new_n519));
  INV_X1    g333(.A(new_n492), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT31), .B1(new_n510), .B2(new_n494), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n503), .B(new_n493), .C1(new_n508), .C2(new_n509), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n516), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT74), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT28), .B1(new_n466), .B2(new_n479), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n465), .A2(new_n444), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n481), .B1(new_n528), .B2(new_n486), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT29), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n442), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n527), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n526), .B1(new_n533), .B2(G902), .ZN(new_n534));
  INV_X1    g348(.A(new_n529), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n482), .A2(new_n535), .A3(new_n531), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(KEYINPUT74), .A3(new_n385), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n443), .B1(new_n510), .B2(new_n486), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n482), .A2(new_n491), .A3(new_n443), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n530), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n534), .B(new_n537), .C1(new_n538), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G472), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n518), .A2(new_n519), .A3(new_n525), .A4(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G221), .B1(new_n396), .B2(G902), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G469), .ZN(new_n546));
  XNOR2_X1  g360(.A(G110), .B(G140), .ZN(new_n547));
  INV_X1    g361(.A(G227), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(G953), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n547), .B(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n194), .A2(new_n191), .A3(new_n189), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n201), .A2(G128), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n473), .B2(new_n474), .ZN(new_n554));
  INV_X1    g368(.A(new_n264), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n241), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n229), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n235), .A2(new_n232), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n242), .B(G101), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n446), .A2(new_n447), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n245), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n197), .A2(new_n200), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n557), .B1(new_n564), .B2(new_n472), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n265), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n558), .A2(new_n563), .A3(new_n460), .A4(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT83), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n562), .A2(new_n245), .B1(new_n565), .B2(new_n265), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n570), .A2(KEYINPUT83), .A3(new_n460), .A4(new_n558), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n550), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n556), .B1(new_n265), .B2(new_n475), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n468), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n550), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT84), .ZN(new_n579));
  AND4_X1   g393(.A1(new_n579), .A2(new_n558), .A3(new_n566), .A4(new_n563), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n579), .B1(new_n570), .B2(new_n558), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n468), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n569), .A2(new_n571), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT85), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n577), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI211_X1 g400(.A(KEYINPUT85), .B(new_n578), .C1(new_n582), .C2(new_n583), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n546), .B(new_n385), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n576), .A2(new_n583), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n589), .A2(new_n550), .B1(new_n582), .B2(new_n572), .ZN(new_n590));
  OAI21_X1  g404(.A(G469), .B1(new_n590), .B2(G902), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n545), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n397), .B1(G234), .B2(new_n385), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n360), .A2(new_n341), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT76), .B1(new_n195), .B2(G119), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n195), .A2(KEYINPUT76), .A3(G119), .ZN(new_n597));
  INV_X1    g411(.A(G119), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G128), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT24), .B(G110), .Z(new_n602));
  NAND3_X1  g416(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n598), .A2(G128), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n599), .B(new_n603), .C1(new_n604), .C2(KEYINPUT23), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n601), .A2(new_n602), .B1(new_n605), .B2(G110), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n595), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n341), .A2(new_n323), .ZN(new_n608));
  OAI22_X1  g422(.A1(new_n601), .A2(new_n602), .B1(new_n605), .B2(G110), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT77), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT22), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G137), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT77), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n607), .A2(new_n610), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n612), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n607), .A2(new_n610), .A3(new_n615), .A4(KEYINPUT78), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT78), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n611), .B2(new_n616), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n619), .A2(new_n385), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n594), .B1(new_n623), .B2(KEYINPUT25), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n622), .A2(new_n620), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT25), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n625), .A2(new_n626), .A3(new_n385), .A4(new_n619), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT79), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT79), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n624), .A2(new_n630), .A3(new_n627), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n593), .A2(G902), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT80), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n625), .A2(new_n619), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n629), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n437), .A2(new_n543), .A3(new_n592), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT97), .B(G101), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G3));
  INV_X1    g453(.A(G472), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n523), .A2(new_n385), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n504), .A2(new_n511), .ZN(new_n644));
  AOI21_X1  g458(.A(G902), .B1(new_n644), .B2(new_n520), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT98), .ZN(new_n646));
  INV_X1    g460(.A(new_n514), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n643), .A2(new_n646), .B1(new_n523), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n592), .A3(new_n636), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n286), .B(new_n287), .C1(new_n296), .C2(new_n297), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n287), .B1(new_n305), .B2(new_n286), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n187), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n386), .A2(new_n387), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n380), .B1(new_n379), .B2(new_n369), .ZN(new_n655));
  AOI211_X1 g469(.A(KEYINPUT20), .B(new_n370), .C1(new_n372), .C2(new_n378), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n658), .B1(new_n424), .B2(new_n428), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n660));
  INV_X1    g474(.A(new_n398), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(KEYINPUT33), .A3(new_n427), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n659), .A2(G478), .A3(new_n663), .A4(new_n385), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n429), .A2(new_n430), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n657), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n653), .A2(new_n394), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n649), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT34), .B(G104), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n654), .B(new_n434), .C1(new_n655), .C2(new_n656), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n674), .B1(new_n675), .B2(new_n394), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n388), .A2(KEYINPUT99), .A3(new_n395), .A4(new_n434), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n673), .B1(new_n653), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n187), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n286), .B1(new_n296), .B2(new_n297), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n288), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n680), .B1(new_n682), .B2(new_n650), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(KEYINPUT100), .A3(new_n676), .A4(new_n677), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n649), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT35), .B(G107), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G9));
  AND3_X1   g502(.A1(new_n624), .A2(new_n630), .A3(new_n627), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n630), .B1(new_n624), .B2(new_n627), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n616), .A2(KEYINPUT36), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n612), .A2(new_n618), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n691), .B1(new_n612), .B2(new_n618), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n633), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(KEYINPUT101), .B(new_n633), .C1(new_n692), .C2(new_n693), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n689), .A2(new_n690), .A3(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n307), .A2(new_n436), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n648), .A2(new_n592), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT37), .B(G110), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G12));
  NAND4_X1  g517(.A1(new_n629), .A2(new_n631), .A3(new_n696), .A4(new_n697), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n704), .B(new_n187), .C1(new_n652), .C2(new_n651), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n512), .A2(KEYINPUT75), .A3(new_n517), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n524), .B1(new_n523), .B2(new_n516), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n523), .A2(new_n647), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n709), .A2(new_n515), .B1(G472), .B2(new_n541), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n705), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(G900), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n390), .B1(new_n392), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n675), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n545), .B(new_n715), .C1(new_n588), .C2(new_n591), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT102), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n195), .ZN(G30));
  XOR2_X1   g533(.A(new_n713), .B(KEYINPUT39), .Z(new_n720));
  NAND2_X1  g534(.A1(new_n592), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n721), .B(KEYINPUT40), .Z(new_n722));
  INV_X1    g536(.A(new_n502), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n443), .B1(new_n528), .B2(new_n486), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n385), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n709), .A2(new_n515), .B1(G472), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n708), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n299), .A2(new_n306), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT38), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n388), .A2(new_n435), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n699), .A2(new_n187), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n722), .A2(new_n727), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT103), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n190), .ZN(G45));
  INV_X1    g548(.A(new_n713), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n657), .A2(new_n666), .A3(new_n735), .ZN(new_n736));
  AOI211_X1 g550(.A(new_n545), .B(new_n736), .C1(new_n588), .C2(new_n591), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n711), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G146), .ZN(G48));
  INV_X1    g553(.A(new_n588), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n558), .A2(new_n566), .A3(new_n563), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT84), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n570), .A2(new_n579), .A3(new_n558), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n744), .A2(new_n468), .B1(new_n569), .B2(new_n571), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT85), .B1(new_n745), .B2(new_n578), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n584), .A2(new_n585), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n577), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n546), .B1(new_n748), .B2(new_n385), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n740), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n544), .A3(new_n543), .A4(new_n636), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n669), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT41), .B(G113), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G15));
  NOR2_X1   g568(.A1(new_n685), .A2(new_n751), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n247), .ZN(G18));
  NOR2_X1   g570(.A1(new_n699), .A2(new_n436), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n543), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n385), .B1(new_n586), .B2(new_n587), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(G469), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n683), .A3(new_n544), .A4(new_n588), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G119), .ZN(G21));
  OAI21_X1  g579(.A(new_n442), .B1(new_n527), .B2(new_n529), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n766), .B1(new_n521), .B2(new_n522), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n641), .A2(G472), .B1(new_n647), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n636), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n683), .A2(new_n395), .A3(new_n730), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n761), .A2(new_n588), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n545), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  NOR2_X1   g589(.A1(new_n762), .A2(new_n736), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n767), .A2(new_n647), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n704), .B(new_n777), .C1(new_n645), .C2(new_n640), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT104), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n641), .A2(G472), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(KEYINPUT104), .A3(new_n704), .A4(new_n777), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n776), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G125), .ZN(G27));
  NAND2_X1  g599(.A1(G469), .A2(G902), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT105), .Z(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n590), .B2(G469), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n545), .B1(new_n588), .B2(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n299), .A2(new_n306), .A3(new_n680), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n543), .A2(new_n789), .A3(new_n636), .A4(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT106), .B1(new_n791), .B2(new_n736), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT42), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n635), .B1(new_n708), .B2(new_n710), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n588), .A2(new_n788), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n795), .A2(new_n790), .A3(new_n544), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT106), .ZN(new_n797));
  INV_X1    g611(.A(new_n736), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n794), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n792), .A2(new_n793), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n523), .A2(new_n516), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n635), .B1(new_n710), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n796), .A2(new_n802), .A3(KEYINPUT42), .A4(new_n798), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G131), .ZN(G33));
  NAND3_X1  g619(.A1(new_n794), .A2(new_n796), .A3(new_n714), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G134), .ZN(G36));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT107), .ZN(new_n809));
  XOR2_X1   g623(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n810));
  NAND2_X1  g624(.A1(new_n388), .A2(new_n666), .ZN(new_n811));
  MUX2_X1   g625(.A(new_n809), .B(new_n810), .S(new_n811), .Z(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n704), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n648), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n814), .A2(KEYINPUT44), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(KEYINPUT44), .ZN(new_n816));
  INV_X1    g630(.A(new_n790), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n590), .A2(KEYINPUT45), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n546), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n590), .A2(KEYINPUT45), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n787), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT46), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n822), .A2(KEYINPUT46), .A3(new_n823), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n588), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n544), .A3(new_n720), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n818), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT108), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(new_n452), .ZN(G39));
  INV_X1    g647(.A(KEYINPUT47), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(new_n834), .A3(new_n544), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n834), .B1(new_n828), .B2(new_n544), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n543), .A2(new_n817), .A3(new_n636), .A4(new_n736), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(G140), .ZN(G42));
  NOR4_X1   g655(.A1(new_n635), .A2(new_n545), .A3(new_n811), .A4(new_n680), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT109), .Z(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(KEYINPUT49), .B2(new_n772), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT110), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n729), .A2(new_n727), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n845), .B(new_n846), .C1(KEYINPUT49), .C2(new_n772), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n544), .A2(new_n750), .A3(new_n390), .A4(new_n790), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n848), .A2(new_n812), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(new_n802), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n850), .A2(KEYINPUT48), .ZN(new_n851));
  INV_X1    g665(.A(new_n727), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n848), .A2(new_n636), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n667), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n640), .B1(new_n523), .B2(new_n385), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n514), .B1(new_n644), .B2(new_n766), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n856), .A2(new_n857), .A3(new_n635), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n812), .A3(new_n390), .ZN(new_n859));
  OAI211_X1 g673(.A(G952), .B(new_n221), .C1(new_n859), .C2(new_n762), .ZN(new_n860));
  OR3_X1    g674(.A1(new_n854), .A2(new_n855), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n855), .B1(new_n854), .B2(new_n860), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n850), .A2(KEYINPUT48), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n851), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n849), .A2(new_n783), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n388), .A2(new_n665), .A3(new_n664), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n866), .B1(new_n853), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n859), .A2(new_n817), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n750), .A2(new_n545), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n836), .B2(new_n837), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n865), .B(new_n868), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n729), .A2(new_n859), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n773), .A2(KEYINPUT114), .A3(new_n680), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT114), .B1(new_n773), .B2(new_n680), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT50), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n873), .B(KEYINPUT50), .C1(new_n876), .C2(new_n877), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n864), .B1(new_n872), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT116), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n870), .B(KEYINPUT113), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n836), .B2(new_n837), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n868), .B1(new_n886), .B2(new_n869), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n882), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n884), .B1(new_n888), .B2(new_n865), .ZN(new_n889));
  AOI211_X1 g703(.A(KEYINPUT116), .B(KEYINPUT51), .C1(new_n887), .C2(new_n882), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n667), .A2(new_n675), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n307), .A2(new_n894), .A3(new_n394), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n648), .A2(new_n592), .A3(new_n895), .A4(new_n636), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n806), .A2(new_n896), .A3(new_n701), .A4(new_n637), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n545), .B(new_n736), .C1(new_n588), .C2(new_n788), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT104), .B1(new_n768), .B2(new_n704), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n856), .A2(new_n857), .A3(new_n699), .A4(new_n779), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR4_X1   g715(.A1(new_n699), .A2(new_n434), .A3(new_n657), .A4(new_n713), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n543), .A2(new_n902), .A3(new_n592), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n817), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT111), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n751), .B1(new_n685), .B2(new_n669), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n858), .A2(new_n395), .A3(new_n683), .A4(new_n730), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n750), .A2(new_n544), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n908), .A2(new_n909), .B1(new_n758), .B2(new_n762), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n906), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n763), .A2(new_n759), .B1(new_n771), .B2(new_n773), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n679), .A2(new_n684), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n794), .B(new_n773), .C1(new_n913), .C2(new_n668), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(KEYINPUT111), .A3(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n905), .A2(new_n804), .A3(new_n911), .A4(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n711), .B1(new_n716), .B2(new_n737), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n683), .A2(new_n730), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n704), .A2(new_n713), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n727), .A2(new_n789), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n784), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT52), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n784), .A2(new_n917), .A3(KEYINPUT52), .A4(new_n920), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n926));
  OR3_X1    g740(.A1(new_n916), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT53), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n916), .B2(new_n925), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n892), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n926), .B1(new_n916), .B2(new_n925), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n923), .A2(new_n924), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n907), .A2(new_n910), .A3(new_n928), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n932), .A2(new_n804), .A3(new_n905), .A4(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n931), .A2(new_n892), .A3(new_n934), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n891), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(G952), .A2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n847), .B1(new_n936), .B2(new_n937), .ZN(G75));
  NAND2_X1  g752(.A1(new_n296), .A2(new_n297), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n305), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n385), .B1(new_n931), .B2(new_n934), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n943), .A2(G210), .ZN(new_n944));
  OR2_X1    g758(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n221), .A2(G952), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n944), .A2(new_n945), .A3(new_n942), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(G51));
  AOI211_X1 g765(.A(new_n385), .B(new_n822), .C1(new_n931), .C2(new_n934), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n787), .B(KEYINPUT57), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n892), .B1(new_n931), .B2(new_n934), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n935), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n955), .B2(new_n748), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT120), .B1(new_n956), .B2(new_n947), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT120), .ZN(new_n958));
  INV_X1    g772(.A(new_n748), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n931), .A2(new_n934), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT54), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n931), .A2(new_n892), .A3(new_n934), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n959), .B1(new_n963), .B2(new_n953), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n958), .B(new_n948), .C1(new_n964), .C2(new_n952), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n957), .A2(new_n965), .ZN(G54));
  AND2_X1   g780(.A1(KEYINPUT58), .A2(G475), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n943), .A2(new_n379), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n968), .A2(KEYINPUT121), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(KEYINPUT121), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n379), .B1(new_n943), .B2(new_n967), .ZN(new_n971));
  NOR4_X1   g785(.A1(new_n969), .A2(new_n970), .A3(new_n947), .A4(new_n971), .ZN(G60));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT59), .Z(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n930), .B2(new_n935), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n659), .A2(new_n663), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(KEYINPUT122), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n974), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n947), .B1(new_n963), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT122), .B1(new_n976), .B2(new_n977), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(G63));
  NAND2_X1  g797(.A1(G217), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT60), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n931), .B2(new_n934), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n625), .A2(new_n619), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT124), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n947), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n692), .A2(new_n693), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n986), .A2(KEYINPUT123), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT123), .B1(new_n986), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n990), .B(KEYINPUT61), .C1(new_n992), .C2(new_n993), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(G66));
  AND3_X1   g812(.A1(new_n896), .A2(new_n637), .A3(new_n701), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n911), .A2(new_n915), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G224), .A2(G953), .ZN(new_n1001));
  OAI22_X1  g815(.A1(new_n1000), .A2(G953), .B1(new_n393), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n296), .B1(G898), .B2(new_n221), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1002), .B(new_n1003), .Z(G69));
  XOR2_X1   g818(.A(new_n500), .B(new_n332), .Z(new_n1005));
  NAND2_X1  g819(.A1(new_n802), .A2(new_n918), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n806), .B1(new_n829), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(new_n818), .B2(new_n830), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n784), .A2(new_n917), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(KEYINPUT125), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(KEYINPUT125), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1008), .A2(new_n840), .A3(new_n804), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n221), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n548), .A2(G900), .A3(G953), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1005), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n733), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n1012), .ZN(new_n1018));
  AOI22_X1  g832(.A1(new_n1018), .A2(KEYINPUT62), .B1(new_n838), .B2(new_n839), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n794), .A2(new_n790), .A3(new_n893), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n831), .B1(new_n721), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(G953), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT126), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n733), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT62), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND4_X1   g840(.A1(new_n1023), .A2(new_n1017), .A3(new_n1025), .A4(new_n1012), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1019), .B(new_n1022), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1016), .B1(new_n1030), .B2(new_n1005), .ZN(G72));
  NAND2_X1  g845(.A1(G472), .A2(G902), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1032), .B(KEYINPUT63), .Z(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(new_n1013), .B2(new_n1000), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n510), .A2(new_n486), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT127), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1034), .A2(new_n442), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n927), .A2(new_n929), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n1039), .B(new_n1033), .C1(new_n723), .C2(new_n538), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1038), .A2(new_n1040), .A3(new_n948), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1021), .A2(new_n1000), .ZN(new_n1042));
  OAI211_X1 g856(.A(new_n1019), .B(new_n1042), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n1033), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1037), .A2(new_n442), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(G57));
endmodule


