//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n550, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G219), .A3(G221), .A4(G220), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(new_n464), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(G2105), .B2(new_n471), .ZN(G160));
  INV_X1    g047(.A(new_n469), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n476), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND4_X1  g059(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n477), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(G2105), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n461), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(new_n477), .B2(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n494), .A2(KEYINPUT68), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n488), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n487), .A2(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT70), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT71), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(new_n500), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G62), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n499), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT72), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n505), .A2(new_n509), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n503), .B1(new_n515), .B2(new_n516), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT69), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n514), .A2(new_n519), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n518), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n501), .A2(new_n504), .B1(new_n506), .B2(new_n508), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n529), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n520), .A2(G51), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n526), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(new_n520), .A2(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n529), .A2(new_n517), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT74), .B(G90), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT73), .Z(new_n539));
  AOI21_X1  g114(.A(new_n537), .B1(new_n539), .B2(G651), .ZN(G171));
  AOI22_X1  g115(.A1(new_n529), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n520), .A2(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n535), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G188));
  XOR2_X1   g129(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n520), .B2(G53), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT78), .B(G65), .Z(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n510), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n556), .B1(new_n559), .B2(G651), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n520), .A2(new_n561), .A3(KEYINPUT9), .A4(G53), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n505), .A2(new_n509), .A3(G91), .A4(new_n517), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n529), .A2(KEYINPUT77), .A3(G91), .A4(new_n517), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n560), .A2(new_n562), .A3(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n510), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(G49), .B2(new_n520), .ZN(new_n572));
  INV_X1    g147(.A(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n573), .B2(new_n535), .ZN(G288));
  AOI22_X1  g149(.A1(new_n529), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n529), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n576));
  INV_X1    g151(.A(new_n517), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n542), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n518), .A2(G85), .B1(G47), .B2(new_n520), .ZN(new_n579));
  NAND2_X1  g154(.A1(G72), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n510), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n579), .B1(new_n583), .B2(new_n542), .ZN(G290));
  NAND2_X1  g159(.A1(new_n518), .A2(G92), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n520), .A2(G54), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n529), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n542), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n592), .B2(G171), .ZN(G284));
  OAI21_X1  g169(.A(new_n593), .B1(new_n592), .B2(G171), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n560), .A2(new_n562), .A3(new_n567), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  XOR2_X1   g173(.A(G280), .B(KEYINPUT79), .Z(G297));
  AND3_X1   g174(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n600));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n475), .A2(G123), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n479), .A2(G135), .ZN(new_n608));
  NOR2_X1   g183(.A1(G99), .A2(G2105), .ZN(new_n609));
  OAI21_X1  g184(.A(G2104), .B1(new_n477), .B2(G111), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND3_X1  g187(.A1(new_n477), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT13), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(G156));
  XNOR2_X1  g192(.A(G2427), .B(G2438), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2430), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT15), .B(G2435), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT14), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2443), .B(G2446), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n624), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(G14), .A3(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g209(.A1(new_n630), .A2(KEYINPUT81), .A3(G14), .A4(new_n631), .ZN(new_n635));
  AND2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(G401));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2067), .B(G2678), .Z(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT17), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(KEYINPUT18), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2072), .B(G2078), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n644), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT82), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XNOR2_X1  g226(.A(G1971), .B(G1976), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XOR2_X1   g228(.A(G1956), .B(G2474), .Z(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n658));
  INV_X1    g233(.A(new_n653), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  AOI22_X1  g235(.A1(new_n657), .A2(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n662), .A2(new_n653), .A3(new_n656), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n661), .B(new_n663), .C1(new_n657), .C2(new_n658), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1986), .B(G1996), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G1981), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1991), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G229));
  INV_X1    g245(.A(G29), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G26), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n475), .A2(G128), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n479), .A2(G140), .ZN(new_n674));
  OR2_X1    g249(.A1(G104), .A2(G2105), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n675), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n672), .B1(new_n678), .B2(new_n671), .ZN(new_n679));
  MUX2_X1   g254(.A(new_n672), .B(new_n679), .S(KEYINPUT28), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G2067), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT92), .B(G1341), .ZN(new_n682));
  INV_X1    g257(.A(G19), .ZN(new_n683));
  OAI21_X1  g258(.A(KEYINPUT91), .B1(new_n683), .B2(G16), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n683), .A2(KEYINPUT91), .A3(G16), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n684), .B(new_n685), .C1(new_n547), .C2(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n681), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n682), .B2(new_n687), .ZN(new_n689));
  NOR2_X1   g264(.A1(G4), .A2(G16), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n600), .B2(G16), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT90), .B(G1348), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n689), .B(new_n694), .C1(G2067), .C2(new_n680), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT93), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n671), .A2(G35), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G162), .B2(new_n671), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT29), .B(G2090), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G29), .A2(G32), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT26), .Z(new_n703));
  INV_X1    g278(.A(G129), .ZN(new_n704));
  INV_X1    g279(.A(G141), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n703), .B1(new_n474), .B2(new_n704), .C1(new_n705), .C2(new_n478), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT96), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n477), .A2(G105), .A3(G2104), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT95), .Z(new_n709));
  OR3_X1    g284(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n707), .B1(new_n706), .B2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n701), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT27), .B(G1996), .Z(new_n715));
  OAI21_X1  g290(.A(new_n700), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n671), .A2(G27), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G164), .B2(new_n671), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n714), .A2(new_n715), .B1(G2078), .B2(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n671), .A2(G33), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT25), .Z(new_n722));
  INV_X1    g297(.A(G139), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n722), .B1(new_n478), .B2(new_n723), .C1(new_n724), .C2(new_n477), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n720), .B1(new_n725), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(G2072), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(KEYINPUT24), .A2(G34), .ZN(new_n729));
  NAND2_X1  g304(.A1(KEYINPUT24), .A2(G34), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n729), .A2(new_n671), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G160), .B2(new_n671), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G2084), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT94), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n726), .A2(new_n727), .B1(new_n732), .B2(G2084), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n719), .A2(new_n728), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  NAND2_X1  g313(.A1(G171), .A2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G5), .B2(G16), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n716), .B(new_n737), .C1(new_n738), .C2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G2078), .B2(new_n718), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT99), .B(KEYINPUT23), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n686), .A2(G20), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n597), .B2(new_n686), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT100), .ZN(new_n747));
  INV_X1    g322(.A(G1956), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n696), .A2(new_n742), .A3(new_n749), .ZN(new_n750));
  MUX2_X1   g325(.A(G24), .B(G290), .S(G16), .Z(new_n751));
  AOI22_X1  g326(.A1(new_n751), .A2(G1986), .B1(KEYINPUT89), .B2(KEYINPUT36), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G1986), .B2(new_n751), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n686), .A2(G23), .ZN(new_n754));
  INV_X1    g329(.A(G288), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(new_n686), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT87), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT33), .B(G1976), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  MUX2_X1   g334(.A(G6), .B(G305), .S(G16), .Z(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT32), .B(G1981), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n686), .A2(G22), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G166), .B2(new_n686), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n762), .B1(new_n764), .B2(G1971), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n759), .B(new_n765), .C1(G1971), .C2(new_n764), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n753), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n671), .A2(G25), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n475), .A2(G119), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT84), .Z(new_n771));
  OR2_X1    g346(.A1(G95), .A2(G2105), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n772), .B(G2104), .C1(G107), .C2(new_n477), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n479), .A2(G131), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n769), .B1(new_n776), .B2(new_n671), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT35), .B(G1991), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT85), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n777), .B(new_n779), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n768), .B(new_n780), .C1(new_n767), .C2(new_n766), .ZN(new_n781));
  AOI21_X1  g356(.A(KEYINPUT89), .B1(KEYINPUT88), .B2(KEYINPUT36), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(G168), .A2(G16), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G16), .B2(G21), .ZN(new_n785));
  INV_X1    g360(.A(G1966), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT97), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT31), .B(G11), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n740), .A2(new_n738), .ZN(new_n790));
  INV_X1    g365(.A(G28), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n791), .B2(KEYINPUT30), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(KEYINPUT30), .B2(new_n791), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n611), .B2(new_n671), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n785), .B2(new_n786), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n788), .A2(new_n789), .A3(new_n790), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT98), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n781), .A2(new_n782), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n750), .A2(new_n783), .A3(new_n797), .A4(new_n798), .ZN(G150));
  INV_X1    g374(.A(G150), .ZN(G311));
  INV_X1    g375(.A(G860), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT39), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n600), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT102), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n542), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n520), .A2(G55), .ZN(new_n809));
  INV_X1    g384(.A(G93), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n535), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(new_n547), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n543), .A2(new_n546), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(new_n812), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n806), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n806), .A2(new_n818), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n804), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n821), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n823), .A2(new_n819), .A3(new_n803), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n802), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n801), .B1(new_n825), .B2(KEYINPUT103), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n822), .A2(new_n824), .A3(new_n802), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT103), .ZN(new_n828));
  AOI211_X1 g403(.A(new_n828), .B(new_n802), .C1(new_n822), .C2(new_n824), .ZN(new_n829));
  OR3_X1    g404(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT104), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n813), .A2(G860), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT37), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT104), .B1(new_n836), .B2(new_n833), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(G145));
  XNOR2_X1  g413(.A(new_n611), .B(G160), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n483), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT106), .ZN(new_n841));
  INV_X1    g416(.A(new_n614), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n840), .A2(KEYINPUT106), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(KEYINPUT106), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(new_n614), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n713), .A2(new_n677), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n475), .A2(G130), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n479), .A2(G142), .ZN(new_n850));
  OR2_X1    g425(.A1(G106), .A2(G2105), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n851), .B(G2104), .C1(G118), .C2(new_n477), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n677), .B1(new_n710), .B2(new_n711), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n848), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n712), .A2(new_n678), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n853), .B1(new_n858), .B2(new_n855), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n859), .A3(new_n775), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n775), .B1(new_n857), .B2(new_n859), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n485), .B(KEYINPUT4), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT68), .B1(new_n494), .B2(new_n495), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n490), .A2(G2105), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n492), .A2(new_n865), .A3(new_n489), .A4(G2104), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n867), .A2(new_n868), .A3(new_n488), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n868), .B1(new_n867), .B2(new_n488), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n863), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n725), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n861), .A2(new_n862), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n857), .A2(new_n859), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n776), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n872), .B1(new_n876), .B2(new_n860), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n847), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n873), .B1(new_n861), .B2(new_n862), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n872), .A3(new_n860), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n846), .A4(new_n843), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(G395));
  XNOR2_X1  g460(.A(G288), .B(G305), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G290), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n887), .A2(G303), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(G303), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n818), .B(new_n603), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(G299), .A2(KEYINPUT108), .ZN(new_n895));
  NAND2_X1  g470(.A1(G299), .A2(KEYINPUT108), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n600), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n591), .A2(KEYINPUT108), .A3(G299), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n900));
  AND2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n899), .A2(KEYINPUT41), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n894), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n893), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n888), .A2(KEYINPUT42), .A3(new_n889), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n892), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n888), .A2(KEYINPUT42), .A3(new_n889), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT42), .B1(new_n888), .B2(new_n889), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n903), .B(new_n905), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n911), .A3(G868), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n813), .A2(new_n592), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT110), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT111), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n918), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n917), .B1(new_n912), .B2(new_n913), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT111), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n919), .A2(new_n922), .ZN(G295));
  NAND2_X1  g498(.A1(new_n915), .A2(new_n918), .ZN(G331));
  NAND2_X1  g499(.A1(new_n904), .A2(new_n900), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n899), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n818), .A2(G301), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n817), .A2(G171), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(G168), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(G168), .B1(new_n928), .B2(new_n929), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n925), .B(new_n927), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n929), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G286), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n904), .A3(new_n930), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n890), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  OAI22_X1  g514(.A1(new_n931), .A2(new_n932), .B1(new_n901), .B2(new_n902), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n890), .A3(new_n936), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n938), .A2(new_n939), .A3(new_n882), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n882), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n890), .B1(new_n940), .B2(new_n936), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT43), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n943), .A2(new_n944), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n938), .A2(KEYINPUT112), .A3(new_n882), .A4(new_n941), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n943), .B2(new_n937), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n950), .B1(new_n954), .B2(KEYINPUT43), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n948), .B1(new_n955), .B2(new_n947), .ZN(G397));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n871), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(KEYINPUT113), .B(KEYINPUT45), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(G160), .A2(G40), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n775), .A2(new_n778), .ZN(new_n965));
  INV_X1    g540(.A(G2067), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n677), .B(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n713), .A2(G1996), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n712), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n965), .B(new_n967), .C1(new_n968), .C2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n678), .A2(new_n966), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n964), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n964), .B1(new_n713), .B2(new_n967), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n963), .A2(KEYINPUT46), .A3(new_n969), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT46), .B1(new_n963), .B2(new_n969), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT47), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n967), .B1(new_n968), .B2(new_n970), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n775), .A2(new_n778), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n979), .A2(new_n980), .A3(new_n965), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n963), .ZN(new_n983));
  OR2_X1    g558(.A1(G290), .A2(G1986), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n964), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT48), .Z(new_n986));
  AOI211_X1 g561(.A(new_n973), .B(new_n978), .C1(new_n983), .C2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(G166), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n988), .A2(new_n989), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n871), .A2(KEYINPUT45), .A3(new_n957), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n957), .B1(new_n487), .B2(new_n497), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n960), .ZN(new_n998));
  INV_X1    g573(.A(new_n467), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n471), .A2(G2105), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n999), .A2(new_n1000), .A3(G40), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1971), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n871), .A2(new_n1005), .A3(new_n957), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n962), .B1(new_n997), .B2(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1004), .B1(G2090), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n995), .B1(G8), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT63), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n995), .A2(G8), .A3(new_n1009), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G305), .B(G1981), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT49), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n497), .A2(KEYINPUT105), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n867), .A2(new_n868), .A3(new_n488), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1384), .B1(new_n1018), .B2(new_n863), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n992), .B1(new_n1019), .B2(new_n1001), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(G288), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n755), .A2(KEYINPUT115), .A3(G1976), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1020), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n755), .A2(G1976), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1026), .A2(KEYINPUT52), .A3(new_n1028), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1021), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT45), .B1(new_n871), .B2(new_n957), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1001), .B1(new_n997), .B2(new_n960), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n786), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2084), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1006), .A2(new_n1007), .A3(new_n1034), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n992), .B(G286), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1012), .A2(new_n1013), .A3(new_n1030), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1005), .B1(new_n871), .B2(new_n957), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT117), .B1(new_n1038), .B2(new_n962), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(new_n1001), .C1(new_n1019), .C2(new_n1005), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1043), .A2(G2090), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n992), .B1(new_n1044), .B2(new_n1004), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1030), .B(new_n1013), .C1(new_n1045), .C2(new_n995), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1036), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1011), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1037), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1030), .A2(G8), .A3(new_n995), .A4(new_n1009), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n755), .A2(new_n1023), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT116), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1015), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G305), .A2(G1981), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1020), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1049), .A2(new_n1050), .A3(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(G168), .A2(new_n992), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1036), .A2(KEYINPUT51), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1033), .A2(new_n1059), .A3(new_n1035), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1061));
  OAI21_X1  g636(.A(G8), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT123), .B(G8), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1057), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1058), .B1(new_n1067), .B2(KEYINPUT51), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT122), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1033), .A2(new_n1059), .A3(new_n1035), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1066), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT62), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1002), .B2(G2078), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT124), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1074), .A2(G2078), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1008), .A2(new_n738), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(new_n1074), .C1(new_n1002), .C2(G2078), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1076), .A2(new_n1079), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1072), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n992), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1057), .B1(new_n1092), .B2(KEYINPUT123), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n1093), .B2(new_n1064), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1089), .B(new_n1090), .C1(new_n1094), .C2(new_n1058), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1073), .A2(new_n1088), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1019), .A2(new_n1097), .A3(new_n966), .A4(new_n1001), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n871), .A2(new_n957), .A3(new_n966), .A4(new_n1001), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT119), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n692), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n591), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1105), .A2(new_n600), .A3(new_n1102), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT60), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n996), .A2(new_n969), .A3(new_n998), .A4(new_n1001), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n958), .B2(new_n962), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n815), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1111), .B(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1043), .A2(new_n748), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n597), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1120));
  NAND3_X1  g695(.A1(G299), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n996), .A2(new_n998), .A3(new_n1001), .A4(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1114), .A2(new_n1115), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  OR4_X1    g701(.A1(KEYINPUT60), .A2(new_n1105), .A3(new_n591), .A4(new_n1102), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1107), .A2(new_n1113), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n600), .B1(new_n1105), .B2(new_n1102), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1125), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1043), .B2(new_n748), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1131), .B2(new_n1123), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1123), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1122), .B(new_n1130), .C1(new_n1043), .C2(new_n748), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(new_n1115), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1133), .A2(KEYINPUT120), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1134), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT121), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1135), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n467), .A2(KEYINPUT126), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n467), .A2(KEYINPUT126), .ZN(new_n1148));
  AND4_X1   g723(.A1(G40), .A2(new_n961), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1149), .A2(new_n1000), .A3(new_n996), .A4(new_n1078), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1150), .A2(new_n1080), .A3(new_n1082), .A4(new_n1076), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(G171), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1146), .B1(new_n1088), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1090), .B1(new_n1094), .B2(new_n1058), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(G171), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1155), .B(KEYINPUT54), .C1(G171), .C2(new_n1083), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1096), .B1(new_n1145), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1046), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1056), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n982), .B1(G1986), .B2(G290), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n964), .B1(new_n1161), .B2(new_n984), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n987), .B1(new_n1160), .B2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g738(.A1(G229), .A2(new_n459), .ZN(new_n1165));
  INV_X1    g739(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1166), .B1(new_n942), .B2(new_n945), .ZN(new_n1167));
  AOI21_X1  g741(.A(G227), .B1(new_n634), .B2(new_n635), .ZN(new_n1168));
  AND2_X1   g742(.A1(new_n883), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1170));
  AND3_X1   g744(.A1(new_n1167), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1171), .A2(new_n1172), .ZN(G308));
  NAND2_X1  g747(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n1167), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1176), .ZN(G225));
endmodule


