//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(new_n202), .A2(new_n203), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n215), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n214), .B(new_n218), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G250), .B(G257), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT67), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n231), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n201), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n203), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n240), .B(new_n245), .Z(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT7), .B1(new_n247), .B2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT7), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(new_n254), .A3(new_n212), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n248), .A2(new_n255), .A3(G68), .ZN(new_n256));
  INV_X1    g0056(.A(G159), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n212), .A2(new_n249), .A3(KEYINPUT70), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT70), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G20), .B2(G33), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G58), .A2(G68), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n212), .B1(new_n208), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT16), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n211), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n261), .A2(new_n263), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n250), .A2(KEYINPUT81), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT81), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(new_n249), .A3(KEYINPUT3), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n252), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n254), .A2(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n251), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT68), .ZN(new_n283));
  AOI21_X1  g0083(.A(G20), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n278), .B1(new_n284), .B2(KEYINPUT7), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n272), .B1(new_n285), .B2(G68), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n270), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT72), .B1(new_n212), .B2(G1), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT72), .ZN(new_n290));
  INV_X1    g0090(.A(G1), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n267), .A2(new_n211), .ZN(new_n294));
  INV_X1    g0094(.A(G13), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G20), .ZN(new_n297));
  AND2_X1   g0097(.A1(KEYINPUT8), .A2(G58), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT8), .A2(G58), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n293), .A2(new_n294), .A3(new_n297), .A4(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT82), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT8), .B(G58), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n295), .A2(new_n212), .A3(G1), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n301), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n302), .B1(new_n301), .B2(new_n305), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n288), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G41), .ZN(new_n310));
  OAI211_X1 g0110(.A(G1), .B(G13), .C1(new_n249), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G1698), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n312), .A2(G226), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n247), .B(new_n313), .C1(G223), .C2(G1698), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G87), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n291), .B1(G41), .B2(G45), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(new_n311), .A3(G274), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n311), .A2(new_n317), .ZN(new_n320));
  INV_X1    g0120(.A(G232), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G179), .ZN(new_n324));
  OAI21_X1  g0124(.A(G169), .B1(new_n316), .B2(new_n322), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n309), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT18), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n288), .A2(new_n308), .B1(new_n325), .B2(new_n324), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT18), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(KEYINPUT83), .A2(G190), .ZN(new_n334));
  NOR2_X1   g0134(.A1(KEYINPUT83), .A2(G190), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n323), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(G200), .B2(new_n323), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n288), .A2(new_n338), .A3(new_n308), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT17), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n288), .A2(new_n338), .A3(KEYINPUT17), .A4(new_n308), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G244), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n319), .B1(new_n320), .B2(new_n345), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT68), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT68), .B1(new_n250), .B2(new_n252), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G238), .A2(G1698), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n321), .B2(G1698), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G107), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n349), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n311), .B1(new_n354), .B2(KEYINPUT73), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT73), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n352), .B(new_n356), .C1(new_n353), .C2(new_n349), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n346), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G179), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n293), .ZN(new_n362));
  INV_X1    g0162(.A(G77), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n304), .A2(new_n268), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(G77), .B2(new_n297), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n258), .A2(new_n260), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n303), .A2(KEYINPUT74), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n303), .A2(KEYINPUT74), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n249), .A2(G20), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(G20), .B2(G77), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n294), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n358), .B2(G169), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n361), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n364), .A2(new_n365), .B1(new_n363), .B2(new_n304), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n371), .A2(new_n375), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n294), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT75), .B1(new_n367), .B2(new_n376), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n354), .A2(KEYINPUT73), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n357), .ZN(new_n391));
  INV_X1    g0191(.A(new_n346), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(G190), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G200), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n388), .B(new_n393), .C1(new_n394), .C2(new_n358), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n333), .A2(new_n344), .A3(new_n381), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n368), .A2(G150), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n212), .A2(G33), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT69), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n398), .B(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n397), .B1(new_n400), .B2(new_n303), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT71), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n205), .A2(G20), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n397), .B(KEYINPUT71), .C1(new_n400), .C2(new_n303), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n268), .ZN(new_n407));
  INV_X1    g0207(.A(new_n365), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n293), .A2(G50), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n408), .A2(new_n409), .B1(G50), .B2(new_n297), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n282), .A2(new_n283), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n311), .B1(new_n413), .B2(new_n363), .ZN(new_n414));
  MUX2_X1   g0214(.A(G222), .B(G223), .S(G1698), .Z(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n319), .ZN(new_n417));
  INV_X1    g0217(.A(new_n320), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(G226), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G169), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n412), .B(new_n422), .C1(G179), .C2(new_n420), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT76), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT9), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n412), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n410), .B1(new_n406), .B2(new_n268), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT76), .B1(new_n427), .B2(KEYINPUT9), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n420), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n427), .A2(KEYINPUT9), .B1(new_n430), .B2(G190), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n420), .A2(G200), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n432), .A2(KEYINPUT77), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT10), .B1(new_n432), .B2(KEYINPUT77), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT10), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n427), .A2(KEYINPUT9), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n430), .A2(G190), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n438), .A2(new_n439), .A3(new_n432), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n426), .A2(new_n428), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n423), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n396), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT84), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n408), .A2(new_n362), .A3(new_n203), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT12), .B1(new_n297), .B2(G68), .ZN(new_n447));
  OR3_X1    g0247(.A1(new_n297), .A2(KEYINPUT12), .A3(G68), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n368), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n363), .B2(new_n400), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n268), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT11), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(KEYINPUT11), .A3(new_n268), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n449), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT13), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n321), .A2(G1698), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(G226), .B2(G1698), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n347), .A2(new_n348), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G97), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n390), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G238), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n319), .B1(new_n320), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n458), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(G226), .A2(G1698), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n321), .B2(G1698), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n282), .A2(new_n283), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n311), .B1(new_n471), .B2(new_n462), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n472), .A2(KEYINPUT13), .A3(new_n466), .ZN(new_n473));
  OAI21_X1  g0273(.A(G169), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT14), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT78), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n464), .A2(new_n476), .A3(new_n467), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT78), .B1(new_n472), .B2(new_n466), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT13), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n464), .A2(new_n458), .A3(new_n467), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(G179), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT13), .B1(new_n472), .B2(new_n466), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT14), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(G169), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n475), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT79), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n475), .A2(new_n481), .A3(KEYINPUT79), .A4(new_n485), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n457), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n456), .B1(G200), .B2(new_n483), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n479), .A2(G190), .A3(new_n480), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n444), .A2(new_n445), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n445), .B1(new_n444), .B2(new_n495), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n250), .A2(new_n252), .A3(G244), .A4(new_n312), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT4), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n500), .A2(new_n501), .B1(G33), .B2(G283), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n312), .A2(KEYINPUT4), .A3(G244), .ZN(new_n503));
  INV_X1    g0303(.A(G250), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(new_n312), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n282), .A2(new_n283), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n311), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(KEYINPUT5), .A2(G41), .ZN(new_n508));
  NOR2_X1   g0308(.A1(KEYINPUT5), .A2(G41), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(G45), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(G1), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n510), .A2(new_n311), .A3(G274), .A4(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n508), .B2(new_n509), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n311), .ZN(new_n515));
  INV_X1    g0315(.A(G257), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n507), .A2(new_n517), .A3(new_n359), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n507), .A2(new_n517), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n518), .B1(new_n520), .B2(G169), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n297), .A2(G97), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n291), .A2(G33), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n294), .A2(new_n297), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n522), .B1(new_n525), .B2(G97), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n368), .A2(G77), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT6), .ZN(new_n528));
  INV_X1    g0328(.A(G97), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n528), .A2(new_n529), .A3(G107), .ZN(new_n530));
  XNOR2_X1  g0330(.A(G97), .B(G107), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n527), .B1(new_n532), .B2(new_n212), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n285), .B2(G107), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n526), .B1(new_n534), .B2(new_n294), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT85), .ZN(new_n536));
  INV_X1    g0336(.A(new_n533), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n212), .B1(new_n347), .B2(new_n348), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(new_n254), .B1(new_n276), .B2(new_n277), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n539), .B2(new_n353), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n268), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT85), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(new_n526), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n521), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n502), .A2(new_n506), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n390), .ZN(new_n546));
  INV_X1    g0346(.A(new_n517), .ZN(new_n547));
  INV_X1    g0347(.A(G190), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n394), .B1(new_n507), .B2(new_n517), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n541), .A3(new_n526), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n544), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n247), .A2(new_n212), .A3(G87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT22), .ZN(new_n556));
  INV_X1    g0356(.A(G87), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n557), .A2(KEYINPUT22), .A3(G20), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n282), .A2(new_n283), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n212), .A2(G107), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT23), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT23), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n212), .B2(G107), .ZN(new_n564));
  INV_X1    g0364(.A(G116), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n249), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n562), .A2(new_n564), .B1(new_n212), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT24), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n560), .A2(KEYINPUT24), .A3(new_n567), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n268), .A3(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n296), .A2(new_n561), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT89), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT25), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n574), .A2(KEYINPUT25), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI221_X1 g0377(.A(new_n577), .B1(new_n575), .B2(new_n573), .C1(new_n524), .C2(new_n353), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n504), .A2(new_n312), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n516), .A2(G1698), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n250), .A2(new_n581), .A3(new_n252), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G294), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n311), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n514), .A2(G264), .A3(new_n311), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT90), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n514), .A2(KEYINPUT90), .A3(G264), .A4(new_n311), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT91), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n590), .A2(new_n591), .A3(G179), .A4(new_n513), .ZN(new_n592));
  INV_X1    g0392(.A(new_n586), .ZN(new_n593));
  INV_X1    g0393(.A(G274), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n514), .A2(new_n390), .A3(new_n594), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n593), .A2(new_n585), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n592), .B1(new_n421), .B2(new_n596), .ZN(new_n597));
  AOI211_X1 g0397(.A(new_n595), .B(new_n585), .C1(new_n588), .C2(new_n589), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n591), .B1(new_n598), .B2(G179), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n580), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n596), .A2(new_n548), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n598), .B2(G200), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(new_n572), .A3(new_n579), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n373), .A2(new_n297), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT19), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n212), .B1(new_n462), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n557), .A2(new_n529), .A3(new_n353), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT87), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT87), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n247), .A2(new_n212), .A3(G68), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n606), .B1(new_n398), .B2(new_n529), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n611), .A2(new_n612), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n605), .B1(new_n615), .B2(new_n268), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n372), .B2(new_n524), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n311), .A2(G274), .A3(new_n512), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT86), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n311), .A2(KEYINPUT86), .A3(G274), .A4(new_n512), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n512), .A2(new_n504), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n311), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n345), .A2(G1698), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n247), .B(new_n625), .C1(G238), .C2(G1698), .ZN(new_n626));
  INV_X1    g0426(.A(new_n566), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n311), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n421), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n624), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n359), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n617), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n524), .A2(new_n557), .ZN(new_n633));
  AOI211_X1 g0433(.A(new_n605), .B(new_n633), .C1(new_n615), .C2(new_n268), .ZN(new_n634));
  OAI21_X1  g0434(.A(G200), .B1(new_n624), .B2(new_n628), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n626), .A2(new_n627), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n390), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n618), .A2(new_n619), .B1(new_n311), .B2(new_n622), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n637), .A2(G190), .A3(new_n621), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n634), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n632), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n365), .A2(G116), .A3(new_n523), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n304), .A2(new_n565), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n267), .A2(new_n211), .B1(G20), .B2(new_n565), .ZN(new_n644));
  AOI21_X1  g0444(.A(G20), .B1(G33), .B2(G283), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(G33), .B2(new_n529), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n644), .A2(new_n646), .A3(KEYINPUT20), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT20), .B1(new_n644), .B2(new_n646), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n642), .B(new_n643), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(G303), .B1(new_n347), .B2(new_n348), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n516), .A2(new_n312), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n312), .A2(G264), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n247), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n311), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G270), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n513), .B1(new_n515), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n649), .B(G169), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT21), .ZN(new_n658));
  INV_X1    g0458(.A(new_n656), .ZN(new_n659));
  INV_X1    g0459(.A(G303), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n282), .B2(new_n283), .ZN(new_n661));
  INV_X1    g0461(.A(new_n653), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n390), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n659), .A2(new_n663), .A3(G179), .ZN(new_n664));
  INV_X1    g0464(.A(new_n649), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n657), .A2(new_n658), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n657), .A2(new_n658), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n336), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n659), .A2(new_n663), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(G200), .B1(new_n654), .B2(new_n656), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(new_n665), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT88), .A4(new_n665), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n641), .A2(new_n668), .A3(new_n676), .ZN(new_n677));
  AND4_X1   g0477(.A1(new_n499), .A2(new_n554), .A3(new_n604), .A4(new_n677), .ZN(G372));
  NAND3_X1  g0478(.A1(new_n544), .A2(KEYINPUT26), .A3(new_n641), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT92), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n624), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n638), .A2(KEYINPUT92), .A3(new_n621), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n628), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n617), .B(new_n631), .C1(new_n683), .C2(G169), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n634), .B(new_n639), .C1(new_n683), .C2(new_n394), .ZN(new_n685));
  INV_X1    g0485(.A(new_n518), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n421), .B2(new_n519), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n684), .A2(new_n685), .A3(new_n687), .A4(new_n535), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n679), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n600), .A2(new_n668), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n536), .A2(new_n543), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n687), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n603), .A2(new_n552), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n684), .A2(new_n685), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n692), .A2(new_n694), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n691), .A2(new_n697), .A3(new_n684), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n499), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n484), .B1(new_n483), .B2(G169), .ZN(new_n700));
  AOI211_X1 g0500(.A(KEYINPUT14), .B(new_n421), .C1(new_n480), .C2(new_n482), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT79), .B1(new_n702), .B2(new_n481), .ZN(new_n703));
  INV_X1    g0503(.A(new_n489), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n456), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n380), .A2(new_n493), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n343), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n707), .A2(new_n332), .B1(new_n442), .B2(new_n436), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n708), .A2(KEYINPUT93), .A3(new_n423), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT93), .B1(new_n708), .B2(new_n423), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n699), .A2(new_n711), .ZN(G369));
  NAND2_X1  g0512(.A1(new_n296), .A2(new_n212), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G213), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G343), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n580), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n604), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n718), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n600), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n721), .A2(new_n665), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n668), .A2(new_n676), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n668), .B2(new_n726), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n668), .A2(new_n718), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n604), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n600), .B2(new_n718), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n730), .A2(new_n733), .ZN(G399));
  NAND2_X1  g0534(.A1(new_n216), .A2(new_n310), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n291), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n608), .A2(G116), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n737), .A2(new_n738), .B1(new_n210), .B2(new_n736), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT94), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT28), .Z(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  INV_X1    g0542(.A(new_n684), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n688), .B2(KEYINPUT26), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n544), .A2(new_n689), .A3(new_n641), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT97), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT97), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n744), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(new_n697), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n742), .B1(new_n750), .B2(new_n721), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n698), .A2(new_n721), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(KEYINPUT29), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n677), .A2(new_n554), .A3(new_n604), .A4(new_n721), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT96), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(KEYINPUT30), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n519), .A2(new_n590), .A3(new_n630), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n758), .B2(new_n664), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n546), .A2(new_n590), .A3(new_n547), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n654), .A2(new_n656), .A3(new_n359), .ZN(new_n761));
  INV_X1    g0561(.A(new_n757), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n760), .A2(new_n761), .A3(new_n630), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n624), .A2(new_n680), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT92), .B1(new_n638), .B2(new_n621), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n637), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n590), .A2(new_n513), .ZN(new_n767));
  AOI21_X1  g0567(.A(G179), .B1(new_n659), .B2(new_n663), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n766), .A2(new_n520), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n759), .A2(new_n763), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n770), .A2(new_n718), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n770), .A2(new_n718), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n755), .B(new_n773), .C1(KEYINPUT31), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G330), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n754), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n741), .B1(new_n778), .B2(G1), .ZN(G364));
  NAND2_X1  g0579(.A1(new_n212), .A2(G13), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT98), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G45), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n737), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n728), .B2(G330), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n728), .A2(G330), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n728), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n211), .B1(G20), .B2(new_n421), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G179), .A2(G200), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n212), .B1(new_n795), .B2(G190), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n529), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n212), .A2(new_n359), .A3(new_n394), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G190), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n797), .B1(new_n800), .B2(G68), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n212), .A2(new_n359), .A3(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n669), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n799), .A2(new_n336), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n801), .B1(new_n202), .B2(new_n803), .C1(new_n201), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n802), .A2(new_n548), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT101), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(KEYINPUT101), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n806), .B1(G77), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n394), .A2(G179), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(G20), .A3(new_n548), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT102), .Z(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G107), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n795), .A2(G20), .A3(new_n548), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G159), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT32), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n815), .A2(G20), .A3(G190), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n557), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n822), .A2(new_n413), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n814), .A2(new_n818), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n823), .A2(new_n660), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n827), .B(new_n349), .C1(G329), .C2(new_n820), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  INV_X1    g0629(.A(G294), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n807), .A2(new_n829), .B1(new_n830), .B2(new_n796), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT33), .B(G317), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(new_n800), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n817), .A2(G283), .ZN(new_n834));
  INV_X1    g0634(.A(new_n803), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(G322), .B1(new_n804), .B2(G326), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n828), .A2(new_n833), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n794), .B1(new_n826), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n790), .A2(new_n793), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT100), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n349), .A2(G355), .A3(new_n216), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n253), .A2(new_n216), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT99), .Z(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(G45), .B2(new_n209), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n245), .A2(new_n511), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n842), .B1(G116), .B2(new_n216), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n783), .B(new_n838), .C1(new_n841), .C2(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n785), .A2(new_n787), .B1(new_n792), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  NAND2_X1  g0650(.A1(new_n391), .A2(new_n392), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n377), .B1(new_n851), .B2(new_n421), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(new_n360), .A3(new_n721), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n377), .A2(new_n721), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n387), .B1(new_n851), .B2(G200), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n393), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n853), .B1(new_n856), .B2(new_n380), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n752), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n854), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n395), .A2(new_n859), .B1(new_n852), .B2(new_n360), .ZN(new_n860));
  INV_X1    g0660(.A(new_n853), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n698), .A2(new_n721), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n784), .B1(new_n864), .B2(new_n776), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n776), .B2(new_n864), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n835), .A2(G143), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G137), .A2(new_n804), .B1(new_n800), .B2(G150), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n867), .B(new_n868), .C1(new_n812), .C2(new_n257), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT34), .Z(new_n870));
  NOR2_X1   g0670(.A1(new_n823), .A2(new_n201), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n253), .B(new_n871), .C1(G132), .C2(new_n820), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n817), .A2(G68), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n872), .B(new_n873), .C1(new_n202), .C2(new_n796), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n803), .A2(new_n830), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n797), .B(new_n875), .C1(G303), .C2(new_n804), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n823), .A2(new_n353), .B1(new_n819), .B2(new_n829), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n349), .B(new_n877), .C1(new_n817), .C2(G87), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n813), .A2(G116), .B1(G283), .B2(new_n800), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT103), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n876), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n879), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(KEYINPUT103), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n870), .A2(new_n874), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n793), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n793), .A2(new_n788), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n783), .B1(new_n363), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n885), .B(new_n887), .C1(new_n862), .C2(new_n789), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n866), .A2(new_n888), .ZN(G384));
  OAI22_X1  g0689(.A1(new_n496), .A2(new_n497), .B1(new_n751), .B2(new_n753), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n711), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT108), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n287), .B1(new_n256), .B2(new_n271), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n308), .B1(new_n269), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT105), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n308), .B(KEYINPUT105), .C1(new_n269), .C2(new_n893), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(new_n326), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(KEYINPUT106), .A3(new_n339), .ZN(new_n899));
  INV_X1    g0699(.A(new_n716), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT106), .B1(new_n898), .B2(new_n339), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT37), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n309), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n329), .B1(new_n905), .B2(new_n338), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT107), .B1(new_n309), .B2(new_n900), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT107), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n909), .B(new_n716), .C1(new_n288), .C2(new_n308), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n906), .B(new_n907), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n328), .A2(new_n331), .A3(new_n341), .A4(new_n342), .ZN(new_n913));
  INV_X1    g0713(.A(new_n901), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n457), .A2(new_n721), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n705), .A2(new_n493), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n921), .B1(new_n490), .B2(new_n494), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n863), .A2(new_n853), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n920), .A2(new_n925), .B1(new_n332), .B2(new_n716), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n918), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  AOI221_X4 g0728(.A(new_n917), .B1(new_n913), .B2(new_n914), .C1(new_n904), .C2(new_n911), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n908), .A2(new_n910), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n327), .A2(new_n339), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT37), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n911), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n913), .A2(new_n930), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT38), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n928), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n705), .A2(new_n718), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n927), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n892), .B(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n935), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n919), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n770), .A2(KEYINPUT31), .A3(new_n718), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n772), .B1(new_n770), .B2(new_n718), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n857), .B1(new_n755), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n922), .B1(new_n705), .B2(new_n493), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n490), .A2(new_n494), .A3(new_n921), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n943), .A2(new_n951), .A3(KEYINPUT40), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT109), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n950), .B1(new_n919), .B2(new_n918), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n953), .B1(new_n954), .B2(KEYINPUT40), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n923), .A2(new_n924), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT38), .B1(new_n912), .B2(new_n915), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n956), .B(new_n947), .C1(new_n929), .C2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT40), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n958), .A2(KEYINPUT109), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n952), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n755), .A2(new_n946), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n499), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(G330), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n962), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n941), .A2(new_n966), .B1(new_n291), .B2(new_n781), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n941), .B2(new_n966), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n210), .A2(G77), .A3(new_n262), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n291), .B(G13), .C1(new_n969), .C2(new_n241), .ZN(new_n970));
  INV_X1    g0770(.A(new_n532), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT35), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT35), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n972), .A2(G116), .A3(new_n213), .A4(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT104), .B(KEYINPUT36), .Z(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n968), .A2(new_n970), .A3(new_n976), .ZN(G367));
  AND3_X1   g0777(.A1(new_n687), .A2(new_n535), .A3(new_n718), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n535), .A2(new_n718), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(new_n554), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n694), .B1(new_n980), .B2(new_n600), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT110), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(new_n721), .A3(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n980), .A2(new_n732), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT42), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n634), .A2(new_n721), .ZN(new_n988));
  MUX2_X1   g0788(.A(new_n696), .B(new_n743), .S(new_n988), .Z(new_n989));
  AOI22_X1  g0789(.A1(new_n985), .A2(new_n987), .B1(KEYINPUT43), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n990), .B(new_n991), .Z(new_n992));
  INV_X1    g0792(.A(new_n730), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n980), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n992), .B1(KEYINPUT111), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(KEYINPUT111), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n782), .A2(G1), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n733), .A2(new_n980), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT44), .Z(new_n1002));
  NOR2_X1   g0802(.A1(new_n733), .A2(new_n980), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n730), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1002), .A2(new_n993), .A3(new_n1004), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n732), .B1(new_n723), .B2(new_n731), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(new_n729), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n777), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n735), .B(KEYINPUT41), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1000), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n992), .A2(KEYINPUT111), .A3(new_n995), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n998), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n844), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n231), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n841), .B1(new_n216), .B2(new_n372), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n784), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n823), .A2(new_n565), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT46), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n660), .B2(new_n803), .C1(new_n829), .C2(new_n805), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n247), .B1(new_n820), .B2(G317), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n529), .B2(new_n816), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n800), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n1027), .A2(new_n830), .B1(new_n353), .B2(new_n796), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1024), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n813), .A2(G283), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n813), .A2(G50), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G143), .A2(new_n804), .B1(new_n800), .B2(G159), .ZN(new_n1032));
  INV_X1    g0832(.A(G150), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n1033), .B2(new_n803), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n823), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1035), .A2(G58), .B1(new_n820), .B2(G137), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n363), .B2(new_n816), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n349), .B1(new_n203), .B2(new_n796), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1029), .A2(new_n1030), .B1(new_n1031), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT47), .Z(new_n1041));
  AOI21_X1  g0841(.A(new_n1020), .B1(new_n1041), .B2(new_n793), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n791), .B2(new_n989), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1016), .A2(new_n1043), .ZN(G387));
  NOR2_X1   g0844(.A1(new_n777), .A2(new_n1010), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(new_n735), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n778), .B2(new_n1011), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n349), .A2(new_n216), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1048), .A2(new_n738), .B1(G107), .B2(new_n216), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT112), .Z(new_n1050));
  NOR2_X1   g0850(.A1(new_n369), .A2(new_n370), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1051), .A2(G50), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT50), .ZN(new_n1053));
  AOI21_X1  g0853(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n738), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1017), .B1(new_n236), .B2(G45), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1050), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n784), .B1(new_n1057), .B2(new_n840), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT113), .Z(new_n1059));
  AOI22_X1  g0859(.A1(new_n835), .A2(G50), .B1(new_n804), .B2(G159), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n203), .B2(new_n807), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n823), .A2(new_n363), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n253), .B(new_n1062), .C1(G150), .C2(new_n820), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n303), .B2(new_n1027), .C1(new_n372), .C2(new_n796), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1061), .B(new_n1064), .C1(G97), .C2(new_n817), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n804), .A2(G322), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n835), .A2(G317), .B1(new_n800), .B2(G311), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n812), .C2(new_n660), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT48), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n796), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1035), .A2(G294), .B1(new_n1072), .B2(G283), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n247), .B1(new_n820), .B2(G326), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n565), .B2(new_n816), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1065), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1059), .B1(new_n1081), .B2(new_n794), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n724), .B2(new_n790), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1011), .B2(new_n999), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1047), .A2(new_n1084), .ZN(G393));
  AOI21_X1  g0885(.A(new_n735), .B1(new_n1008), .B2(new_n1045), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1006), .A2(KEYINPUT115), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1007), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1086), .B1(new_n1089), .B2(new_n1045), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n844), .A2(new_n240), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1091), .B(new_n841), .C1(new_n529), .C2(new_n216), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n807), .A2(new_n830), .B1(new_n565), .B2(new_n796), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n835), .A2(G311), .B1(new_n804), .B2(G317), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT52), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(G303), .C2(new_n800), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1035), .A2(G283), .B1(new_n820), .B2(G322), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n818), .A2(new_n413), .A3(new_n1097), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT116), .Z(new_n1099));
  OAI22_X1  g0899(.A1(new_n805), .A2(new_n1033), .B1(new_n257), .B2(new_n803), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT51), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n247), .B1(new_n823), .B2(new_n203), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G143), .B2(new_n820), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n363), .B2(new_n796), .C1(new_n201), .C2(new_n1027), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n812), .A2(new_n1051), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G87), .C2(new_n817), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1096), .A2(new_n1099), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n784), .B(new_n1092), .C1(new_n1107), .C2(new_n794), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n980), .B2(new_n790), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n1089), .B2(new_n999), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1090), .A2(new_n1110), .ZN(G390));
  NAND2_X1  g0911(.A1(new_n927), .A2(new_n936), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n788), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT54), .B(G143), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n813), .A2(new_n1115), .B1(G137), .B2(new_n800), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1116), .A2(KEYINPUT120), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(KEYINPUT120), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n823), .A2(KEYINPUT53), .A3(new_n1033), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G128), .B2(new_n804), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n257), .B2(new_n796), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n835), .A2(G132), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n816), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1123), .A2(G50), .B1(new_n820), .B2(G125), .ZN(new_n1124));
  OAI21_X1  g0924(.A(KEYINPUT53), .B1(new_n823), .B2(new_n1033), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1122), .A2(new_n349), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  NOR4_X1   g0926(.A1(new_n1117), .A2(new_n1118), .A3(new_n1121), .A4(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n824), .B(new_n349), .C1(G294), .C2(new_n820), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n796), .A2(new_n363), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n804), .B2(G283), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n835), .A2(G116), .B1(new_n800), .B2(G107), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1128), .A2(new_n873), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n812), .A2(new_n529), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n793), .B1(new_n1127), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n783), .B1(new_n303), .B2(new_n886), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1113), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n937), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n929), .B2(new_n935), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n750), .A2(new_n721), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n853), .B1(new_n1140), .B2(new_n860), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1139), .B1(new_n1141), .B2(new_n956), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT117), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n603), .A2(new_n552), .A3(new_n684), .A4(new_n685), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1144), .A2(new_n544), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n743), .B1(new_n1145), .B2(new_n692), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n718), .B1(new_n1146), .B2(new_n691), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n861), .B1(new_n1147), .B2(new_n862), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n948), .A2(new_n949), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1138), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1143), .A2(new_n1150), .B1(new_n927), .B2(new_n936), .ZN(new_n1151));
  OAI211_X1 g0951(.A(KEYINPUT117), .B(new_n1138), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1142), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n947), .A2(G330), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT118), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT118), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n956), .A2(new_n1156), .A3(G330), .A4(new_n947), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(KEYINPUT119), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n956), .A2(new_n775), .A3(G330), .A4(new_n862), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1153), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1142), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1143), .B1(new_n925), .B2(new_n937), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1112), .A2(new_n1152), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT119), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n1158), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1160), .A2(new_n1162), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1137), .B1(new_n1169), .B2(new_n1000), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1149), .B1(new_n776), .B2(new_n857), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1155), .A2(new_n1171), .A3(new_n1157), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1148), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1174), .A2(new_n1161), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n750), .A2(new_n721), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n860), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n861), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1172), .A2(new_n1173), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(G330), .B(new_n963), .C1(new_n496), .C2(new_n497), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n890), .C1(new_n710), .C2(new_n709), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1160), .A2(new_n1162), .A3(new_n1168), .A4(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1182), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n735), .B1(new_n1169), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1170), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G378));
  NAND3_X1  g0987(.A1(new_n943), .A2(new_n951), .A3(KEYINPUT40), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n954), .A2(new_n953), .A3(KEYINPUT40), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT109), .B1(new_n958), .B2(new_n959), .ZN(new_n1190));
  OAI211_X1 g0990(.A(G330), .B(new_n1188), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n427), .A2(new_n716), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n443), .B(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1193), .B(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1195), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n961), .B2(G330), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n939), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n961), .A2(G330), .A3(new_n1197), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1200), .A2(new_n1201), .A3(new_n940), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1000), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1195), .A2(new_n788), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n886), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n784), .B1(G50), .B2(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n835), .A2(G128), .B1(G137), .B2(new_n808), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G125), .A2(new_n804), .B1(new_n800), .B2(G132), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1035), .A2(new_n1115), .B1(new_n1072), .B2(G150), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1123), .A2(G159), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G33), .B(G41), .C1(new_n820), .C2(G124), .ZN(new_n1214));
  AND4_X1   g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n804), .A2(G116), .B1(new_n808), .B2(new_n373), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n529), .B2(new_n1027), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1062), .B1(G283), .B2(new_n820), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n247), .A2(G41), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n202), .C2(new_n816), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n803), .A2(new_n353), .B1(new_n203), .B2(new_n796), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1217), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT121), .Z(new_n1223));
  AOI21_X1  g1023(.A(new_n1215), .B1(new_n1223), .B2(KEYINPUT58), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1224), .B1(KEYINPUT58), .B2(new_n1223), .C1(new_n1219), .C2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1206), .B1(new_n1226), .B2(new_n793), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1204), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT122), .B1(new_n1203), .B2(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1200), .A2(new_n940), .A3(new_n1201), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n940), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n999), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT122), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1228), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1230), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1181), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1183), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1239), .A3(KEYINPUT57), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1202), .A2(new_n1199), .B1(new_n1183), .B2(new_n1238), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n736), .C1(KEYINPUT57), .C2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT123), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1236), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1243), .B1(new_n1236), .B2(new_n1242), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(G375));
  INV_X1    g1047(.A(new_n1013), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1184), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1149), .A2(new_n788), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n784), .B1(G68), .B2(new_n1205), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n823), .A2(new_n257), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n247), .B1(new_n816), .B2(new_n202), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(G128), .C2(new_n820), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n835), .A2(G137), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n804), .A2(G132), .B1(new_n808), .B2(G150), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n800), .A2(new_n1115), .B1(new_n1072), .B2(G50), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n796), .A2(new_n372), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n565), .A2(new_n1027), .B1(new_n805), .B2(new_n830), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(G283), .C2(new_n835), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n817), .A2(G77), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1035), .A2(G97), .B1(new_n820), .B2(G303), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1262), .A2(new_n413), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n812), .A2(new_n353), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1259), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1252), .B1(new_n1267), .B2(new_n793), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1251), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1179), .B2(new_n1000), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1250), .A2(new_n1271), .ZN(G381));
  NOR2_X1   g1072(.A1(G393), .A2(G396), .ZN(new_n1273));
  INV_X1    g1073(.A(G384), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1090), .A2(new_n1110), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(G378), .A2(G387), .A3(new_n1275), .A4(G381), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1245), .B2(new_n1246), .ZN(G407));
  NAND2_X1  g1077(.A1(new_n1236), .A2(new_n1242), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(KEYINPUT123), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G378), .B1(new_n1279), .B2(new_n1244), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n717), .A2(G213), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(G213), .A3(G407), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT124), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(KEYINPUT124), .A3(G213), .A4(G407), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(G409));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1236), .A2(new_n1242), .A3(G378), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1241), .A2(new_n1248), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1233), .A2(new_n1228), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1186), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1282), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1274), .A2(KEYINPUT125), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1274), .A2(KEYINPUT125), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1179), .A2(new_n1181), .A3(KEYINPUT60), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n736), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT60), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1249), .B2(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1295), .B(new_n1296), .C1(new_n1300), .C2(new_n1270), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1249), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n736), .A3(new_n1297), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1303), .A2(KEYINPUT125), .A3(new_n1274), .A4(new_n1271), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1301), .A2(new_n1304), .A3(KEYINPUT126), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT126), .B1(new_n1301), .B2(new_n1304), .ZN(new_n1306));
  INV_X1    g1106(.A(G2897), .ZN(new_n1307));
  OAI22_X1  g1107(.A1(new_n1305), .A2(new_n1306), .B1(new_n1307), .B2(new_n1281), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1281), .A2(new_n1307), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1301), .A2(new_n1304), .A3(KEYINPUT126), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1308), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1289), .B1(new_n1294), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1294), .A2(new_n1309), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT127), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1016), .B2(new_n1043), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1016), .A2(new_n1321), .A3(new_n1043), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n849), .B1(new_n1047), .B2(new_n1084), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1273), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G390), .A2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1090), .B(new_n1110), .C1(new_n1273), .C2(new_n1325), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1323), .A2(new_n1324), .A3(new_n1327), .A4(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1324), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1330), .B1(new_n1331), .B2(new_n1322), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1294), .A2(KEYINPUT63), .A3(new_n1309), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1317), .A2(new_n1320), .A3(new_n1334), .A4(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1294), .A2(new_n1337), .A3(new_n1309), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1337), .B1(new_n1294), .B2(new_n1309), .ZN(new_n1339));
  NOR3_X1   g1139(.A1(new_n1338), .A2(new_n1316), .A3(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1336), .B1(new_n1340), .B2(new_n1334), .ZN(G405));
  NAND2_X1  g1141(.A1(new_n1278), .A2(G378), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  NOR3_X1   g1143(.A1(new_n1280), .A2(new_n1334), .A3(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1186), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1333), .B1(new_n1345), .B2(new_n1342), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1309), .B1(new_n1344), .B2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1334), .B1(new_n1280), .B2(new_n1343), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1345), .A2(new_n1333), .A3(new_n1342), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1348), .A2(new_n1304), .A3(new_n1301), .A4(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1347), .A2(new_n1350), .ZN(G402));
endmodule


