//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n598, new_n599, new_n600, new_n601, new_n603,
    new_n604, new_n605, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT80), .B(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G155gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT2), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G141gat), .B(G148gat), .Z(new_n210));
  XNOR2_X1  g009(.A(G155gat), .B(G162gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n211), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G197gat), .B(G204gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT22), .ZN(new_n219));
  XNOR2_X1  g018(.A(G211gat), .B(G218gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G211gat), .ZN(new_n223));
  INV_X1    g022(.A(G218gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n220), .B(new_n218), .C1(KEYINPUT22), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT29), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n217), .B1(KEYINPUT3), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT86), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT74), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n226), .B1(new_n222), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT74), .B1(new_n219), .B2(new_n221), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n212), .A2(new_n236), .A3(new_n216), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n235), .B1(new_n238), .B2(KEYINPUT29), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n230), .A2(new_n231), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G228gat), .ZN(new_n241));
  INV_X1    g040(.A(G233gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n236), .B1(new_n235), .B2(KEYINPUT29), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n217), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(new_n239), .A3(new_n243), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G22gat), .ZN(new_n250));
  INV_X1    g049(.A(G22gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n251), .A3(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT85), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n205), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI211_X1 g054(.A(KEYINPUT85), .B(new_n204), .C1(new_n250), .C2(new_n252), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n258));
  NAND2_X1  g057(.A1(G225gat), .A2(G233gat), .ZN(new_n259));
  XOR2_X1   g058(.A(G113gat), .B(G120gat), .Z(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G134gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G127gat), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n264), .B(KEYINPUT70), .Z(new_n265));
  INV_X1    g064(.A(G127gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G134gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT71), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n262), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n260), .A2(new_n261), .A3(new_n267), .A4(new_n264), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n217), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n269), .A2(new_n212), .A3(new_n270), .A4(new_n216), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n259), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n258), .B1(new_n274), .B2(KEYINPUT81), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(new_n237), .A3(new_n271), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n276), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n277), .A2(new_n279), .A3(new_n259), .A4(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n275), .B(new_n281), .C1(KEYINPUT81), .C2(new_n274), .ZN(new_n282));
  INV_X1    g081(.A(new_n258), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G57gat), .B(G85gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT84), .ZN(new_n287));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT6), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n285), .B2(new_n291), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n296), .B2(new_n293), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n298));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT23), .ZN(new_n300));
  AND2_X1   g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT23), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT66), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT23), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n301), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n300), .B1(new_n306), .B2(new_n299), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n311));
  NAND3_X1  g110(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n310), .B2(new_n312), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n307), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n298), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n314), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n320));
  INV_X1    g119(.A(G169gat), .ZN(new_n321));
  INV_X1    g120(.A(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n301), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n319), .A2(new_n320), .A3(new_n300), .A4(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(KEYINPUT67), .A3(new_n316), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n318), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(KEYINPUT68), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n299), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(KEYINPUT23), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n310), .A2(new_n312), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n325), .A2(new_n332), .A3(KEYINPUT25), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT69), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n329), .A2(new_n337), .A3(new_n331), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n323), .B1(new_n301), .B2(KEYINPUT26), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n336), .B1(new_n340), .B2(new_n309), .ZN(new_n341));
  INV_X1    g140(.A(new_n309), .ZN(new_n342));
  AOI211_X1 g141(.A(KEYINPUT69), .B(new_n342), .C1(new_n338), .C2(new_n339), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT27), .B(G183gat), .ZN(new_n344));
  INV_X1    g143(.A(G190gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT28), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n341), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n335), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G226gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(new_n242), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n352), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n348), .B1(new_n328), .B2(new_n334), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(KEYINPUT29), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n235), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G8gat), .B(G36gat), .Z(new_n360));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT75), .B1(new_n355), .B2(new_n354), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n364));
  INV_X1    g163(.A(new_n334), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n318), .B2(new_n327), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n364), .B(new_n352), .C1(new_n366), .C2(new_n348), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n356), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n368), .A2(KEYINPUT76), .A3(new_n235), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT76), .B1(new_n368), .B2(new_n235), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n359), .B(new_n362), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n297), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n359), .B1(new_n369), .B2(new_n370), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT77), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n377), .B(new_n359), .C1(new_n369), .C2(new_n370), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n362), .B(KEYINPUT78), .Z(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n371), .A2(new_n372), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n374), .B1(new_n382), .B2(KEYINPUT79), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n380), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n257), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(G15gat), .B(G43gat), .Z(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT72), .ZN(new_n388));
  XNOR2_X1  g187(.A(G71gat), .B(G99gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n355), .A2(new_n271), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n270), .B(new_n269), .C1(new_n366), .C2(new_n348), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(new_n392), .A3(G227gat), .A4(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT33), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(KEYINPUT32), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n393), .B(KEYINPUT32), .C1(new_n394), .C2(new_n390), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n391), .A2(new_n392), .ZN(new_n400));
  INV_X1    g199(.A(G227gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n401), .B2(new_n242), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(KEYINPUT34), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n403), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT36), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT73), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT36), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n399), .A2(new_n403), .A3(KEYINPUT73), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n409), .A2(new_n404), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT87), .B1(new_n386), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n415));
  INV_X1    g214(.A(new_n413), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n380), .A2(new_n381), .A3(new_n384), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n384), .B1(new_n380), .B2(new_n381), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n417), .A2(new_n418), .A3(new_n374), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n415), .B(new_n416), .C1(new_n419), .C2(new_n257), .ZN(new_n420));
  INV_X1    g219(.A(new_n257), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n380), .A2(new_n381), .A3(new_n373), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n292), .A2(KEYINPUT88), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(G225gat), .A3(G233gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n272), .A2(new_n259), .A3(new_n273), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(KEYINPUT39), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n291), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n427), .B(new_n428), .C1(KEYINPUT39), .C2(new_n425), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT40), .ZN(new_n430));
  OR2_X1    g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n292), .A2(KEYINPUT88), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n430), .ZN(new_n433));
  AND4_X1   g232(.A1(new_n423), .A2(new_n431), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n421), .B1(new_n422), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT38), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n376), .A2(KEYINPUT37), .A3(new_n378), .ZN(new_n437));
  INV_X1    g236(.A(new_n375), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n362), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n436), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n379), .A2(new_n436), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n357), .B2(new_n235), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n368), .A2(new_n358), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n375), .B2(KEYINPUT37), .ZN(new_n446));
  INV_X1    g245(.A(new_n296), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n447), .A3(new_n423), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n446), .A2(new_n448), .A3(new_n294), .A4(new_n371), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n435), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n414), .A2(new_n420), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n382), .A2(KEYINPUT79), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n257), .A2(new_n404), .A3(new_n405), .ZN(new_n453));
  INV_X1    g252(.A(new_n374), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n452), .A2(new_n385), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n404), .A2(new_n411), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT35), .B1(new_n448), .B2(new_n294), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n457), .A2(new_n257), .A3(new_n409), .A4(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n459), .A2(new_n422), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n451), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G57gat), .B(G64gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n463), .B(KEYINPUT92), .Z(new_n464));
  NAND2_X1  g263(.A1(G71gat), .A2(G78gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(G71gat), .A2(G78gat), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT9), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n465), .B(new_n467), .C1(new_n463), .C2(new_n468), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT91), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n471), .A2(new_n472), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT21), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G231gat), .A2(G233gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G127gat), .B(G155gat), .Z(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT20), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT94), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n481), .B(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(G1gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488));
  MUX2_X1   g287(.A(G1gat), .B(new_n487), .S(new_n488), .Z(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(G8gat), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n475), .B2(new_n476), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n485), .B(new_n491), .Z(new_n492));
  XOR2_X1   g291(.A(G183gat), .B(G211gat), .Z(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n485), .B(new_n491), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT98), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G85gat), .ZN(new_n502));
  INV_X1    g301(.A(G92gat), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n501), .A2(KEYINPUT8), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G85gat), .A2(G92gat), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT97), .B1(new_n505), .B2(KEYINPUT7), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT97), .A3(KEYINPUT7), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(KEYINPUT7), .B2(new_n505), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n504), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G99gat), .B(G106gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT99), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OR3_X1    g312(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n514), .A2(new_n515), .B1(G29gat), .B2(G36gat), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n516), .A2(KEYINPUT15), .ZN(new_n517));
  XNOR2_X1  g316(.A(G43gat), .B(G50gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n516), .B2(KEYINPUT15), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n519), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n513), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G232gat), .A2(G233gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT95), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT41), .ZN(new_n528));
  INV_X1    g327(.A(new_n522), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n524), .B(new_n528), .C1(new_n513), .C2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G190gat), .B(G218gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT96), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n527), .A2(KEYINPUT41), .ZN(new_n534));
  XOR2_X1   g333(.A(G134gat), .B(G162gat), .Z(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n533), .A2(new_n536), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n498), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT100), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT10), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n475), .A2(new_n542), .ZN(new_n543));
  OR3_X1    g342(.A1(new_n513), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n513), .B2(new_n543), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n511), .B(new_n475), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n542), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n547), .A2(new_n550), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G120gat), .B(G148gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(G176gat), .B(G204gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n551), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n529), .A2(new_n490), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n523), .B2(new_n490), .ZN(new_n563));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(KEYINPUT89), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT90), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(KEYINPUT18), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(KEYINPUT18), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n522), .B(new_n490), .Z(new_n570));
  XOR2_X1   g369(.A(new_n565), .B(KEYINPUT13), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT11), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n321), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(G197gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT12), .Z(new_n578));
  OR2_X1    g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n540), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n462), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(new_n297), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT101), .B(G1gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(G1324gat));
  INV_X1    g386(.A(new_n422), .ZN(new_n588));
  OAI21_X1  g387(.A(G8gat), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT102), .Z(new_n590));
  XOR2_X1   g389(.A(KEYINPUT16), .B(G8gat), .Z(new_n591));
  NAND4_X1  g390(.A1(new_n462), .A2(new_n422), .A3(new_n583), .A4(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT42), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT103), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n593), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(G1325gat));
  OAI21_X1  g396(.A(G15gat), .B1(new_n584), .B2(new_n416), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n457), .A2(new_n409), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n600), .A2(G15gat), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n598), .B1(new_n584), .B2(new_n601), .ZN(G1326gat));
  NOR2_X1   g401(.A1(new_n584), .A2(new_n257), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT104), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT43), .B(G22gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(G1327gat));
  INV_X1    g405(.A(new_n539), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n498), .A2(new_n582), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n462), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n609), .A2(G29gat), .A3(new_n297), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT45), .Z(new_n611));
  NAND3_X1  g410(.A1(new_n462), .A2(KEYINPUT44), .A3(new_n607), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT44), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n452), .A2(new_n385), .A3(new_n454), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n413), .B1(new_n614), .B2(new_n421), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n615), .A2(new_n450), .B1(new_n456), .B2(new_n460), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n613), .B1(new_n616), .B2(new_n539), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n608), .B(KEYINPUT105), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(G29gat), .B1(new_n620), .B2(new_n297), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n611), .A2(new_n621), .ZN(G1328gat));
  OAI21_X1  g421(.A(G36gat), .B1(new_n620), .B2(new_n588), .ZN(new_n623));
  OR3_X1    g422(.A1(new_n609), .A2(G36gat), .A3(new_n588), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT46), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n625), .A2(KEYINPUT106), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(KEYINPUT106), .ZN(new_n627));
  OAI221_X1 g426(.A(new_n623), .B1(KEYINPUT46), .B2(new_n624), .C1(new_n626), .C2(new_n627), .ZN(G1329gat));
  NAND2_X1  g427(.A1(new_n413), .A2(G43gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n609), .A2(new_n600), .ZN(new_n630));
  OAI22_X1  g429(.A1(new_n620), .A2(new_n629), .B1(G43gat), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g431(.A1(new_n421), .A2(G50gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n609), .A2(new_n257), .ZN(new_n634));
  OAI22_X1  g433(.A1(new_n620), .A2(new_n633), .B1(G50gat), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g435(.A1(new_n616), .A2(new_n540), .A3(new_n581), .A4(new_n561), .ZN(new_n637));
  INV_X1    g436(.A(new_n297), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT107), .B(G57gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1332gat));
  AOI21_X1  g440(.A(new_n588), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(G1333gat));
  INV_X1    g444(.A(new_n637), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n646), .A2(G71gat), .A3(new_n600), .ZN(new_n647));
  OAI21_X1  g446(.A(G71gat), .B1(new_n646), .B2(new_n416), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g449(.A1(new_n637), .A2(new_n421), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT108), .B(G78gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1335gat));
  NOR2_X1   g452(.A1(new_n498), .A2(new_n581), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n561), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n612), .A2(new_n617), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT109), .B1(new_n658), .B2(new_n297), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(G85gat), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n658), .A2(KEYINPUT109), .A3(new_n297), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n615), .A2(new_n450), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n539), .B1(new_n662), .B2(new_n461), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n655), .B1(new_n663), .B2(KEYINPUT110), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT110), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n616), .B2(new_n539), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT51), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n614), .A2(new_n421), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n668), .A2(new_n450), .A3(new_n416), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n459), .A2(new_n422), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(KEYINPUT35), .B2(new_n455), .ZN(new_n671));
  OAI211_X1 g470(.A(KEYINPUT110), .B(new_n607), .C1(new_n669), .C2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n666), .A2(new_n672), .A3(KEYINPUT51), .A4(new_n654), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n664), .A2(KEYINPUT111), .A3(KEYINPUT51), .A4(new_n666), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n667), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n560), .A2(new_n502), .A3(new_n638), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT112), .Z(new_n679));
  OAI22_X1  g478(.A1(new_n660), .A2(new_n661), .B1(new_n677), .B2(new_n679), .ZN(G1336gat));
  NOR2_X1   g479(.A1(new_n588), .A2(G92gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n677), .A2(new_n561), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n503), .B1(new_n657), .B2(new_n422), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT52), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n675), .A2(new_n676), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n560), .B(new_n681), .C1(new_n686), .C2(new_n667), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT52), .ZN(new_n688));
  INV_X1    g487(.A(new_n684), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n685), .A2(new_n690), .ZN(G1337gat));
  OR4_X1    g490(.A1(G99gat), .A2(new_n677), .A3(new_n600), .A4(new_n561), .ZN(new_n692));
  OAI21_X1  g491(.A(G99gat), .B1(new_n658), .B2(new_n416), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(G1338gat));
  INV_X1    g493(.A(KEYINPUT115), .ZN(new_n695));
  OR3_X1    g494(.A1(new_n561), .A2(G106gat), .A3(new_n257), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n677), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n612), .A2(new_n421), .A3(new_n617), .A4(new_n656), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT113), .B(G106gat), .Z(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT114), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT114), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n698), .A2(new_n702), .A3(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT53), .B1(new_n697), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT53), .B1(new_n698), .B2(new_n699), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n695), .A2(KEYINPUT53), .ZN(new_n707));
  OAI22_X1  g506(.A1(new_n677), .A2(new_n696), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(G1339gat));
  NOR2_X1   g508(.A1(new_n540), .A2(new_n581), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n561), .ZN(new_n711));
  INV_X1    g510(.A(new_n498), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n546), .A2(new_n548), .B1(G230gat), .B2(G233gat), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT54), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n558), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n551), .A2(KEYINPUT54), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n549), .A2(new_n550), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT55), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n715), .B(KEYINPUT55), .C1(new_n716), .C2(new_n717), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n720), .A2(new_n581), .A3(new_n559), .A4(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n563), .A2(new_n565), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n570), .A2(new_n571), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n577), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n560), .A2(new_n579), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n607), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n720), .A2(new_n559), .A3(new_n721), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n579), .A2(new_n725), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n728), .A2(new_n539), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n712), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n711), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n600), .A2(new_n421), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n732), .A2(new_n638), .A3(new_n588), .A4(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n581), .ZN(new_n735));
  OAI21_X1  g534(.A(G113gat), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n638), .ZN(new_n737));
  INV_X1    g536(.A(new_n453), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n588), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n735), .A2(G113gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT116), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n736), .B1(new_n740), .B2(new_n742), .ZN(G1340gat));
  INV_X1    g542(.A(G120gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n734), .A2(new_n744), .A3(new_n561), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n739), .A2(new_n588), .A3(new_n560), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n744), .ZN(G1341gat));
  NOR3_X1   g546(.A1(new_n734), .A2(new_n266), .A3(new_n712), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n740), .A2(new_n712), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n749), .A2(KEYINPUT117), .ZN(new_n750));
  AOI21_X1  g549(.A(G127gat), .B1(new_n749), .B2(KEYINPUT117), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(G1342gat));
  OAI21_X1  g551(.A(G134gat), .B1(new_n734), .B2(new_n539), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n539), .A2(G134gat), .A3(new_n422), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n739), .A2(KEYINPUT56), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT56), .B1(new_n739), .B2(new_n754), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT118), .ZN(G1343gat));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n413), .A2(new_n297), .A3(new_n422), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(G141gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n735), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n257), .A2(new_n765), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n722), .A2(KEYINPUT119), .A3(new_n726), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT119), .B1(new_n722), .B2(new_n726), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n539), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n730), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n498), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT120), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n711), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n766), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n732), .A2(new_n421), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n765), .ZN(new_n777));
  AOI211_X1 g576(.A(new_n761), .B(new_n764), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n413), .A2(new_n257), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT121), .Z(new_n780));
  NOR3_X1   g579(.A1(new_n737), .A2(new_n422), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(G141gat), .B1(new_n781), .B2(new_n581), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n759), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n761), .B1(new_n775), .B2(new_n777), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n763), .ZN(new_n785));
  INV_X1    g584(.A(new_n782), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(KEYINPUT58), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(G1344gat));
  INV_X1    g587(.A(G148gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n781), .A2(new_n789), .A3(new_n560), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT59), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G148gat), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n784), .B2(new_n560), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n257), .A2(KEYINPUT57), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n711), .B(KEYINPUT122), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n771), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n776), .A2(KEYINPUT57), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n796), .A2(new_n560), .A3(new_n760), .A4(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n791), .B1(new_n798), .B2(G148gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n790), .B1(new_n793), .B2(new_n799), .ZN(G1345gat));
  NAND3_X1  g599(.A1(new_n781), .A2(new_n208), .A3(new_n498), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n784), .A2(new_n498), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n208), .ZN(G1346gat));
  NAND3_X1  g602(.A1(new_n781), .A2(new_n207), .A3(new_n607), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n784), .A2(new_n607), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n207), .ZN(G1347gat));
  AOI211_X1 g605(.A(new_n638), .B(new_n588), .C1(new_n711), .C2(new_n731), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(new_n453), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n321), .A3(new_n581), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n733), .ZN(new_n810));
  OAI21_X1  g609(.A(G169gat), .B1(new_n810), .B2(new_n735), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(KEYINPUT123), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(KEYINPUT123), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n809), .B1(new_n812), .B2(new_n813), .ZN(G1348gat));
  NAND3_X1  g613(.A1(new_n808), .A2(new_n322), .A3(new_n560), .ZN(new_n815));
  OAI21_X1  g614(.A(G176gat), .B1(new_n810), .B2(new_n561), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1349gat));
  INV_X1    g616(.A(KEYINPUT124), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n498), .A2(new_n344), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n807), .A2(new_n453), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n807), .A2(new_n733), .A3(new_n498), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n818), .A2(new_n820), .B1(new_n821), .B2(G183gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n808), .A2(KEYINPUT124), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n825));
  NAND2_X1  g624(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT125), .A4(KEYINPUT60), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(G1350gat));
  NAND3_X1  g628(.A1(new_n807), .A2(new_n733), .A3(new_n607), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT126), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n830), .A2(new_n831), .A3(G190gat), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n830), .B2(G190gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT61), .ZN(new_n834));
  OR3_X1    g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n834), .B1(new_n832), .B2(new_n833), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n808), .A2(new_n345), .A3(new_n607), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(G1351gat));
  AND2_X1   g637(.A1(new_n796), .A2(new_n797), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n413), .A2(new_n588), .A3(new_n638), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(G197gat), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n841), .A2(new_n842), .A3(new_n735), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n807), .A2(new_n779), .ZN(new_n844));
  AOI21_X1  g643(.A(G197gat), .B1(new_n844), .B2(new_n581), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n845), .ZN(G1352gat));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n561), .A2(G204gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT127), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n839), .A2(new_n560), .A3(new_n840), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(G204gat), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n844), .A2(new_n848), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n850), .B(new_n852), .C1(new_n847), .C2(new_n853), .ZN(G1353gat));
  NAND3_X1  g653(.A1(new_n844), .A2(new_n223), .A3(new_n498), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n796), .A2(new_n498), .A3(new_n797), .A4(new_n840), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n856), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT63), .B1(new_n856), .B2(G211gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(G1354gat));
  OAI21_X1  g658(.A(G218gat), .B1(new_n841), .B2(new_n539), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n224), .A3(new_n607), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1355gat));
endmodule


