//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1228, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g0026(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT65), .B(G20), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n209), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT0), .ZN(new_n235));
  NAND4_X1  g0035(.A1(new_n222), .A2(new_n223), .A3(new_n232), .A4(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(G361));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  INV_X1    g0042(.A(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT2), .B(G226), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT69), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(KEYINPUT82), .ZN(new_n256));
  INV_X1    g0056(.A(G13), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n259), .A2(new_n226), .A3(new_n227), .A4(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(KEYINPUT8), .B(G58), .Z(new_n262));
  NAND2_X1  g0062(.A1(new_n206), .A2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n261), .A2(new_n264), .B1(new_n259), .B2(new_n262), .ZN(new_n265));
  XNOR2_X1  g0065(.A(G58), .B(G68), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n266), .A2(G20), .B1(G159), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n272));
  AOI21_X1  g0072(.A(G20), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT7), .ZN(new_n274));
  OAI21_X1  g0074(.A(G68), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n229), .A2(new_n276), .A3(KEYINPUT7), .ZN(new_n277));
  OAI211_X1 g0077(.A(KEYINPUT16), .B(new_n268), .C1(new_n275), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n226), .A2(new_n227), .A3(new_n260), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT79), .ZN(new_n282));
  INV_X1    g0082(.A(new_n273), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT78), .B1(new_n271), .B2(KEYINPUT3), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT78), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(new_n269), .A3(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n286), .A3(new_n272), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT65), .A2(G20), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT65), .A2(G20), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n288), .A2(new_n289), .A3(new_n274), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n283), .A2(new_n274), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G68), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n268), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT16), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n282), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n287), .A2(new_n290), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n274), .B1(new_n276), .B2(G20), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n268), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n282), .B(new_n294), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n281), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT80), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT79), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n300), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(KEYINPUT80), .A3(new_n281), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n265), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  INV_X1    g0110(.A(G274), .ZN(new_n311));
  INV_X1    g0111(.A(new_n224), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G41), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G41), .ZN(new_n315));
  INV_X1    g0115(.A(G45), .ZN(new_n316));
  AOI21_X1  g0116(.A(G1), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n317), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n312), .A2(new_n313), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n319), .B1(G232), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G1698), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n276), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G223), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n326), .A2(new_n327), .B1(new_n271), .B2(new_n211), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT81), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n276), .A2(G1698), .ZN(new_n330));
  INV_X1    g0130(.A(G226), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n276), .A2(KEYINPUT81), .A3(G226), .A4(G1698), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n328), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n228), .A2(new_n313), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n310), .B(new_n324), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n335), .ZN(new_n337));
  INV_X1    g0137(.A(new_n324), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n336), .B1(new_n339), .B2(G200), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT17), .B1(new_n309), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n265), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT80), .B1(new_n307), .B2(new_n281), .ZN(new_n343));
  AOI211_X1 g0143(.A(new_n303), .B(new_n280), .C1(new_n306), .C2(new_n300), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n340), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT17), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n256), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT18), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n339), .A2(G179), .ZN(new_n351));
  INV_X1    g0151(.A(G169), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n339), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n349), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n350), .B1(new_n349), .B2(new_n353), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n345), .A2(new_n346), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n304), .A2(new_n308), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n358), .A2(KEYINPUT17), .A3(new_n342), .A4(new_n340), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n359), .A3(KEYINPUT82), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n348), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n279), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n288), .A2(new_n289), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n262), .A2(G33), .A3(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n267), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n257), .A2(new_n207), .A3(G1), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n366), .B1(new_n202), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT9), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n279), .A2(new_n367), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(G50), .A3(new_n263), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n368), .B2(new_n371), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n318), .B1(new_n322), .B2(new_n331), .ZN(new_n376));
  XOR2_X1   g0176(.A(KEYINPUT70), .B(G223), .Z(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G1698), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G222), .B2(G1698), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n276), .ZN(new_n380));
  INV_X1    g0180(.A(G77), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n270), .A2(new_n272), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n335), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n376), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G190), .ZN(new_n385));
  INV_X1    g0185(.A(G200), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(new_n384), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT10), .B1(new_n375), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT10), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n385), .B(new_n389), .C1(new_n386), .C2(new_n384), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT72), .B1(new_n373), .B2(new_n374), .ZN(new_n391));
  INV_X1    g0191(.A(new_n374), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(new_n372), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT73), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI211_X1 g0197(.A(KEYINPUT73), .B(new_n390), .C1(new_n391), .C2(new_n394), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n388), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G179), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n384), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n368), .A2(new_n371), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n401), .B(new_n402), .C1(G169), .C2(new_n384), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n367), .A2(new_n292), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT12), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n370), .A2(KEYINPUT71), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT71), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n261), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n409), .A3(new_n263), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n406), .B1(new_n410), .B2(new_n292), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT77), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n412), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n267), .A2(G50), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT76), .B1(new_n207), .B2(G68), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT76), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n363), .A2(G33), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n417), .B1(new_n418), .B2(new_n415), .C1(new_n419), .C2(new_n381), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n279), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT11), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n413), .A2(new_n414), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G97), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G226), .A2(G1698), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n243), .B2(G1698), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n276), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n335), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT74), .ZN(new_n430));
  INV_X1    g0230(.A(G238), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n318), .B1(new_n322), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT75), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n430), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n430), .B2(new_n434), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n424), .B(G169), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n438), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(G179), .A3(new_n436), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n436), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n424), .B1(new_n443), .B2(G169), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n423), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n423), .ZN(new_n446));
  OAI21_X1  g0246(.A(G200), .B1(new_n437), .B2(new_n438), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(G190), .A3(new_n436), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n262), .A2(new_n267), .B1(new_n229), .B2(G77), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT15), .B(G87), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n419), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n279), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n367), .A2(new_n381), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n453), .B(new_n454), .C1(new_n381), .C2(new_n410), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n382), .A2(G107), .ZN(new_n456));
  OAI221_X1 g0256(.A(new_n456), .B1(new_n330), .B2(new_n431), .C1(new_n243), .C2(new_n326), .ZN(new_n457));
  INV_X1    g0257(.A(new_n335), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n319), .B1(G244), .B2(new_n323), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(new_n310), .ZN(new_n462));
  AOI211_X1 g0262(.A(new_n455), .B(new_n462), .C1(G200), .C2(new_n461), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n352), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n459), .A2(new_n400), .A3(new_n460), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n455), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n445), .A2(new_n449), .A3(new_n468), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n361), .A2(new_n404), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT89), .ZN(new_n472));
  INV_X1    g0272(.A(G283), .ZN(new_n473));
  MUX2_X1   g0273(.A(new_n213), .B(new_n473), .S(G33), .Z(new_n474));
  INV_X1    g0274(.A(G116), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n474), .A2(new_n363), .B1(G20), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n476), .A2(KEYINPUT20), .A3(new_n279), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT20), .B1(new_n476), .B2(new_n279), .ZN(new_n478));
  OAI22_X1  g0278(.A1(new_n477), .A2(new_n478), .B1(G116), .B2(new_n259), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n475), .B1(new_n206), .B2(G33), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n407), .A2(new_n409), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT88), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT88), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n407), .A2(new_n409), .A3(new_n483), .A4(new_n480), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n479), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g0285(.A(KEYINPUT5), .B(G41), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n316), .A2(G1), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n486), .A2(new_n487), .B1(new_n312), .B2(new_n313), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n314), .A2(new_n489), .B1(new_n490), .B2(G270), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n382), .A2(G303), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G264), .A2(G1698), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n214), .B2(G1698), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n276), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n495), .A3(KEYINPUT87), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n458), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT87), .B1(new_n492), .B2(new_n495), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n491), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G169), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n472), .B1(new_n485), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n485), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n492), .A2(new_n495), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT87), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n458), .A3(new_n496), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G179), .A3(new_n491), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n501), .A2(KEYINPUT21), .B1(new_n502), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT90), .ZN(new_n510));
  NOR2_X1   g0310(.A1(KEYINPUT23), .A2(G107), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n229), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n271), .B2(new_n475), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n207), .ZN(new_n515));
  INV_X1    g0315(.A(G107), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n512), .B(new_n515), .C1(new_n513), .C2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n363), .A2(new_n276), .A3(G87), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT22), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT22), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n363), .A2(new_n276), .A3(new_n521), .A4(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n510), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n518), .A2(new_n523), .A3(new_n510), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(KEYINPUT24), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT24), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n362), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n367), .A2(new_n516), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT25), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n531), .B(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n370), .B1(G1), .B2(new_n271), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n516), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n276), .A2(G257), .A3(G1698), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT91), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n276), .A2(G250), .A3(new_n325), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n541), .A2(KEYINPUT92), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n541), .A2(KEYINPUT92), .B1(G33), .B2(G294), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n458), .B1(G264), .B2(new_n490), .ZN(new_n545));
  INV_X1    g0345(.A(new_n314), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(new_n488), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(G169), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n542), .A2(new_n543), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n538), .B(KEYINPUT91), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n458), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n490), .A2(G264), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(G179), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n537), .A2(new_n550), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT21), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n472), .B(new_n559), .C1(new_n485), .C2(new_n500), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n509), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT84), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G283), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n276), .A2(G244), .A3(new_n325), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT4), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n563), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n458), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n547), .B1(G257), .B2(new_n490), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n562), .B1(new_n571), .B2(new_n310), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT84), .A4(G190), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(G200), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n296), .A2(new_n297), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G107), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT6), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n213), .A2(new_n516), .ZN(new_n578));
  NOR2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(KEYINPUT6), .A2(G97), .ZN(new_n581));
  OR3_X1    g0381(.A1(new_n581), .A2(KEYINPUT83), .A3(G107), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT83), .B1(new_n581), .B2(G107), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n584), .A2(new_n229), .B1(G77), .B2(new_n267), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n362), .B1(new_n576), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n367), .A2(new_n213), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n534), .B2(new_n213), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n589), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n586), .A2(new_n588), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n569), .A2(new_n570), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n400), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n571), .A2(new_n352), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n535), .B1(new_n527), .B2(new_n529), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n555), .A2(G200), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n545), .A2(G190), .A3(new_n548), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n579), .A2(new_n211), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n425), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n601), .B1(new_n229), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n363), .A2(new_n276), .A3(G68), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n363), .A2(G33), .A3(G97), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n602), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT85), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(KEYINPUT85), .A3(new_n602), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n451), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n612), .A2(new_n362), .B1(new_n259), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT86), .B1(new_n534), .B2(new_n211), .ZN(new_n615));
  INV_X1    g0415(.A(new_n534), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT86), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(G87), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n614), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n321), .B(G250), .C1(G1), .C2(new_n316), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n314), .A2(new_n487), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n276), .A2(G244), .A3(G1698), .ZN(new_n623));
  OAI221_X1 g0423(.A(new_n623), .B1(new_n271), .B2(new_n475), .C1(new_n326), .C2(new_n431), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n622), .B1(new_n624), .B2(new_n458), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G190), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n386), .B2(new_n625), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI211_X1 g0428(.A(G179), .B(new_n622), .C1(new_n624), .C2(new_n458), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n624), .A2(new_n458), .ZN(new_n630));
  INV_X1    g0430(.A(new_n622), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n352), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n616), .A2(new_n613), .ZN(new_n634));
  OAI221_X1 g0434(.A(new_n634), .B1(new_n259), .B2(new_n613), .C1(new_n612), .C2(new_n362), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n619), .A2(new_n628), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n499), .A2(G200), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n485), .B(new_n637), .C1(new_n310), .C2(new_n499), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n596), .A2(new_n600), .A3(new_n636), .A4(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n471), .A2(new_n561), .A3(new_n639), .ZN(G372));
  INV_X1    g0440(.A(KEYINPUT93), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n509), .A2(new_n558), .A3(new_n641), .A4(new_n560), .ZN(new_n642));
  INV_X1    g0442(.A(new_n479), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n482), .A2(new_n484), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n500), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT21), .B1(new_n645), .B2(KEYINPUT89), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n502), .A2(new_n508), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n560), .A3(new_n647), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n597), .A2(new_n549), .A3(new_n556), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT93), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n596), .A2(new_n600), .A3(new_n636), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n642), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n633), .A2(new_n635), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n618), .A2(new_n615), .ZN(new_n655));
  OAI221_X1 g0455(.A(new_n655), .B1(new_n259), .B2(new_n613), .C1(new_n362), .C2(new_n612), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n656), .B2(new_n627), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n653), .B1(new_n657), .B2(new_n595), .ZN(new_n658));
  INV_X1    g0458(.A(new_n595), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n636), .A2(new_n659), .A3(KEYINPUT26), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n658), .A2(new_n660), .B1(new_n635), .B2(new_n633), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n652), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n470), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT94), .ZN(new_n664));
  INV_X1    g0464(.A(new_n403), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n357), .A2(new_n359), .A3(KEYINPUT82), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT82), .B1(new_n357), .B2(new_n359), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n449), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n445), .B1(new_n669), .B2(new_n466), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n356), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n665), .B1(new_n672), .B2(new_n399), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n664), .A2(new_n673), .ZN(G369));
  NAND2_X1  g0474(.A1(new_n363), .A2(new_n258), .ZN(new_n675));
  XOR2_X1   g0475(.A(new_n675), .B(KEYINPUT95), .Z(new_n676));
  INV_X1    g0476(.A(KEYINPUT27), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  AND4_X1   g0479(.A1(G213), .A2(new_n678), .A3(G343), .A4(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n485), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n648), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n638), .ZN(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n537), .A2(new_n680), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n649), .B1(new_n600), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n558), .A2(new_n680), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n680), .B1(new_n509), .B2(new_n560), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n689), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(G399));
  NAND2_X1  g0494(.A1(new_n233), .A2(new_n315), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n206), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n601), .A2(G116), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n697), .A2(new_n698), .B1(new_n231), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n590), .A2(new_n595), .A3(KEYINPUT98), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT98), .B1(new_n590), .B2(new_n595), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n636), .A2(new_n600), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n561), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n680), .B1(new_n706), .B2(new_n661), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n680), .B1(new_n652), .B2(new_n661), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(KEYINPUT29), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n648), .A2(new_n649), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n651), .A2(new_n711), .A3(new_n638), .A4(new_n681), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n507), .A2(new_n632), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n545), .A3(new_n592), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT97), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(KEYINPUT30), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(G179), .B1(new_n506), .B2(new_n491), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n555), .A2(new_n718), .A3(new_n571), .A4(new_n632), .ZN(new_n719));
  INV_X1    g0519(.A(new_n716), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n713), .A2(new_n545), .A3(new_n592), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n717), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n680), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n712), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n710), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n701), .B1(new_n730), .B2(G1), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n229), .A2(new_n257), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G45), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n697), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n686), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(G330), .B1(new_n683), .B2(new_n638), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n684), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n233), .A2(new_n276), .ZN(new_n743));
  INV_X1    g0543(.A(G355), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n743), .A2(new_n744), .B1(G116), .B2(new_n233), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n233), .A2(new_n382), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n316), .B2(new_n231), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n254), .A2(G45), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n228), .B1(new_n207), .B2(G169), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n741), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n735), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G311), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n363), .A2(new_n400), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G190), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n310), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G322), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n755), .A2(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR4_X1   g0562(.A1(new_n207), .A2(new_n310), .A3(new_n386), .A4(G179), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n276), .B1(new_n763), .B2(G303), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT99), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n756), .A2(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G190), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT33), .B(G317), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n766), .A2(new_n310), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G326), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n363), .B1(new_n400), .B2(new_n759), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G179), .A2(G190), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n229), .A2(new_n386), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n773), .A2(G294), .B1(new_n776), .B2(G329), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n765), .A2(new_n769), .A3(new_n771), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n229), .A2(G200), .A3(new_n774), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n762), .B(new_n778), .C1(G283), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT100), .ZN(new_n783));
  INV_X1    g0583(.A(G58), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n784), .A2(new_n760), .B1(new_n758), .B2(new_n381), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(G97), .B2(new_n773), .ZN(new_n786));
  INV_X1    g0586(.A(new_n763), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n276), .B1(new_n779), .B2(new_n516), .C1(new_n787), .C2(new_n211), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G50), .B2(new_n770), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n776), .A2(G159), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n790), .A2(KEYINPUT32), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n767), .A2(G68), .B1(new_n790), .B2(KEYINPUT32), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n786), .A2(new_n789), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n782), .A2(KEYINPUT100), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n783), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n754), .B1(new_n795), .B2(new_n751), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n736), .A2(new_n738), .B1(new_n742), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  AND2_X1   g0598(.A1(new_n680), .A2(new_n455), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n466), .B1(new_n463), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n681), .A2(new_n467), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n709), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n728), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n735), .B1(new_n804), .B2(new_n728), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n751), .A2(new_n739), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n734), .B1(new_n381), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n276), .B1(new_n763), .B2(G107), .ZN(new_n811));
  INV_X1    g0611(.A(new_n770), .ZN(new_n812));
  INV_X1    g0612(.A(G303), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(new_n213), .B2(new_n772), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n758), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G116), .B1(G311), .B2(new_n776), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n211), .B2(new_n779), .C1(new_n817), .C2(new_n760), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n814), .B(new_n818), .C1(G283), .C2(new_n767), .ZN(new_n819));
  INV_X1    g0619(.A(new_n760), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G159), .A2(new_n815), .B1(new_n820), .B2(G143), .ZN(new_n821));
  INV_X1    g0621(.A(new_n767), .ZN(new_n822));
  INV_X1    g0622(.A(G150), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n821), .B1(new_n822), .B2(new_n823), .C1(new_n824), .C2(new_n812), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT34), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n292), .A2(new_n779), .B1(new_n775), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n276), .B1(new_n787), .B2(new_n202), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(G58), .C2(new_n773), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n819), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n810), .B1(new_n750), .B2(new_n831), .C1(new_n803), .C2(new_n740), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n808), .A2(new_n832), .ZN(G384));
  OR2_X1    g0633(.A1(new_n584), .A2(KEYINPUT35), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n584), .A2(KEYINPUT35), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n228), .A2(G116), .A3(new_n229), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT36), .Z(new_n838));
  OAI211_X1 g0638(.A(new_n231), .B(G77), .C1(new_n784), .C2(new_n292), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n202), .A2(G68), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n206), .B(G13), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n678), .A2(new_n679), .A3(G213), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n268), .B1(new_n275), .B2(new_n277), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n846), .A2(new_n294), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n342), .B1(new_n847), .B2(new_n280), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n668), .B2(new_n356), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n353), .A2(new_n848), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(new_n345), .A3(new_n849), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n349), .A2(new_n353), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n349), .A2(new_n845), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n345), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n844), .B1(new_n850), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n339), .A2(new_n352), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G179), .B2(new_n339), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT18), .B1(new_n309), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n349), .A2(new_n350), .A3(new_n353), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n666), .A2(new_n667), .A3(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(KEYINPUT38), .B(new_n858), .C1(new_n866), .C2(new_n849), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(G169), .B1(new_n437), .B2(new_n438), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT14), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n441), .A3(new_n439), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n423), .B(new_n680), .C1(new_n871), .C2(new_n669), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n423), .A2(new_n680), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n445), .A2(new_n449), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n727), .A2(new_n803), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n843), .B1(new_n868), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n854), .A2(new_n855), .A3(new_n345), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n857), .ZN(new_n880));
  INV_X1    g0680(.A(new_n855), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n357), .A2(new_n359), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n881), .B1(new_n865), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n844), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n867), .A2(new_n885), .ZN(new_n886));
  AND4_X1   g0686(.A1(KEYINPUT40), .A2(new_n727), .A3(new_n803), .A4(new_n875), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n877), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n470), .A2(new_n727), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n685), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n470), .B(new_n708), .C1(KEYINPUT29), .C2(new_n709), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n673), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT103), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n886), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n860), .A2(KEYINPUT39), .A3(new_n867), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n871), .A2(new_n423), .A3(new_n681), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n356), .A2(new_n845), .ZN(new_n901));
  INV_X1    g0701(.A(new_n875), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n662), .A2(new_n681), .A3(new_n803), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n801), .B(KEYINPUT102), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n901), .B1(new_n868), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n894), .B(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n891), .A2(KEYINPUT105), .A3(new_n908), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n909), .B1(new_n206), .B2(new_n732), .C1(new_n908), .C2(new_n891), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT105), .B1(new_n891), .B2(new_n908), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n842), .B1(new_n910), .B2(new_n911), .ZN(G367));
  OAI21_X1  g0712(.A(new_n704), .B1(new_n589), .B2(new_n681), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n659), .A2(new_n680), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n915), .A2(new_n690), .A3(new_n692), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT42), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(KEYINPUT106), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT106), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n916), .B2(new_n917), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT43), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n636), .B1(new_n619), .B2(new_n681), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n680), .A2(new_n656), .A3(new_n635), .A4(new_n633), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n916), .A2(new_n917), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n913), .A2(new_n558), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n680), .B1(new_n929), .B2(new_n595), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n922), .A2(new_n923), .A3(new_n927), .A4(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n915), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n691), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n931), .B1(new_n919), .B2(new_n921), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n927), .A2(new_n923), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n932), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n934), .B1(new_n932), .B2(new_n938), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n695), .B(KEYINPUT41), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n690), .B(new_n692), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(new_n686), .Z(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n729), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT109), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT109), .B1(new_n944), .B2(new_n729), .ZN(new_n948));
  INV_X1    g0748(.A(new_n693), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n949), .A2(new_n950), .A3(new_n933), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT45), .B1(new_n693), .B2(new_n915), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n954));
  OR2_X1    g0754(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n949), .A2(new_n933), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(KEYINPUT107), .B(KEYINPUT44), .C1(new_n693), .C2(new_n915), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT108), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n691), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR4_X1   g0762(.A1(new_n953), .A2(new_n958), .A3(new_n960), .A4(new_n691), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n947), .B(new_n948), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n942), .B1(new_n964), .B2(new_n730), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n733), .A2(G1), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n941), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n241), .A2(new_n746), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n752), .B1(new_n233), .B2(new_n451), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n779), .A2(new_n381), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n202), .A2(new_n758), .B1(new_n760), .B2(new_n823), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n970), .B(new_n971), .C1(G137), .C2(new_n776), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n773), .A2(G68), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n973), .B(new_n276), .C1(new_n784), .C2(new_n787), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G143), .B2(new_n770), .ZN(new_n975));
  INV_X1    g0775(.A(G159), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n972), .B(new_n975), .C1(new_n976), .C2(new_n822), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n763), .A2(G116), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT46), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT110), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n776), .A2(G317), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n276), .B1(new_n978), .B2(new_n979), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G294), .A2(new_n767), .B1(new_n770), .B2(G311), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n773), .A2(G107), .B1(new_n780), .B2(G97), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n473), .B2(new_n758), .C1(new_n813), .C2(new_n760), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n977), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT111), .Z(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n735), .B1(new_n968), .B2(new_n969), .C1(new_n990), .C2(new_n750), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n993));
  INV_X1    g0793(.A(new_n741), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n992), .B(new_n993), .C1(new_n994), .C2(new_n926), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n967), .A2(new_n995), .ZN(G387));
  NAND2_X1  g0796(.A1(new_n947), .A2(new_n948), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n695), .B1(new_n944), .B2(new_n729), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n690), .A2(new_n994), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n743), .A2(new_n698), .B1(G107), .B2(new_n233), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n246), .A2(new_n316), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n262), .A2(new_n202), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT50), .Z(new_n1004));
  INV_X1    g0804(.A(new_n698), .ZN(new_n1005));
  AOI211_X1 g0805(.A(G45), .B(new_n1005), .C1(G68), .C2(G77), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n746), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1001), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n735), .B1(new_n1008), .B2(new_n753), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n276), .B1(new_n779), .B2(new_n213), .C1(new_n787), .C2(new_n381), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n262), .B2(new_n767), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G68), .A2(new_n815), .B1(new_n820), .B2(G50), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n772), .A2(new_n451), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G150), .B2(new_n776), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n770), .A2(G159), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n276), .B1(new_n776), .B2(G326), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n755), .A2(new_n822), .B1(new_n812), .B2(new_n761), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT114), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(KEYINPUT114), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G303), .A2(new_n815), .B1(new_n820), .B2(G317), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n773), .A2(G283), .B1(new_n763), .B2(G294), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1017), .B1(new_n475), .B2(new_n779), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1016), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1000), .B(new_n1009), .C1(new_n1031), .C2(new_n751), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n966), .ZN(new_n1033));
  OR3_X1    g0833(.A1(new_n944), .A2(KEYINPUT113), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT113), .B1(new_n944), .B2(new_n1033), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n999), .A2(new_n1036), .ZN(G393));
  OR2_X1    g0837(.A1(new_n959), .A2(new_n691), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n959), .A2(new_n691), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n966), .A3(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n251), .A2(new_n746), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n752), .B1(new_n213), .B2(new_n233), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n735), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n770), .A2(G317), .B1(new_n820), .B2(G311), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n773), .A2(G116), .B1(new_n776), .B2(G322), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n817), .B2(new_n758), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n276), .B1(new_n763), .B2(G283), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n516), .B2(new_n779), .C1(new_n822), .C2(new_n813), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1045), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(KEYINPUT115), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(KEYINPUT115), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n770), .A2(G150), .B1(new_n820), .B2(G159), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT51), .Z(new_n1054));
  NAND2_X1  g0854(.A1(new_n776), .A2(G143), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n772), .A2(new_n381), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n262), .B2(new_n815), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n276), .B1(new_n779), .B2(new_n211), .C1(new_n787), .C2(new_n292), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G50), .B2(new_n767), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1051), .A2(new_n1052), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1043), .B1(new_n1061), .B2(new_n751), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n915), .B2(new_n994), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n964), .A2(new_n696), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n947), .A2(new_n948), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1040), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(G390));
  NAND4_X1  g0866(.A1(new_n727), .A2(new_n875), .A3(G330), .A4(new_n803), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n903), .A2(new_n904), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n899), .B1(new_n1069), .B2(new_n875), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n896), .B2(new_n897), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n707), .A2(new_n800), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n801), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n899), .B1(new_n1073), .B2(new_n875), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n886), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1068), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT39), .B1(new_n867), .B2(new_n885), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n849), .ZN(new_n1079));
  AOI221_X4 g0879(.A(new_n844), .B1(new_n857), .B2(new_n853), .C1(new_n361), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n361), .A2(new_n1079), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT38), .B1(new_n1081), .B2(new_n858), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1078), .B1(new_n1083), .B2(KEYINPUT39), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1067), .B(new_n1075), .C1(new_n1084), .C2(new_n1070), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1077), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n1033), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1084), .A2(new_n740), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n809), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n735), .B1(new_n262), .B2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n213), .A2(new_n758), .B1(new_n760), .B2(new_n475), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1056), .B(new_n1091), .C1(G294), .C2(new_n776), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n382), .B1(new_n779), .B2(new_n292), .C1(new_n787), .C2(new_n211), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G107), .B2(new_n767), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(new_n473), .C2(new_n812), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT54), .B(G143), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n758), .A2(new_n1096), .B1(new_n772), .B2(new_n976), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n382), .B(new_n1097), .C1(G132), .C2(new_n820), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n763), .A2(G150), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT53), .Z(new_n1100));
  AOI22_X1  g0900(.A1(G50), .A2(new_n780), .B1(new_n776), .B2(G125), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G128), .A2(new_n770), .B1(new_n767), .B2(G137), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT117), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1104), .A2(new_n750), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1095), .A2(KEYINPUT117), .A3(new_n1103), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1090), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1087), .B1(new_n1088), .B2(new_n1107), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n561), .A2(new_n639), .A3(new_n680), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n725), .A2(new_n726), .ZN(new_n1110));
  OAI211_X1 g0910(.A(G330), .B(new_n803), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n902), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n801), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n707), .B2(new_n800), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1112), .A2(new_n1067), .A3(new_n1114), .A4(KEYINPUT116), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1067), .A3(new_n1114), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1112), .A2(new_n1067), .B1(new_n903), .B2(new_n904), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1115), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n892), .B(new_n673), .C1(new_n471), .C2(new_n728), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1086), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1077), .A2(new_n1085), .A3(new_n1122), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n696), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1108), .A2(new_n1126), .ZN(G378));
  AND2_X1   g0927(.A1(new_n900), .A2(new_n906), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT38), .B1(new_n880), .B2(new_n883), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n859), .B1(new_n361), .B2(new_n1079), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(KEYINPUT38), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n876), .A2(KEYINPUT40), .ZN(new_n1132));
  OAI21_X1  g0932(.A(G330), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n845), .A2(new_n402), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n404), .B(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n877), .A2(new_n1133), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1136), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1135), .B(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n876), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n843), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n685), .B1(new_n886), .B2(new_n887), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1140), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1128), .B1(new_n1138), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT120), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1137), .B1(new_n877), .B2(new_n1133), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1143), .A2(new_n1144), .A3(new_n1140), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n907), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1146), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1121), .B(KEYINPUT121), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1125), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1128), .B(KEYINPUT120), .C1(new_n1138), .C2(new_n1145), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1146), .A2(KEYINPUT122), .A3(new_n1150), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT122), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1128), .B(new_n1159), .C1(new_n1138), .C2(new_n1145), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1158), .A2(new_n1153), .A3(KEYINPUT57), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n696), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1151), .A2(new_n966), .A3(new_n1154), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n735), .B1(G50), .B2(new_n1089), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT119), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n760), .A2(new_n1167), .B1(new_n787), .B2(new_n1096), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT118), .Z(new_n1169));
  AOI22_X1  g0969(.A1(new_n815), .A2(G137), .B1(new_n773), .B2(G150), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n770), .A2(G125), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n827), .C2(new_n822), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n271), .B(new_n315), .C1(new_n779), .C2(new_n976), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G124), .B2(new_n776), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n776), .A2(G283), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n780), .A2(G58), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n516), .B2(new_n760), .C1(new_n451), .C2(new_n758), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n767), .A2(G97), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n382), .A2(new_n315), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G77), .B2(new_n763), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n973), .A3(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1183), .B(new_n1187), .C1(G116), .C2(new_n770), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1185), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1191));
  AND4_X1   g0991(.A1(new_n1179), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1166), .B1(new_n750), .B2(new_n1192), .C1(new_n1137), .C2(new_n740), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1164), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1163), .A2(new_n1194), .ZN(G375));
  OAI21_X1  g0995(.A(new_n735), .B1(G68), .B2(new_n1089), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1181), .B(new_n276), .C1(new_n976), .C2(new_n787), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1096), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n767), .B2(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n815), .A2(G150), .B1(new_n773), .B2(G50), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n820), .A2(G137), .B1(G128), .B2(new_n776), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n770), .A2(G132), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n760), .A2(new_n473), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1013), .B(new_n1204), .C1(G107), .C2(new_n815), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n276), .B(new_n970), .C1(new_n767), .C2(G116), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(new_n817), .C2(new_n812), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n787), .A2(new_n213), .B1(new_n775), .B2(new_n813), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT123), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1203), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1196), .B1(new_n1210), .B2(new_n751), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n875), .B2(new_n740), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1120), .B2(new_n1033), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT124), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n942), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1123), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1218), .ZN(G381));
  INV_X1    g1019(.A(G375), .ZN(new_n1220));
  INV_X1    g1020(.A(G378), .ZN(new_n1221));
  INV_X1    g1021(.A(G390), .ZN(new_n1222));
  INV_X1    g1022(.A(G384), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1225), .A2(G387), .A3(G381), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1220), .A2(new_n1221), .A3(new_n1226), .ZN(G407));
  INV_X1    g1027(.A(G213), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(G343), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1220), .A2(new_n1221), .A3(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(G407), .A2(new_n1230), .A3(G213), .ZN(G409));
  AOI21_X1  g1031(.A(new_n797), .B1(new_n999), .B2(new_n1036), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1224), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n967), .A2(G390), .A3(new_n995), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G390), .B1(new_n967), .B2(new_n995), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G387), .A2(new_n1222), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G378), .B(new_n1194), .C1(new_n1157), .C2(new_n1162), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1158), .A2(new_n966), .A3(new_n1160), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1193), .B(new_n1243), .C1(new_n1155), .C2(new_n942), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1221), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1229), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT125), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1246), .A2(KEYINPUT125), .A3(new_n1247), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1120), .A2(KEYINPUT60), .A3(new_n1121), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n696), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1123), .A2(KEYINPUT60), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n1254), .B2(new_n1217), .ZN(new_n1255));
  OR3_X1    g1055(.A1(new_n1255), .A2(new_n1214), .A3(new_n1223), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1223), .B1(new_n1255), .B2(new_n1214), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT62), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1250), .A2(KEYINPUT127), .A3(new_n1251), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1229), .A2(G2897), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1258), .B(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT125), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1249), .B(new_n1229), .C1(new_n1242), .C2(new_n1245), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1262), .A2(new_n1263), .A3(new_n1268), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1260), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT127), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1229), .B(new_n1258), .C1(new_n1242), .C2(new_n1245), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(KEYINPUT62), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1241), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1238), .A2(new_n1240), .A3(new_n1263), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1248), .B2(new_n1265), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1248), .B2(new_n1258), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1259), .A2(KEYINPUT63), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1266), .A2(new_n1267), .A3(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT126), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1250), .A2(KEYINPUT63), .A3(new_n1251), .A4(new_n1259), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1284), .A2(new_n1285), .A3(new_n1279), .A4(new_n1277), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1275), .A2(new_n1287), .ZN(G405));
  NOR2_X1   g1088(.A1(new_n1220), .A2(G378), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1242), .ZN(new_n1290));
  OR3_X1    g1090(.A1(new_n1289), .A2(new_n1290), .A3(new_n1259), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1259), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1241), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(new_n1240), .A3(new_n1238), .A4(new_n1292), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(G402));
endmodule


