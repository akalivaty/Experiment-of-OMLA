//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OR3_X1    g0013(.A1(new_n213), .A2(KEYINPUT65), .A3(G13), .ZN(new_n214));
  OAI21_X1  g0014(.A(KEYINPUT65), .B1(new_n213), .B2(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n207), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n202), .C2(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n223), .B(new_n228), .C1(G97), .C2(G257), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n212), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT1), .Z(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n211), .ZN(new_n233));
  AND3_X1   g0033(.A1(new_n203), .A2(new_n205), .A3(G50), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n218), .B(new_n231), .C1(new_n233), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  INV_X1    g0041(.A(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT66), .B(G250), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n240), .B(new_n245), .Z(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND2_X1  g0053(.A1(G58), .A2(G68), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n203), .A2(new_n205), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT76), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G159), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT76), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n255), .A2(new_n260), .A3(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT77), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n257), .A2(KEYINPUT77), .A3(new_n259), .A4(new_n261), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n266), .A2(new_n267), .A3(G20), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT78), .B1(new_n268), .B2(KEYINPUT7), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(KEYINPUT7), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n211), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT78), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT7), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n269), .A2(new_n270), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G68), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n264), .A2(new_n265), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT16), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n232), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT75), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n275), .A2(new_n277), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n270), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n275), .A2(KEYINPUT75), .A3(new_n277), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G68), .A3(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n264), .A2(KEYINPUT16), .A3(new_n265), .A4(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n283), .A2(new_n285), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n285), .B1(new_n210), .B2(G20), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n299), .B2(new_n294), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n273), .A2(new_n274), .ZN(new_n302));
  INV_X1    g0102(.A(G1698), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(G226), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G223), .A2(G1698), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n304), .A2(new_n305), .B1(new_n272), .B2(new_n221), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G41), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(G1), .A3(G13), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n210), .B(G274), .C1(G41), .C2(G45), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(G232), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G200), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT80), .B(G190), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n310), .A2(new_n316), .A3(new_n311), .A4(new_n313), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n292), .A2(new_n301), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT17), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT18), .ZN(new_n320));
  AND4_X1   g0120(.A1(G179), .A2(new_n310), .A3(new_n311), .A4(new_n313), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(G169), .B2(new_n314), .ZN(new_n322));
  AOI211_X1 g0122(.A(new_n320), .B(new_n322), .C1(new_n292), .C2(new_n301), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n281), .A2(new_n282), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n291), .A2(new_n285), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n301), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n322), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT18), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT79), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n325), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n300), .B1(new_n330), .B2(new_n283), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n320), .B1(new_n331), .B2(new_n322), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT79), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n326), .A2(KEYINPUT18), .A3(new_n327), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n319), .A2(new_n329), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n311), .B(KEYINPUT73), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n308), .A2(new_n312), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n266), .A2(new_n267), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n237), .B2(G1698), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n226), .A2(new_n303), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n340), .A2(new_n341), .B1(G33), .B2(G97), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n337), .B1(new_n227), .B2(new_n338), .C1(new_n342), .C2(new_n308), .ZN(new_n343));
  XOR2_X1   g0143(.A(new_n343), .B(KEYINPUT13), .Z(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT14), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(G179), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n343), .B(KEYINPUT13), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(G169), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n258), .A2(G50), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(KEYINPUT74), .B1(G20), .B2(new_n202), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n211), .A2(G33), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n353), .B1(KEYINPUT74), .B2(new_n352), .C1(new_n207), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n202), .B2(new_n299), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n210), .A2(new_n202), .A3(G13), .A4(G20), .ZN(new_n358));
  XOR2_X1   g0158(.A(new_n358), .B(KEYINPUT12), .Z(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT11), .B1(new_n355), .B2(new_n285), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n351), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n344), .A2(G190), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n348), .A2(G200), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n336), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n303), .A2(G222), .ZN(new_n369));
  AND2_X1   g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n302), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n207), .B2(new_n302), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT68), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n309), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n311), .B1(new_n338), .B2(new_n226), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT67), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(G50), .B1(new_n211), .B2(G1), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT69), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n284), .A2(new_n232), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT69), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(G50), .C1(new_n211), .C2(G1), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n381), .A2(new_n382), .A3(new_n295), .A4(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(G50), .B2(new_n295), .ZN(new_n386));
  XOR2_X1   g0186(.A(new_n386), .B(KEYINPUT70), .Z(new_n387));
  NAND2_X1  g0187(.A1(new_n258), .A2(G150), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n388), .B1(new_n354), .B2(new_n293), .C1(new_n206), .C2(new_n211), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n387), .B1(new_n382), .B2(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n391), .A2(KEYINPUT9), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(KEYINPUT9), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n379), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT10), .B1(new_n394), .B2(KEYINPUT72), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n377), .A2(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n394), .B(new_n396), .C1(KEYINPUT72), .C2(KEYINPUT10), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n377), .A2(new_n345), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n400), .B(new_n391), .C1(G179), .C2(new_n377), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G20), .A2(G77), .ZN(new_n403));
  INV_X1    g0203(.A(new_n258), .ZN(new_n404));
  OR2_X1    g0204(.A1(KEYINPUT15), .A2(G87), .ZN(new_n405));
  NAND2_X1  g0205(.A1(KEYINPUT15), .A2(G87), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n403), .B1(new_n293), .B2(new_n404), .C1(new_n407), .C2(new_n354), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n285), .B1(new_n207), .B2(new_n296), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n207), .B2(new_n299), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT71), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G238), .A2(G1698), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n302), .B(new_n413), .C1(new_n237), .C2(G1698), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n309), .C1(G107), .C2(new_n302), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(new_n311), .C1(new_n220), .C2(new_n338), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n378), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(G200), .B2(new_n416), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n345), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n416), .A2(G179), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n411), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n368), .A2(new_n402), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT6), .ZN(new_n426));
  INV_X1    g0226(.A(G97), .ZN(new_n427));
  INV_X1    g0227(.A(G107), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(G97), .A2(G107), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(KEYINPUT6), .A3(G97), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n211), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n279), .B2(G107), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n404), .A2(new_n207), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n285), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n210), .A2(G33), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n295), .A2(new_n439), .A3(new_n232), .A4(new_n284), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(G97), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n296), .A2(new_n427), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G45), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G1), .ZN(new_n448));
  NOR2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  AND2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n448), .B(G274), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n448), .B1(new_n450), .B2(new_n449), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n308), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n453), .B2(new_n242), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT85), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT84), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT84), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G33), .A3(G283), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(G250), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n461));
  OAI211_X1 g0261(.A(G244), .B(new_n303), .C1(new_n266), .C2(new_n267), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT83), .A2(KEYINPUT4), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n460), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n309), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT85), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n451), .C1(new_n453), .C2(new_n242), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n455), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G169), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n455), .A2(new_n467), .A3(G179), .A4(new_n469), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n438), .A2(new_n446), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT82), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n382), .B1(new_n434), .B2(new_n436), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(new_n445), .ZN(new_n476));
  AOI211_X1 g0276(.A(new_n435), .B(new_n433), .C1(new_n279), .C2(G107), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n446), .B(KEYINPUT82), .C1(new_n477), .C2(new_n382), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G200), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(G190), .B2(new_n470), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n473), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n211), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT22), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT22), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n302), .A2(new_n486), .A3(new_n211), .A4(G87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n272), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n211), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n211), .A2(G107), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT23), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n488), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(KEYINPUT24), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT24), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n485), .A2(new_n487), .B1(new_n211), .B2(new_n490), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(new_n493), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n285), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n441), .A2(new_n442), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G107), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT89), .B1(new_n295), .B2(G107), .ZN(new_n502));
  XOR2_X1   g0302(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n295), .A2(KEYINPUT89), .A3(G107), .ZN(new_n505));
  XOR2_X1   g0305(.A(new_n504), .B(new_n505), .Z(new_n506));
  NAND2_X1  g0306(.A1(new_n242), .A2(G1698), .ZN(new_n507));
  OAI221_X1 g0307(.A(new_n507), .B1(G250), .B2(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G294), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n308), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n452), .A2(G264), .A3(new_n308), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n511), .A2(new_n513), .A3(new_n378), .A4(new_n451), .ZN(new_n514));
  INV_X1    g0314(.A(new_n451), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n510), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(G200), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n499), .A2(new_n501), .A3(new_n506), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT90), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n494), .A2(KEYINPUT24), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n497), .A2(new_n496), .A3(new_n493), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(new_n285), .B1(new_n500), .B2(G107), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT90), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(new_n506), .A4(new_n517), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n506), .ZN(new_n527));
  INV_X1    g0327(.A(G179), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n516), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n516), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n345), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n452), .A2(G270), .A3(new_n308), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G303), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n308), .B1(new_n339), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n303), .A2(G257), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G264), .A2(G1698), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n538), .C1(new_n266), .C2(new_n267), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT87), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n273), .A2(new_n535), .A3(new_n274), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n539), .A2(new_n309), .A3(new_n541), .A4(KEYINPUT87), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n451), .B(new_n534), .C1(new_n540), .C2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n295), .A2(G116), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n440), .A2(new_n489), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n211), .B1(new_n427), .B2(G33), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n457), .B2(new_n459), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT20), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n489), .A2(G20), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n285), .A2(new_n552), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n549), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n460), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n284), .A2(new_n232), .B1(G20), .B2(new_n489), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT20), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n546), .B(new_n548), .C1(new_n554), .C2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n544), .A2(new_n559), .A3(G169), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n539), .A2(new_n309), .A3(new_n541), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n542), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n566), .A2(new_n451), .A3(new_n534), .A4(new_n316), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n551), .B1(new_n550), .B2(new_n553), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n556), .A2(KEYINPUT20), .A3(new_n557), .ZN(new_n569));
  AOI211_X1 g0369(.A(new_n545), .B(new_n547), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  AOI211_X1 g0370(.A(new_n515), .B(new_n533), .C1(new_n565), .C2(new_n542), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n567), .B(new_n570), .C1(new_n571), .C2(new_n480), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(G179), .A3(new_n559), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n544), .A2(new_n559), .A3(KEYINPUT21), .A4(G169), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n562), .A2(new_n572), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n221), .A2(new_n427), .A3(new_n428), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G97), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n211), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n578), .A3(KEYINPUT19), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n211), .B(G68), .C1(new_n266), .C2(new_n267), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n354), .B2(new_n427), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n285), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n295), .B1(new_n405), .B2(new_n406), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT86), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n584), .A2(KEYINPUT86), .A3(new_n586), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n448), .A2(G274), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n308), .B(G250), .C1(G1), .C2(new_n447), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n273), .A2(new_n274), .B1(new_n220), .B2(G1698), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n227), .A2(new_n303), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n490), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n592), .B(new_n593), .C1(new_n596), .C2(new_n308), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G190), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n500), .A2(G87), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(G200), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n591), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n407), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n441), .A2(new_n442), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT86), .B1(new_n584), .B2(new_n586), .ZN(new_n605));
  AOI211_X1 g0405(.A(new_n588), .B(new_n585), .C1(new_n583), .C2(new_n285), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n598), .A2(new_n528), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n597), .A2(new_n345), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n575), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n483), .A2(new_n526), .A3(new_n532), .A4(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n425), .A2(new_n613), .ZN(G372));
  INV_X1    g0414(.A(new_n366), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n363), .B1(new_n422), .B2(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n616), .A2(new_n319), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n332), .A2(new_n334), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n399), .B(new_n398), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n620), .A2(new_n401), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n562), .A2(new_n573), .A3(new_n574), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n532), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT91), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(new_n609), .B1(new_n598), .B2(new_n528), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n625), .B(new_n607), .C1(new_n624), .C2(new_n609), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(new_n602), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n623), .A2(new_n526), .A3(new_n483), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n471), .A2(new_n472), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n476), .A2(new_n629), .A3(new_n478), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT26), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n473), .A2(new_n602), .A3(new_n610), .ZN(new_n633));
  XOR2_X1   g0433(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n628), .B(new_n626), .C1(new_n632), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n424), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n621), .A2(new_n637), .ZN(G369));
  NAND3_X1  g0438(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT93), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n642));
  INV_X1    g0442(.A(G213), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n640), .B2(KEYINPUT93), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n523), .B2(new_n506), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT95), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT95), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n650), .A2(new_n526), .A3(new_n532), .A4(new_n651), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT96), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT96), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n532), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n623), .B(new_n648), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n653), .B(new_n654), .C1(new_n532), .C2(new_n648), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n622), .A2(new_n570), .A3(new_n648), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n575), .B1(new_n559), .B2(new_n647), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(KEYINPUT94), .B(G330), .Z(new_n662));
  AND2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n657), .A2(new_n664), .ZN(G399));
  INV_X1    g0465(.A(new_n216), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n576), .A2(G116), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n667), .A2(new_n210), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n234), .B2(new_n667), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT28), .Z(new_n671));
  NAND2_X1  g0471(.A1(new_n636), .A2(new_n648), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT29), .ZN(new_n673));
  INV_X1    g0473(.A(new_n470), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n597), .A2(new_n510), .A3(new_n512), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(G179), .A4(new_n571), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT30), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n571), .A2(G179), .A3(new_n598), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n679), .A2(new_n530), .A3(new_n470), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n647), .ZN(new_n683));
  OAI211_X1 g0483(.A(KEYINPUT31), .B(new_n683), .C1(new_n613), .C2(new_n647), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n683), .A2(KEYINPUT31), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n684), .A2(new_n662), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n627), .A2(new_n631), .A3(KEYINPUT26), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n633), .A2(new_n634), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n628), .A3(new_n626), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n648), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT29), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n673), .A2(new_n687), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n671), .B1(new_n695), .B2(G1), .ZN(G364));
  INV_X1    g0496(.A(G13), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G20), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n210), .B1(new_n698), .B2(G45), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n667), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n663), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n662), .B2(new_n661), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n234), .A2(new_n447), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n339), .B(new_n704), .C1(new_n249), .C2(new_n447), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n302), .A2(G355), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n216), .A3(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(G1), .B(G13), .C1(new_n211), .C2(G169), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT97), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(KEYINPUT97), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n707), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(G116), .B2(new_n666), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n528), .A2(new_n480), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n211), .A2(G190), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G317), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT33), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n722), .A2(KEYINPUT33), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G283), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n480), .A2(G179), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(G20), .A3(new_n378), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G20), .A3(G190), .ZN(new_n729));
  OAI221_X1 g0529(.A(new_n725), .B1(new_n726), .B2(new_n728), .C1(new_n535), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G179), .A2(G200), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n211), .B1(new_n731), .B2(G190), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n302), .B(new_n730), .C1(G294), .C2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n316), .A2(G20), .A3(new_n718), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT98), .B(G326), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n528), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n719), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G311), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n719), .A2(new_n731), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT99), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n316), .A2(G20), .A3(new_n739), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n745), .A2(G329), .B1(G322), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n734), .A2(new_n738), .A3(new_n742), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n728), .A2(new_n428), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n729), .A2(new_n221), .B1(new_n740), .B2(new_n207), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n750), .B(new_n751), .C1(G68), .C2(new_n721), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n732), .A2(new_n427), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n339), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G50), .A2(new_n736), .B1(new_n747), .B2(G58), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G159), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n743), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT32), .Z(new_n759));
  OAI21_X1  g0559(.A(new_n749), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n717), .B1(new_n760), .B2(new_n711), .ZN(new_n761));
  INV_X1    g0561(.A(new_n714), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n701), .B(new_n761), .C1(new_n661), .C2(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n703), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(G396));
  INV_X1    g0565(.A(KEYINPUT102), .ZN(new_n766));
  OR3_X1    g0566(.A1(new_n422), .A2(new_n766), .A3(new_n648), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n419), .B(new_n422), .C1(new_n412), .C2(new_n648), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n766), .B1(new_n422), .B2(new_n648), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n672), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n636), .A2(new_n648), .A3(new_n770), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n687), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT103), .ZN(new_n776));
  INV_X1    g0576(.A(new_n701), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n774), .A2(new_n687), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(KEYINPUT103), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n711), .A2(new_n712), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n207), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n720), .A2(new_n726), .B1(new_n740), .B2(new_n489), .ZN(new_n783));
  INV_X1    g0583(.A(new_n729), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n753), .B(new_n783), .C1(G107), .C2(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n745), .A2(G311), .B1(G294), .B2(new_n747), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n736), .A2(G303), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n728), .A2(new_n221), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n302), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n785), .A2(new_n786), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n728), .A2(new_n202), .B1(new_n732), .B2(new_n201), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n339), .B1(new_n745), .B2(G132), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT101), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n794), .B1(new_n793), .B2(new_n792), .C1(new_n225), .C2(new_n729), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n747), .A2(G143), .B1(G150), .B2(new_n721), .ZN(new_n796));
  INV_X1    g0596(.A(G137), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n796), .B1(new_n797), .B2(new_n735), .C1(new_n757), .C2(new_n740), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n790), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n777), .B1(new_n801), .B2(new_n711), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n782), .B(new_n802), .C1(new_n770), .C2(new_n713), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n780), .A2(new_n803), .ZN(G384));
  NAND3_X1  g0604(.A1(new_n234), .A2(G77), .A3(new_n254), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT104), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G50), .B2(new_n202), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(G1), .A3(new_n697), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n431), .A2(new_n432), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n489), .B1(new_n809), .B2(KEYINPUT35), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n810), .B(new_n233), .C1(KEYINPUT35), .C2(new_n809), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT36), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT40), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n645), .B(KEYINPUT106), .Z(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n326), .B1(new_n327), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n816), .A2(new_n318), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n264), .A2(new_n265), .A3(new_n290), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n818), .A2(new_n282), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n301), .B1(new_n819), .B2(new_n325), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n327), .ZN(new_n821));
  INV_X1    g0621(.A(new_n645), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n821), .A2(new_n823), .A3(new_n318), .ZN(new_n824));
  MUX2_X1   g0624(.A(new_n817), .B(new_n824), .S(KEYINPUT37), .Z(new_n825));
  INV_X1    g0625(.A(new_n823), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n336), .A2(KEYINPUT105), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT105), .B1(new_n336), .B2(new_n826), .ZN(new_n828));
  OAI211_X1 g0628(.A(KEYINPUT38), .B(new_n825), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT38), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n331), .B(new_n814), .C1(new_n319), .C2(new_n618), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n817), .B(KEYINPUT37), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT108), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n684), .A2(new_n835), .A3(new_n685), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n684), .B2(new_n685), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n363), .B(new_n366), .C1(new_n361), .C2(new_n648), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n362), .B(new_n647), .C1(new_n615), .C2(new_n351), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n771), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n813), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n838), .A2(new_n813), .A3(new_n841), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n830), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n844), .B1(new_n846), .B2(new_n829), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n424), .A2(new_n838), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n662), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n846), .A2(KEYINPUT39), .A3(new_n829), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT39), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n834), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n363), .A2(new_n647), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n619), .A2(new_n814), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n846), .A2(new_n829), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n839), .A2(new_n840), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n422), .A2(new_n647), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n773), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n856), .A2(new_n857), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT107), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n673), .A2(new_n693), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(new_n866), .B2(new_n424), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n865), .A3(new_n424), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n621), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n864), .B(new_n871), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n851), .A2(new_n872), .B1(new_n210), .B2(new_n698), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT109), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n851), .A2(new_n872), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n808), .B(new_n812), .C1(new_n874), .C2(new_n875), .ZN(G367));
  AOI22_X1  g0676(.A1(G143), .A2(new_n736), .B1(new_n747), .B2(G150), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n202), .B2(new_n732), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G58), .A2(new_n784), .B1(new_n721), .B2(G159), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n879), .B1(new_n225), .B2(new_n740), .C1(new_n797), .C2(new_n743), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n728), .A2(new_n207), .ZN(new_n881));
  NOR4_X1   g0681(.A1(new_n878), .A2(new_n880), .A3(new_n339), .A4(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT115), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n784), .A2(KEYINPUT46), .A3(G116), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT46), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n729), .B2(new_n489), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n884), .B(new_n886), .C1(new_n428), .C2(new_n732), .ZN(new_n887));
  INV_X1    g0687(.A(new_n728), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n302), .B(new_n887), .C1(G97), .C2(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(G294), .A2(new_n721), .B1(new_n741), .B2(G283), .ZN(new_n890));
  INV_X1    g0690(.A(G311), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n735), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(G303), .B2(new_n747), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n889), .B(new_n893), .C1(new_n722), .C2(new_n743), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n883), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT47), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n777), .B1(new_n896), .B2(new_n711), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n216), .A2(new_n339), .ZN(new_n898));
  OAI221_X1 g0698(.A(new_n715), .B1(new_n216), .B2(new_n407), .C1(new_n245), .C2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT114), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n648), .B1(new_n591), .B2(new_n600), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n626), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n627), .B2(new_n901), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT110), .Z(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n897), .B(new_n900), .C1(new_n905), .C2(new_n762), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n622), .A2(new_n647), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n655), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n483), .B1(new_n479), .B2(new_n648), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n631), .A2(new_n647), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n914), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n912), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n912), .A2(new_n656), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n648), .B1(new_n921), .B2(new_n473), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n918), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT112), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n658), .A2(new_n663), .A3(new_n912), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n919), .B1(new_n918), .B2(new_n922), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT43), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n929), .B2(new_n904), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n925), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n927), .B1(new_n925), .B2(new_n930), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n667), .B(KEYINPUT41), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n657), .A2(new_n483), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT44), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n657), .A2(new_n912), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT45), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n938), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n664), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n937), .A2(new_n664), .A3(new_n940), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT113), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n908), .B1(new_n663), .B2(new_n944), .C1(new_n658), .C2(new_n907), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n663), .A2(new_n944), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n942), .A2(new_n695), .A3(new_n943), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n935), .B1(new_n951), .B2(new_n695), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n700), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n906), .B1(new_n933), .B2(new_n953), .ZN(G387));
  OAI21_X1  g0754(.A(new_n339), .B1(new_n728), .B2(new_n489), .ZN(new_n955));
  INV_X1    g0755(.A(G322), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n735), .A2(new_n956), .B1(new_n891), .B2(new_n720), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT116), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n535), .B2(new_n740), .C1(new_n722), .C2(new_n746), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT48), .ZN(new_n960));
  INV_X1    g0760(.A(G294), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n960), .B1(new_n726), .B2(new_n732), .C1(new_n961), .C2(new_n729), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT49), .Z(new_n963));
  INV_X1    g0763(.A(new_n743), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n955), .B(new_n963), .C1(new_n737), .C2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G50), .A2(new_n747), .B1(new_n736), .B2(G159), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n427), .B2(new_n728), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G68), .A2(new_n741), .B1(new_n964), .B2(G150), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n207), .B2(new_n729), .C1(new_n293), .C2(new_n720), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n732), .A2(new_n407), .ZN(new_n970));
  NOR4_X1   g0770(.A1(new_n967), .A2(new_n969), .A3(new_n339), .A4(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n711), .B1(new_n965), .B2(new_n971), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n240), .A2(G45), .A3(new_n339), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n293), .A2(KEYINPUT50), .A3(G50), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT50), .B1(new_n293), .B2(G50), .ZN(new_n975));
  NAND2_X1  g0775(.A1(G68), .A2(G77), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n974), .A2(new_n975), .A3(new_n447), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n668), .B1(new_n977), .B2(new_n339), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n216), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n979), .B(new_n715), .C1(new_n428), .C2(new_n216), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n972), .A2(new_n701), .A3(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT117), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n658), .B2(new_n762), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n950), .A2(new_n700), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n950), .A2(new_n695), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n948), .A2(new_n694), .A3(new_n949), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n667), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n983), .A2(new_n984), .A3(new_n987), .ZN(G393));
  OAI221_X1 g0788(.A(new_n715), .B1(new_n427), .B2(new_n216), .C1(new_n898), .C2(new_n252), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n720), .A2(new_n535), .B1(new_n732), .B2(new_n489), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n990), .A2(KEYINPUT119), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(KEYINPUT119), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n339), .B1(new_n728), .B2(new_n428), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n729), .A2(new_n726), .B1(new_n740), .B2(new_n961), .ZN(new_n994));
  NOR4_X1   g0794(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n891), .A2(new_n746), .B1(new_n735), .B2(new_n722), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT52), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n995), .B(new_n997), .C1(new_n956), .C2(new_n743), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G50), .A2(new_n721), .B1(new_n741), .B2(new_n294), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n964), .A2(G143), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n202), .C2(new_n729), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G77), .B2(new_n733), .ZN(new_n1002));
  INV_X1    g0802(.A(G150), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n1003), .A2(new_n735), .B1(new_n746), .B2(new_n757), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT51), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n302), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n998), .B1(new_n1006), .B2(new_n788), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n777), .B1(new_n1007), .B2(new_n711), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n989), .B(new_n1008), .C1(new_n912), .C2(new_n762), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT118), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n942), .B2(new_n943), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n943), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1013), .A2(KEYINPUT118), .A3(new_n941), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1010), .B1(new_n1015), .B2(new_n700), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n985), .B1(new_n1013), .B2(new_n941), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n951), .A2(new_n1017), .A3(new_n667), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(G390));
  NAND2_X1  g0819(.A1(new_n849), .A2(G330), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n869), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n621), .C1(new_n1021), .C2(new_n867), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n770), .A2(G330), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n859), .B1(new_n838), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n686), .A2(new_n770), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n859), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n861), .B1(new_n692), .B2(new_n771), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1025), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT120), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n838), .A2(new_n1032), .A3(new_n859), .A4(new_n1024), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n684), .A2(new_n685), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT108), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n684), .A2(new_n685), .A3(new_n835), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1035), .A2(new_n859), .A3(new_n1036), .A4(new_n1024), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT120), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1033), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1040), .A2(KEYINPUT121), .A3(new_n862), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(KEYINPUT121), .B1(new_n1040), .B2(new_n862), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1031), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n852), .A2(new_n854), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n855), .B1(new_n862), .B2(new_n859), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n855), .B1(new_n1029), .B2(new_n859), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n834), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1045), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1047), .B1(new_n852), .B2(new_n854), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1051), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1028), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1023), .B(new_n1044), .C1(new_n1052), .C2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1033), .B(new_n1038), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1049), .A2(new_n1051), .A3(new_n1028), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1040), .A2(new_n862), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT121), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1030), .B1(new_n1062), .B2(new_n1041), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1058), .B(new_n1059), .C1(new_n1063), .C2(new_n1022), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1057), .A2(new_n1064), .A3(new_n667), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n781), .A2(new_n293), .ZN(new_n1067));
  INV_X1    g0867(.A(G125), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n302), .B1(new_n225), .B2(new_n728), .C1(new_n744), .C2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT122), .ZN(new_n1070));
  XOR2_X1   g0870(.A(KEYINPUT54), .B(G143), .Z(new_n1071));
  NAND2_X1  g0871(.A1(new_n741), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n729), .A2(new_n1003), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT53), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G128), .A2(new_n736), .B1(new_n747), .B2(G132), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n721), .A2(G137), .B1(new_n733), .B2(G159), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1070), .A2(new_n1072), .A3(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT123), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n729), .A2(new_n221), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n728), .A2(new_n202), .B1(new_n740), .B2(new_n427), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(G107), .C2(new_n721), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n745), .A2(G294), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n302), .B1(new_n733), .B2(G77), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G116), .A2(new_n747), .B1(new_n736), .B2(G283), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1079), .A2(new_n1086), .B1(new_n709), .B2(new_n710), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n777), .B(new_n1087), .C1(new_n1046), .C2(new_n712), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1066), .A2(new_n700), .B1(new_n1067), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1065), .A2(new_n1089), .ZN(G378));
  INV_X1    g0890(.A(KEYINPUT57), .ZN(new_n1091));
  OAI21_X1  g0891(.A(G330), .B1(new_n843), .B2(new_n847), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT125), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n402), .A2(KEYINPUT55), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n402), .A2(KEYINPUT55), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n391), .A2(new_n822), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT56), .Z(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1093), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1093), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1092), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1103), .B(G330), .C1(new_n843), .C2(new_n847), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1105), .A2(new_n864), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n864), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1022), .B1(new_n1066), .B2(new_n1044), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1091), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1057), .A2(new_n1023), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n864), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1105), .A2(new_n864), .A3(new_n1106), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1112), .A2(new_n1117), .A3(KEYINPUT57), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1111), .A2(new_n1118), .A3(new_n667), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n700), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1120));
  OR3_X1    g0920(.A1(new_n1100), .A2(new_n713), .A3(new_n1101), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n781), .A2(new_n225), .ZN(new_n1122));
  INV_X1    g0922(.A(G128), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1068), .A2(new_n735), .B1(new_n746), .B2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G132), .A2(new_n721), .B1(new_n741), .B2(G137), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1003), .B2(new_n732), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1124), .B(new_n1126), .C1(new_n784), .C2(new_n1071), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT59), .ZN(new_n1128));
  AOI21_X1  g0928(.A(G41), .B1(new_n888), .B2(G159), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT124), .B(G124), .ZN(new_n1130));
  AOI21_X1  g0930(.A(G33), .B1(new_n964), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G58), .A2(new_n888), .B1(new_n741), .B2(new_n603), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n202), .B2(new_n732), .C1(new_n427), .C2(new_n720), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n339), .B1(new_n729), .B2(new_n207), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1134), .A2(G41), .A3(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n745), .A2(G283), .B1(G116), .B2(new_n736), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(new_n428), .C2(new_n746), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT58), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n225), .B1(new_n266), .B2(G41), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1132), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n777), .B1(new_n1141), .B2(new_n711), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1121), .A2(new_n1122), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1120), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1119), .A2(new_n1145), .ZN(G375));
  NAND2_X1  g0946(.A1(new_n1044), .A2(new_n1023), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1022), .B(new_n1031), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n934), .A3(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G97), .A2(new_n784), .B1(new_n741), .B2(G107), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n489), .B2(new_n720), .ZN(new_n1151));
  NOR4_X1   g0951(.A1(new_n1151), .A2(new_n302), .A3(new_n881), .A4(new_n970), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n745), .A2(G303), .B1(G283), .B2(new_n747), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n961), .C2(new_n735), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n746), .A2(new_n797), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n732), .A2(new_n225), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n729), .A2(new_n757), .B1(new_n740), .B2(new_n1003), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(new_n721), .C2(new_n1071), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n745), .A2(G128), .B1(G132), .B2(new_n736), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n339), .B1(new_n888), .B2(G58), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1154), .B1(new_n1155), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n777), .B1(new_n1162), .B2(new_n711), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n859), .B2(new_n713), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n202), .B2(new_n781), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1044), .B2(new_n700), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1149), .A2(new_n1166), .ZN(G381));
  AND4_X1   g0967(.A1(new_n1089), .A2(new_n1065), .A3(new_n1120), .A4(new_n1143), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1119), .A2(new_n1168), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1169), .A2(G396), .A3(G393), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n931), .A2(new_n932), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n952), .B2(new_n700), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1172), .A2(new_n1016), .A3(new_n906), .A4(new_n1018), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1173), .A2(G384), .A3(G381), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(new_n1174), .ZN(G407));
  OAI211_X1 g0975(.A(G407), .B(G213), .C1(G343), .C2(new_n1169), .ZN(G409));
  NAND2_X1  g0976(.A1(G387), .A2(G390), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(G393), .B(G396), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1177), .A2(new_n1178), .A3(new_n1173), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n1177), .B2(new_n1173), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n643), .A2(G343), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(G2897), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n667), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1148), .A2(KEYINPUT126), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1186), .B2(KEYINPUT60), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT60), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1148), .A2(KEYINPUT126), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1187), .A2(new_n1147), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(G384), .A3(new_n1166), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(G384), .B1(new_n1190), .B2(new_n1166), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1184), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1190), .A2(new_n1166), .ZN(new_n1195));
  INV_X1    g0995(.A(G384), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1197), .A2(G2897), .A3(new_n1191), .A4(new_n1183), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT127), .ZN(new_n1200));
  INV_X1    g1000(.A(G378), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1119), .B2(new_n1145), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1065), .A2(new_n1120), .A3(new_n1089), .A4(new_n1143), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1109), .A2(new_n1110), .A3(new_n935), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1203), .A2(new_n1204), .B1(new_n643), .B2(G343), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1200), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1023), .A2(new_n1057), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n934), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1183), .B1(new_n1168), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1185), .B1(new_n1207), .B2(KEYINPUT57), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1144), .B1(new_n1210), .B2(new_n1111), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1209), .B(KEYINPUT127), .C1(new_n1211), .C2(new_n1201), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1199), .A2(new_n1206), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT61), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1202), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT62), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1209), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1213), .A2(new_n1214), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1206), .A2(new_n1212), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1217), .B1(new_n1220), .B2(new_n1216), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1182), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1215), .A2(new_n1216), .A3(new_n1209), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1215), .A2(new_n1209), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT63), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1220), .A2(KEYINPUT63), .A3(new_n1216), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n1214), .A4(new_n1181), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1222), .A2(new_n1228), .ZN(G405));
  NAND2_X1  g1029(.A1(new_n1215), .A2(new_n1169), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1181), .A2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1169), .B(new_n1215), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1216), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1216), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(G402));
endmodule


