

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  XNOR2_X2 U321 ( .A(n396), .B(n395), .ZN(n551) );
  XNOR2_X1 U322 ( .A(n306), .B(n442), .ZN(n526) );
  XNOR2_X1 U323 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U324 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U325 ( .A(n451), .B(G176GAT), .ZN(n452) );
  XNOR2_X1 U326 ( .A(n453), .B(n452), .ZN(G1349GAT) );
  XOR2_X1 U327 ( .A(G120GAT), .B(G71GAT), .Z(n402) );
  XOR2_X1 U328 ( .A(G127GAT), .B(KEYINPUT0), .Z(n290) );
  XNOR2_X1 U329 ( .A(G113GAT), .B(G134GAT), .ZN(n289) );
  XNOR2_X1 U330 ( .A(n290), .B(n289), .ZN(n329) );
  XOR2_X1 U331 ( .A(n402), .B(n329), .Z(n292) );
  XNOR2_X1 U332 ( .A(G43GAT), .B(G190GAT), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U334 ( .A(G15GAT), .B(KEYINPUT85), .Z(n294) );
  NAND2_X1 U335 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U337 ( .A(n296), .B(n295), .Z(n301) );
  XOR2_X1 U338 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n298) );
  XNOR2_X1 U339 ( .A(G99GAT), .B(G176GAT), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(n299), .ZN(n300) );
  XNOR2_X1 U342 ( .A(n301), .B(n300), .ZN(n306) );
  XOR2_X1 U343 ( .A(G183GAT), .B(KEYINPUT84), .Z(n303) );
  XNOR2_X1 U344 ( .A(KEYINPUT19), .B(KEYINPUT83), .ZN(n302) );
  XNOR2_X1 U345 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U346 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n304) );
  XNOR2_X1 U347 ( .A(n305), .B(n304), .ZN(n442) );
  XOR2_X1 U348 ( .A(KEYINPUT21), .B(G211GAT), .Z(n308) );
  XNOR2_X1 U349 ( .A(KEYINPUT86), .B(G204GAT), .ZN(n307) );
  XNOR2_X1 U350 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U351 ( .A(G197GAT), .B(n309), .Z(n438) );
  XOR2_X1 U352 ( .A(KEYINPUT3), .B(KEYINPUT87), .Z(n311) );
  XNOR2_X1 U353 ( .A(KEYINPUT88), .B(G155GAT), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U355 ( .A(KEYINPUT2), .B(n312), .Z(n328) );
  XNOR2_X1 U356 ( .A(n438), .B(n328), .ZN(n325) );
  XOR2_X1 U357 ( .A(KEYINPUT90), .B(G106GAT), .Z(n314) );
  XNOR2_X1 U358 ( .A(G50GAT), .B(G218GAT), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U360 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n316) );
  XNOR2_X1 U361 ( .A(KEYINPUT23), .B(KEYINPUT89), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U363 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U364 ( .A(G141GAT), .B(G22GAT), .Z(n348) );
  XOR2_X1 U365 ( .A(G148GAT), .B(G78GAT), .Z(n401) );
  XOR2_X1 U366 ( .A(KEYINPUT75), .B(G162GAT), .Z(n390) );
  XOR2_X1 U367 ( .A(n401), .B(n390), .Z(n320) );
  NAND2_X1 U368 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n348), .B(n321), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n461) );
  XOR2_X1 U373 ( .A(KEYINPUT92), .B(KEYINPUT1), .Z(n327) );
  XNOR2_X1 U374 ( .A(G1GAT), .B(G57GAT), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n333) );
  XOR2_X1 U376 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n331) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U379 ( .A(n333), .B(n332), .ZN(n345) );
  NAND2_X1 U380 ( .A1(G225GAT), .A2(G233GAT), .ZN(n339) );
  XOR2_X1 U381 ( .A(G85GAT), .B(G148GAT), .Z(n335) );
  XNOR2_X1 U382 ( .A(G141GAT), .B(G120GAT), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n337) );
  XOR2_X1 U384 ( .A(G29GAT), .B(G162GAT), .Z(n336) );
  XNOR2_X1 U385 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U386 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U387 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n341) );
  XNOR2_X1 U388 ( .A(KEYINPUT94), .B(KEYINPUT91), .ZN(n340) );
  XNOR2_X1 U389 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U390 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U391 ( .A(n345), .B(n344), .ZN(n524) );
  XOR2_X1 U392 ( .A(G169GAT), .B(G8GAT), .Z(n439) );
  XOR2_X1 U393 ( .A(G15GAT), .B(G1GAT), .Z(n366) );
  XOR2_X1 U394 ( .A(n439), .B(n366), .Z(n347) );
  NAND2_X1 U395 ( .A1(G229GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U396 ( .A(n347), .B(n346), .ZN(n349) );
  XOR2_X1 U397 ( .A(n349), .B(n348), .Z(n357) );
  XOR2_X1 U398 ( .A(KEYINPUT66), .B(KEYINPUT64), .Z(n351) );
  XNOR2_X1 U399 ( .A(G197GAT), .B(G113GAT), .ZN(n350) );
  XNOR2_X1 U400 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U401 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n353) );
  XNOR2_X1 U402 ( .A(KEYINPUT67), .B(KEYINPUT65), .ZN(n352) );
  XNOR2_X1 U403 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U404 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U405 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U406 ( .A(G29GAT), .B(KEYINPUT8), .Z(n359) );
  XNOR2_X1 U407 ( .A(G43GAT), .B(G36GAT), .ZN(n358) );
  XNOR2_X1 U408 ( .A(n359), .B(n358), .ZN(n361) );
  XOR2_X1 U409 ( .A(G50GAT), .B(KEYINPUT7), .Z(n360) );
  XNOR2_X1 U410 ( .A(n361), .B(n360), .ZN(n382) );
  XNOR2_X1 U411 ( .A(n362), .B(n382), .ZN(n564) );
  XNOR2_X1 U412 ( .A(n564), .B(KEYINPUT68), .ZN(n553) );
  XOR2_X1 U413 ( .A(G78GAT), .B(G211GAT), .Z(n364) );
  XNOR2_X1 U414 ( .A(G183GAT), .B(G127GAT), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U416 ( .A(n365), .B(G155GAT), .Z(n368) );
  XNOR2_X1 U417 ( .A(G22GAT), .B(n366), .ZN(n367) );
  XNOR2_X1 U418 ( .A(n368), .B(n367), .ZN(n381) );
  XOR2_X1 U419 ( .A(KEYINPUT81), .B(KEYINPUT12), .Z(n370) );
  NAND2_X1 U420 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U422 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n372) );
  XNOR2_X1 U423 ( .A(KEYINPUT80), .B(KEYINPUT78), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U425 ( .A(n374), .B(n373), .Z(n379) );
  XOR2_X1 U426 ( .A(G57GAT), .B(KEYINPUT13), .Z(n400) );
  XOR2_X1 U427 ( .A(KEYINPUT79), .B(G64GAT), .Z(n376) );
  XNOR2_X1 U428 ( .A(G8GAT), .B(G71GAT), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U430 ( .A(n400), .B(n377), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U432 ( .A(n381), .B(n380), .Z(n573) );
  INV_X1 U433 ( .A(n573), .ZN(n481) );
  INV_X1 U434 ( .A(KEYINPUT36), .ZN(n397) );
  INV_X1 U435 ( .A(n382), .ZN(n396) );
  XOR2_X1 U436 ( .A(G92GAT), .B(G85GAT), .Z(n384) );
  XNOR2_X1 U437 ( .A(G99GAT), .B(G106GAT), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n405) );
  INV_X1 U439 ( .A(KEYINPUT10), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n405), .B(n385), .ZN(n387) );
  NAND2_X1 U441 ( .A1(G232GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n394) );
  XOR2_X1 U443 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n389) );
  XNOR2_X1 U444 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n388) );
  XOR2_X1 U445 ( .A(n389), .B(n388), .Z(n392) );
  XOR2_X1 U446 ( .A(G190GAT), .B(G218GAT), .Z(n431) );
  XNOR2_X1 U447 ( .A(n390), .B(n431), .ZN(n391) );
  XOR2_X2 U448 ( .A(KEYINPUT77), .B(n551), .Z(n536) );
  XNOR2_X1 U449 ( .A(n397), .B(n536), .ZN(n479) );
  NOR2_X1 U450 ( .A1(n481), .A2(n479), .ZN(n398) );
  XOR2_X1 U451 ( .A(KEYINPUT45), .B(n398), .Z(n399) );
  NOR2_X1 U452 ( .A1(n553), .A2(n399), .ZN(n418) );
  XOR2_X1 U453 ( .A(G176GAT), .B(G64GAT), .Z(n430) );
  XOR2_X1 U454 ( .A(n400), .B(n430), .Z(n404) );
  XNOR2_X1 U455 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U456 ( .A(n404), .B(n403), .ZN(n409) );
  XOR2_X1 U457 ( .A(n405), .B(KEYINPUT70), .Z(n407) );
  NAND2_X1 U458 ( .A1(G230GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U459 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U460 ( .A(n409), .B(n408), .Z(n417) );
  XOR2_X1 U461 ( .A(KEYINPUT71), .B(KEYINPUT69), .Z(n411) );
  XNOR2_X1 U462 ( .A(G204GAT), .B(KEYINPUT73), .ZN(n410) );
  XNOR2_X1 U463 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U464 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n413) );
  XNOR2_X1 U465 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n412) );
  XNOR2_X1 U466 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n417), .B(n416), .ZN(n569) );
  NAND2_X1 U469 ( .A1(n418), .A2(n569), .ZN(n419) );
  XNOR2_X1 U470 ( .A(n419), .B(KEYINPUT112), .ZN(n428) );
  XNOR2_X1 U471 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n426) );
  XOR2_X1 U472 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n421) );
  XOR2_X1 U473 ( .A(KEYINPUT41), .B(n569), .Z(n494) );
  INV_X1 U474 ( .A(n494), .ZN(n545) );
  NAND2_X1 U475 ( .A1(n564), .A2(n545), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n423) );
  NOR2_X1 U477 ( .A1(n551), .A2(n573), .ZN(n422) );
  NAND2_X1 U478 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(KEYINPUT47), .B(n424), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n427) );
  NAND2_X1 U481 ( .A1(n428), .A2(n427), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n429), .B(KEYINPUT48), .ZN(n522) );
  XOR2_X1 U483 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U484 ( .A1(G226GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U486 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n435) );
  XNOR2_X1 U487 ( .A(G36GAT), .B(G92GAT), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U489 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U491 ( .A(n441), .B(n440), .ZN(n443) );
  XNOR2_X1 U492 ( .A(n443), .B(n442), .ZN(n457) );
  NAND2_X1 U493 ( .A1(n522), .A2(n457), .ZN(n445) );
  XOR2_X1 U494 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n444) );
  XNOR2_X1 U495 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U496 ( .A1(n524), .A2(n446), .ZN(n562) );
  NOR2_X1 U497 ( .A1(n461), .A2(n562), .ZN(n448) );
  XNOR2_X1 U498 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U500 ( .A(KEYINPUT119), .B(n449), .Z(n450) );
  NOR2_X2 U501 ( .A1(n526), .A2(n450), .ZN(n557) );
  NAND2_X1 U502 ( .A1(n557), .A2(n545), .ZN(n453) );
  XOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n451) );
  INV_X1 U504 ( .A(n524), .ZN(n456) );
  XOR2_X1 U505 ( .A(n457), .B(KEYINPUT27), .Z(n523) );
  XNOR2_X1 U506 ( .A(n461), .B(KEYINPUT28), .ZN(n529) );
  NOR2_X1 U507 ( .A1(n523), .A2(n529), .ZN(n454) );
  NAND2_X1 U508 ( .A1(n454), .A2(n526), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n456), .A2(n455), .ZN(n467) );
  INV_X1 U510 ( .A(n457), .ZN(n513) );
  OR2_X1 U511 ( .A1(n513), .A2(n526), .ZN(n458) );
  XNOR2_X1 U512 ( .A(KEYINPUT97), .B(n458), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n461), .A2(n459), .ZN(n460) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n460), .Z(n464) );
  NAND2_X1 U515 ( .A1(n461), .A2(n526), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n462), .B(KEYINPUT26), .ZN(n563) );
  NOR2_X1 U517 ( .A1(n523), .A2(n563), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n524), .A2(n465), .ZN(n466) );
  NAND2_X1 U520 ( .A1(n467), .A2(n466), .ZN(n480) );
  NOR2_X1 U521 ( .A1(n481), .A2(n536), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT16), .B(n468), .Z(n469) );
  NOR2_X1 U523 ( .A1(n480), .A2(n469), .ZN(n495) );
  NAND2_X1 U524 ( .A1(n553), .A2(n569), .ZN(n470) );
  XOR2_X1 U525 ( .A(KEYINPUT74), .B(n470), .Z(n484) );
  NAND2_X1 U526 ( .A1(n495), .A2(n484), .ZN(n476) );
  NOR2_X1 U527 ( .A1(n524), .A2(n476), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT34), .B(n471), .Z(n472) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n472), .ZN(G1324GAT) );
  NOR2_X1 U530 ( .A1(n513), .A2(n476), .ZN(n473) );
  XOR2_X1 U531 ( .A(G8GAT), .B(n473), .Z(G1325GAT) );
  NOR2_X1 U532 ( .A1(n526), .A2(n476), .ZN(n475) );
  XNOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  INV_X1 U535 ( .A(n529), .ZN(n519) );
  NOR2_X1 U536 ( .A1(n519), .A2(n476), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT98), .B(n477), .Z(n478) );
  XNOR2_X1 U538 ( .A(G22GAT), .B(n478), .ZN(G1327GAT) );
  XNOR2_X1 U539 ( .A(KEYINPUT99), .B(KEYINPUT39), .ZN(n487) );
  NOR2_X1 U540 ( .A1(n479), .A2(n480), .ZN(n482) );
  NAND2_X1 U541 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(n483), .ZN(n510) );
  NAND2_X1 U543 ( .A1(n484), .A2(n510), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(KEYINPUT38), .ZN(n492) );
  NOR2_X1 U545 ( .A1(n524), .A2(n492), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U547 ( .A(G29GAT), .B(n488), .Z(G1328GAT) );
  NOR2_X1 U548 ( .A1(n492), .A2(n513), .ZN(n489) );
  XOR2_X1 U549 ( .A(G36GAT), .B(n489), .Z(G1329GAT) );
  NOR2_X1 U550 ( .A1(n526), .A2(n492), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT40), .B(n490), .Z(n491) );
  XNOR2_X1 U552 ( .A(G43GAT), .B(n491), .ZN(G1330GAT) );
  NOR2_X1 U553 ( .A1(n519), .A2(n492), .ZN(n493) );
  XOR2_X1 U554 ( .A(G50GAT), .B(n493), .Z(G1331GAT) );
  NOR2_X1 U555 ( .A1(n564), .A2(n494), .ZN(n509) );
  NAND2_X1 U556 ( .A1(n509), .A2(n495), .ZN(n505) );
  NOR2_X1 U557 ( .A1(n524), .A2(n505), .ZN(n497) );
  XNOR2_X1 U558 ( .A(KEYINPUT42), .B(KEYINPUT100), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U560 ( .A(G57GAT), .B(n498), .Z(G1332GAT) );
  NOR2_X1 U561 ( .A1(n513), .A2(n505), .ZN(n500) );
  XNOR2_X1 U562 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(n501), .ZN(G1333GAT) );
  NOR2_X1 U565 ( .A1(n526), .A2(n505), .ZN(n503) );
  XNOR2_X1 U566 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G71GAT), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U569 ( .A1(n519), .A2(n505), .ZN(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U572 ( .A(G78GAT), .B(n508), .Z(G1335GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n509), .ZN(n518) );
  NOR2_X1 U574 ( .A1(n524), .A2(n518), .ZN(n511) );
  XOR2_X1 U575 ( .A(G85GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT106), .B(n512), .ZN(G1336GAT) );
  NOR2_X1 U577 ( .A1(n513), .A2(n518), .ZN(n514) );
  XOR2_X1 U578 ( .A(G92GAT), .B(n514), .Z(G1337GAT) );
  NOR2_X1 U579 ( .A1(n526), .A2(n518), .ZN(n515) );
  XOR2_X1 U580 ( .A(G99GAT), .B(n515), .Z(G1338GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n517) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(KEYINPUT108), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(n521) );
  NOR2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U585 ( .A(n521), .B(n520), .Z(G1339GAT) );
  NOR2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U587 ( .A1(n522), .A2(n525), .ZN(n540) );
  NOR2_X1 U588 ( .A1(n526), .A2(n540), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(KEYINPUT113), .ZN(n528) );
  NOR2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n553), .A2(n537), .ZN(n530) );
  XNOR2_X1 U592 ( .A(n530), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n532) );
  NAND2_X1 U594 ( .A1(n537), .A2(n545), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(n533), .ZN(G1341GAT) );
  NAND2_X1 U597 ( .A1(n537), .A2(n573), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NOR2_X1 U603 ( .A1(n563), .A2(n540), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n564), .A2(n550), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(n541), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n543) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT52), .B(n544), .Z(n547) );
  NAND2_X1 U610 ( .A1(n550), .A2(n545), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  XOR2_X1 U612 ( .A(G155GAT), .B(KEYINPUT117), .Z(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n573), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1346GAT) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n552), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U617 ( .A(G169GAT), .B(KEYINPUT121), .Z(n555) );
  NAND2_X1 U618 ( .A1(n557), .A2(n553), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(G1348GAT) );
  NAND2_X1 U620 ( .A1(n557), .A2(n573), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n536), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(KEYINPUT58), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n561) );
  XNOR2_X1 U626 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n568) );
  XOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT59), .Z(n566) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n574), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n571) );
  INV_X1 U634 ( .A(n574), .ZN(n578) );
  OR2_X1 U635 ( .A1(n578), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n577) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n580) );
  NOR2_X1 U643 ( .A1(n479), .A2(n578), .ZN(n579) );
  XOR2_X1 U644 ( .A(n580), .B(n579), .Z(G1355GAT) );
endmodule

