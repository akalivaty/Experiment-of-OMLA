//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954;
  XNOR2_X1  g000(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n203), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n203), .B1(KEYINPUT66), .B2(G183gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n202), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT28), .A3(new_n205), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NOR3_X1   g015(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n212), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221));
  INV_X1    g020(.A(G169gat), .ZN(new_n222));
  INV_X1    g021(.A(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT23), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n212), .A2(KEYINPUT24), .ZN(new_n227));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n224), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n231), .A2(new_n233), .A3(KEYINPUT25), .A4(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n221), .B1(new_n229), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n213), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n229), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n229), .A2(new_n235), .A3(new_n221), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n220), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G134gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(KEYINPUT68), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(KEYINPUT1), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247));
  INV_X1    g046(.A(G113gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(G120gat), .ZN(new_n249));
  INV_X1    g048(.A(G120gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(G113gat), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n247), .B(new_n243), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G127gat), .ZN(new_n254));
  INV_X1    g053(.A(G127gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n246), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n257), .ZN(new_n258));
  AND4_X1   g057(.A1(KEYINPUT25), .A2(new_n231), .A3(new_n233), .A4(new_n234), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n227), .A2(new_n228), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n224), .A2(new_n226), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n259), .A2(KEYINPUT65), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(new_n239), .A3(new_n236), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n263), .A2(new_n254), .A3(new_n256), .A4(new_n220), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G227gat), .ZN(new_n266));
  INV_X1    g065(.A(G233gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT34), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT32), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n266), .A2(new_n267), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n258), .A2(new_n271), .A3(new_n264), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n271), .A4(new_n264), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT33), .B1(new_n274), .B2(new_n275), .ZN(new_n277));
  XNOR2_X1  g076(.A(G15gat), .B(G43gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(G71gat), .B(G99gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n276), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n280), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n283), .A2(KEYINPUT33), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n276), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n269), .B1(new_n281), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT83), .B(G22gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G228gat), .A2(G233gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT22), .ZN(new_n294));
  INV_X1    g093(.A(G211gat), .ZN(new_n295));
  INV_X1    g094(.A(G218gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G211gat), .B(G218gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n293), .A3(new_n297), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n304));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  INV_X1    g105(.A(G141gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(G148gat), .ZN(new_n308));
  INV_X1    g107(.A(G148gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(G141gat), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n304), .B(new_n306), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G155gat), .B(G162gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G141gat), .B(G148gat), .Z(new_n315));
  NAND4_X1  g114(.A1(new_n315), .A2(new_n312), .A3(new_n304), .A4(new_n306), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT77), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT77), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n314), .A2(new_n316), .A3(new_n320), .A4(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n303), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n314), .A2(new_n316), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT78), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT29), .B1(new_n301), .B2(new_n302), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n324), .A2(KEYINPUT80), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n333));
  AOI211_X1 g132(.A(new_n333), .B(new_n303), .C1(new_n322), .C2(new_n323), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n292), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G78gat), .B(G106gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT31), .B(G50gat), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n336), .B(new_n337), .Z(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n314), .A2(new_n316), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT81), .B1(new_n331), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n345), .B(new_n325), .C1(new_n330), .C2(KEYINPUT3), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n292), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n322), .A2(new_n323), .ZN(new_n348));
  INV_X1    g147(.A(new_n303), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n347), .A2(new_n350), .B1(new_n340), .B2(new_n339), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n335), .A2(new_n342), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n342), .B1(new_n335), .B2(new_n351), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n291), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n274), .A2(new_n275), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT32), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT33), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n358), .A3(new_n282), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n268), .B(KEYINPUT34), .Z(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n360), .A3(new_n287), .ZN(new_n361));
  INV_X1    g160(.A(new_n292), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n329), .A2(new_n331), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n350), .B2(new_n333), .ZN(new_n364));
  INV_X1    g163(.A(new_n334), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n351), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n341), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n335), .A2(new_n342), .A3(new_n351), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n290), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n289), .A2(new_n354), .A3(new_n361), .A4(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n317), .B1(new_n314), .B2(new_n316), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n246), .A2(new_n252), .A3(new_n255), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n255), .B1(new_n246), .B2(new_n252), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n322), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n257), .A2(new_n327), .A3(KEYINPUT4), .A4(new_n328), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n343), .B1(new_n374), .B2(new_n373), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n376), .A2(new_n377), .A3(new_n378), .A4(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n254), .A2(new_n325), .A3(new_n256), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n377), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT0), .ZN(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  NAND2_X1  g191(.A1(new_n379), .A2(KEYINPUT4), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n257), .A2(new_n327), .A3(new_n380), .A4(new_n328), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n395), .A2(new_n383), .A3(new_n377), .A4(new_n376), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n388), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n388), .A2(new_n396), .ZN(new_n400));
  INV_X1    g199(.A(new_n392), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n388), .A2(KEYINPUT79), .A3(new_n392), .A4(new_n396), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n399), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(KEYINPUT6), .A3(new_n401), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n263), .A2(new_n408), .A3(new_n220), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n263), .B2(new_n220), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n349), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n263), .A2(new_n408), .A3(new_n220), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n218), .B1(new_n208), .B2(new_n210), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n236), .A2(new_n239), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(new_n262), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n303), .B(new_n413), .C1(new_n416), .C2(new_n410), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n417), .A3(KEYINPUT71), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n409), .A2(new_n411), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT71), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n303), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(KEYINPUT30), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT75), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n418), .B2(new_n421), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT75), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT30), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n431), .A2(KEYINPUT30), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n422), .A2(KEYINPUT72), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT72), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n437), .A3(new_n421), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n435), .B1(new_n439), .B2(new_n427), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n407), .A2(new_n434), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT35), .B1(new_n371), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n444));
  AOI211_X1 g243(.A(KEYINPUT5), .B(new_n386), .C1(new_n322), .C2(new_n375), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n382), .A2(new_n387), .B1(new_n445), .B2(new_n395), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n446), .B2(new_n392), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n400), .A2(KEYINPUT86), .A3(new_n401), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n406), .B1(new_n443), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT35), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(new_n371), .ZN(new_n453));
  INV_X1    g252(.A(new_n438), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n437), .B1(new_n418), .B2(new_n421), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n427), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n435), .ZN(new_n457));
  INV_X1    g256(.A(new_n433), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n432), .B1(new_n431), .B2(KEYINPUT30), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n440), .A2(KEYINPUT84), .A3(new_n434), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g263(.A1(KEYINPUT88), .A2(new_n442), .B1(new_n453), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n466), .B(KEYINPUT35), .C1(new_n371), .C2(new_n441), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT39), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n385), .A2(new_n386), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(KEYINPUT85), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n395), .A2(new_n376), .ZN(new_n471));
  OAI221_X1 g270(.A(new_n470), .B1(KEYINPUT85), .B2(new_n469), .C1(new_n471), .C2(new_n377), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n377), .B1(new_n395), .B2(new_n376), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n401), .B1(new_n473), .B2(new_n468), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT40), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n449), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n354), .A2(new_n370), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n431), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n406), .B(new_n483), .C1(new_n443), .C2(new_n449), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n436), .B2(new_n438), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n422), .A2(new_n485), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n427), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT38), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n412), .A2(new_n417), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT38), .B1(new_n490), .B2(KEYINPUT37), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n487), .A2(new_n427), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n492), .A2(new_n493), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n489), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n480), .B(new_n482), .C1(new_n484), .C2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  INV_X1    g297(.A(new_n361), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n360), .B1(new_n359), .B2(new_n287), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n289), .A2(KEYINPUT36), .A3(new_n361), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n501), .A2(new_n502), .B1(new_n441), .B2(new_n481), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n465), .A2(new_n467), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G43gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G50gat), .ZN(new_n506));
  INV_X1    g305(.A(G50gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G43gat), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT15), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT14), .B(G29gat), .Z(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(G36gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT14), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n512), .A2(new_n513), .A3(G29gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n509), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n511), .A2(new_n514), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT90), .B(G50gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n505), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT91), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT91), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n520), .A3(new_n505), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n508), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n515), .B1(new_n524), .B2(new_n509), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT17), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(G1gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(G1gat), .B2(new_n527), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G8gat), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n529), .B(new_n532), .C1(G1gat), .C2(new_n527), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n509), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n518), .A2(KEYINPUT91), .B1(G43gat), .B2(new_n507), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT15), .B1(new_n537), .B2(new_n521), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n538), .B2(new_n516), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n540), .A3(new_n515), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n535), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n534), .B(new_n515), .C1(new_n524), .C2(new_n509), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT92), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n539), .A2(new_n545), .A3(new_n534), .A4(new_n515), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT93), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT18), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n542), .A2(new_n547), .A3(new_n552), .A4(new_n548), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n542), .A2(new_n547), .A3(new_n548), .ZN(new_n555));
  INV_X1    g354(.A(new_n525), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n547), .B1(new_n534), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n548), .B(KEYINPUT13), .Z(new_n558));
  AOI22_X1  g357(.A1(new_n555), .A2(KEYINPUT18), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G113gat), .B(G141gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G169gat), .B(G197gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT12), .Z(new_n568));
  NAND3_X1  g367(.A1(new_n560), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n554), .B(new_n559), .C1(new_n561), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n504), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n407), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT95), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n582), .B(KEYINPUT95), .C1(new_n578), .C2(new_n577), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n586), .A2(KEYINPUT21), .ZN(new_n587));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(new_n255), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n584), .A2(KEYINPUT96), .A3(new_n585), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT96), .B1(new_n584), .B2(new_n585), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT21), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(new_n593), .A3(new_n535), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n589), .B(G127gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n535), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT97), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  INV_X1    g400(.A(G155gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n600), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n594), .A2(new_n597), .A3(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT8), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(G85gat), .B2(G92gat), .ZN(new_n614));
  XOR2_X1   g413(.A(G99gat), .B(G106gat), .Z(new_n615));
  OR3_X1    g414(.A1(new_n611), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(new_n611), .B2(new_n614), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n556), .A2(new_n618), .B1(KEYINPUT41), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n617), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT100), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n526), .A2(new_n541), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G190gat), .B(G218gat), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n620), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n620), .B2(new_n623), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n619), .A2(KEYINPUT41), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT98), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n626), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n626), .B2(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n615), .A2(KEYINPUT101), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n586), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n621), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n586), .A2(new_n616), .A3(new_n617), .A4(new_n636), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n644), .A3(new_n639), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n618), .B(KEYINPUT10), .C1(new_n591), .C2(new_n592), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT102), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n608), .A2(new_n635), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n576), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT103), .B(G1gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1324gat));
  INV_X1    g459(.A(new_n464), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  NAND4_X1  g461(.A1(new_n574), .A2(new_n656), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n574), .A2(new_n656), .A3(new_n661), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n664), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT104), .B1(new_n664), .B2(KEYINPUT42), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n663), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT105), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n666), .A2(new_n667), .A3(new_n673), .A4(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(G1325gat));
  NOR3_X1   g474(.A1(new_n504), .A2(new_n657), .A3(new_n573), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n501), .A2(new_n502), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n499), .A2(new_n500), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n504), .A2(new_n573), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n657), .A2(G15gat), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n679), .A2(G15gat), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT106), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n676), .A2(new_n481), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT107), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT43), .B(G22gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  NOR2_X1   g488(.A1(new_n608), .A2(new_n635), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n655), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n576), .A2(G29gat), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT45), .Z(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(new_n504), .B2(new_n635), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n442), .A2(KEYINPUT88), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n453), .A2(new_n464), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n467), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n480), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n482), .B1(new_n496), .B2(new_n484), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n503), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n635), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(KEYINPUT44), .A3(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n698), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n608), .B(KEYINPUT108), .Z(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n692), .A3(new_n573), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n575), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G29gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n712), .ZN(G1328gat));
  NAND3_X1  g512(.A1(new_n708), .A2(new_n661), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G36gat), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n574), .A2(new_n513), .A3(new_n661), .A4(new_n693), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n715), .A2(new_n718), .A3(KEYINPUT109), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1329gat));
  NAND4_X1  g522(.A1(new_n698), .A2(new_n678), .A3(new_n707), .A4(new_n710), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n694), .A2(G43gat), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n724), .A2(G43gat), .B1(new_n682), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1330gat));
  NAND4_X1  g529(.A1(new_n698), .A2(new_n481), .A3(new_n707), .A4(new_n710), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n517), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n482), .A2(new_n517), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n693), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n574), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g538(.A1(new_n705), .A2(new_n573), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n608), .A2(new_n635), .A3(new_n692), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n575), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n661), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT49), .B(G64gat), .Z(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n745), .B2(new_n747), .ZN(G1333gat));
  NOR4_X1   g547(.A1(new_n740), .A2(G71gat), .A3(new_n681), .A4(new_n741), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(G71gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n740), .A2(new_n677), .A3(new_n741), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n750), .B(KEYINPUT113), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n752), .A2(new_n751), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(new_n749), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n753), .A2(new_n756), .A3(new_n758), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n742), .A2(new_n481), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g563(.A1(new_n572), .A2(new_n608), .A3(new_n655), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n708), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n407), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n573), .A4(new_n690), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n705), .A2(new_n573), .A3(new_n690), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n572), .B1(new_n701), .B2(new_n704), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n774), .A2(KEYINPUT114), .A3(KEYINPUT51), .A4(new_n690), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n770), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n407), .A2(G85gat), .A3(new_n655), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n767), .B1(new_n777), .B2(new_n778), .ZN(G1336gat));
  NOR3_X1   g578(.A1(new_n464), .A2(G92gat), .A3(new_n655), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n698), .A2(new_n661), .A3(new_n707), .A4(new_n765), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(new_n782), .B2(G92gat), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n773), .A2(new_n768), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n780), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(G92gat), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT115), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n781), .A2(new_n783), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n787), .A2(new_n788), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(new_n785), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n794), .ZN(G1337gat));
  OAI21_X1  g594(.A(G99gat), .B1(new_n766), .B2(new_n677), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n681), .A2(G99gat), .A3(new_n655), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n777), .B2(new_n797), .ZN(G1338gat));
  NAND3_X1  g597(.A1(new_n708), .A2(new_n481), .A3(new_n765), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G106gat), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n482), .A2(G106gat), .A3(new_n655), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n776), .A2(new_n803), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n799), .A2(G106gat), .B1(new_n786), .B2(new_n803), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n802), .A2(new_n804), .B1(new_n805), .B2(new_n801), .ZN(G1339gat));
  NOR2_X1   g605(.A1(new_n657), .A2(new_n572), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n645), .A2(new_n646), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n641), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n645), .A2(new_n646), .A3(new_n643), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n651), .B1(new_n647), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT117), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT55), .B1(new_n811), .B2(new_n813), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n809), .B(new_n651), .C1(new_n641), .C2(new_n640), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n822), .B1(new_n821), .B2(new_n823), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n817), .B(new_n820), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n548), .B1(new_n542), .B2(new_n547), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n828), .A2(new_n829), .B1(new_n557), .B2(new_n558), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n567), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n554), .A2(new_n559), .A3(new_n570), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n827), .A2(new_n706), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n692), .A2(new_n833), .A3(new_n832), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n827), .B2(new_n572), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n836), .B2(new_n706), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n608), .B(KEYINPUT108), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n807), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n680), .A2(new_n482), .A3(new_n575), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n839), .A2(new_n661), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n572), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g642(.A1(new_n692), .A2(new_n250), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT119), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n841), .A2(new_n692), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n250), .ZN(G1341gat));
  NAND2_X1  g647(.A1(new_n841), .A2(new_n608), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT68), .B(G127gat), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n838), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n849), .A2(new_n850), .B1(new_n841), .B2(new_n851), .ZN(G1342gat));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n841), .B(new_n706), .C1(new_n853), .C2(new_n243), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n243), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1343gat));
  NOR3_X1   g655(.A1(new_n678), .A2(new_n661), .A3(new_n407), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n858), .B(new_n859), .C1(new_n839), .C2(new_n482), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n816), .A2(new_n823), .A3(new_n821), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n569), .B2(new_n571), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n635), .B1(new_n862), .B2(new_n835), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n608), .B1(new_n863), .B2(new_n834), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT57), .B(new_n481), .C1(new_n864), .C2(new_n807), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n826), .B1(new_n571), .B2(new_n569), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n635), .B1(new_n867), .B2(new_n835), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n709), .B1(new_n868), .B2(new_n834), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n481), .B1(new_n869), .B2(new_n807), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n858), .B1(new_n870), .B2(new_n859), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n572), .B(new_n857), .C1(new_n866), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G141gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n677), .A2(new_n481), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n575), .B(new_n464), .C1(new_n874), .C2(KEYINPUT121), .ZN(new_n875));
  AOI211_X1 g674(.A(new_n875), .B(new_n839), .C1(KEYINPUT121), .C2(new_n874), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n573), .A2(G141gat), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT122), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n873), .A2(new_n881), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1344gat));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n857), .B1(new_n866), .B2(new_n871), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n884), .B(G148gat), .C1(new_n885), .C2(new_n655), .ZN(new_n886));
  INV_X1    g685(.A(new_n870), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n481), .B1(new_n864), .B2(new_n807), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n859), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n857), .A2(new_n692), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n309), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n886), .B1(new_n884), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n876), .A2(new_n309), .A3(new_n692), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1345gat));
  OAI21_X1  g695(.A(G155gat), .B1(new_n885), .B2(new_n838), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n602), .A3(new_n608), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1346gat));
  OAI211_X1 g698(.A(new_n706), .B(new_n857), .C1(new_n866), .C2(new_n871), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G162gat), .ZN(new_n901));
  INV_X1    g700(.A(G162gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n876), .A2(new_n902), .A3(new_n706), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n901), .A2(KEYINPUT123), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1347gat));
  NAND2_X1  g707(.A1(new_n661), .A2(new_n407), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n371), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n869), .B2(new_n807), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n222), .A3(new_n573), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n572), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n912), .B1(new_n916), .B2(new_n222), .ZN(G1348gat));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n223), .A3(new_n692), .ZN(new_n918));
  OAI21_X1  g717(.A(G176gat), .B1(new_n911), .B2(new_n655), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1349gat));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(new_n911), .B2(new_n838), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G183gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n911), .A2(new_n921), .A3(new_n838), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n608), .A2(new_n209), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n923), .A2(new_n924), .B1(new_n911), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g726(.A1(new_n913), .A2(new_n205), .A3(new_n706), .A4(new_n914), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT126), .Z(new_n929));
  OAI21_X1  g728(.A(G190gat), .B1(new_n911), .B2(new_n635), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n909), .A2(new_n678), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n887), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n572), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n933), .B(KEYINPUT127), .Z(new_n937));
  AOI21_X1  g736(.A(new_n937), .B1(new_n888), .B2(new_n890), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n572), .A2(G197gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  INV_X1    g739(.A(new_n938), .ZN(new_n941));
  OAI21_X1  g740(.A(G204gat), .B1(new_n941), .B2(new_n655), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n934), .A2(G204gat), .A3(new_n655), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n935), .A2(new_n295), .A3(new_n608), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n938), .A2(new_n608), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1354gat));
  OAI21_X1  g751(.A(G218gat), .B1(new_n941), .B2(new_n635), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n935), .A2(new_n296), .A3(new_n706), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1355gat));
endmodule


