//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n187));
  OAI21_X1  g001(.A(G214), .B1(G237), .B2(G902), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G122), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT3), .A2(G107), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT3), .A2(G107), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(G104), .B2(new_n194), .ZN(new_n195));
  OR2_X1    g009(.A1(KEYINPUT77), .A2(G104), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT77), .A2(G104), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n195), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n196), .A2(new_n198), .A3(new_n200), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n202), .B1(G104), .B2(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G113), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT66), .A2(G119), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT66), .A2(G119), .ZN(new_n210));
  INV_X1    g024(.A(G116), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT5), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n208), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT66), .A2(G119), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(G116), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n216), .A2(G116), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(KEYINPUT5), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n212), .A2(new_n220), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT2), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G113), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n214), .A2(new_n222), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n229));
  INV_X1    g043(.A(new_n200), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT77), .A2(G104), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n230), .A2(new_n231), .A3(new_n194), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G107), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n199), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(G101), .B(new_n229), .C1(new_n232), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n202), .B1(new_n195), .B2(new_n201), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT79), .A3(new_n229), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n195), .A2(new_n201), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G101), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n238), .A2(new_n240), .B1(new_n243), .B2(new_n203), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n224), .A2(new_n226), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n212), .B2(new_n220), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n219), .A2(new_n221), .A3(new_n227), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(KEYINPUT67), .B(new_n245), .C1(new_n212), .C2(new_n220), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI221_X4 g065(.A(new_n192), .B1(new_n207), .B2(new_n228), .C1(new_n244), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n238), .A2(new_n240), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n242), .A2(G101), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n253), .A2(new_n250), .A3(new_n249), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n228), .A2(new_n207), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n191), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n190), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n236), .A2(new_n237), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT79), .B1(new_n239), .B2(new_n229), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n249), .A2(new_n250), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n257), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n192), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n189), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT83), .ZN(new_n267));
  INV_X1    g081(.A(G143), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT64), .B1(new_n268), .B2(G146), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n270));
  INV_X1    g084(.A(G146), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G143), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n268), .A2(G146), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n269), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(G143), .B(G146), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n279), .A2(new_n275), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n267), .B(G125), .C1(new_n278), .C2(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n274), .A2(new_n277), .B1(new_n279), .B2(new_n275), .ZN(new_n282));
  INV_X1    g096(.A(G125), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT83), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT84), .ZN(new_n286));
  INV_X1    g100(.A(G953), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G224), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n288), .B(KEYINPUT85), .Z(new_n289));
  INV_X1    g103(.A(KEYINPUT84), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n281), .A2(new_n284), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n268), .A2(G146), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n293));
  OAI21_X1  g107(.A(G128), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G128), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(KEYINPUT1), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n274), .A2(new_n294), .B1(new_n279), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n283), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n286), .A2(new_n289), .A3(new_n291), .A4(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n286), .A2(new_n291), .A3(new_n298), .ZN(new_n300));
  INV_X1    g114(.A(new_n289), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n259), .A2(new_n266), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G210), .B1(G237), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n256), .A2(new_n257), .A3(new_n191), .ZN(new_n306));
  INV_X1    g120(.A(new_n222), .ZN(new_n307));
  OAI21_X1  g121(.A(G113), .B1(new_n219), .B2(KEYINPUT5), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n248), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n203), .A2(new_n206), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n257), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n191), .B(KEYINPUT86), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT8), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n281), .A2(new_n284), .A3(new_n298), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT7), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT87), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n316), .A2(KEYINPUT87), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n289), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n312), .A2(new_n314), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n306), .B(new_n320), .C1(new_n299), .C2(new_n316), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n303), .A2(new_n305), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n302), .A2(new_n299), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n189), .B1(new_n265), .B2(new_n306), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n258), .A2(new_n190), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n320), .A2(new_n306), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n285), .A2(KEYINPUT84), .B1(new_n283), .B2(new_n297), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n330), .A2(KEYINPUT7), .A3(new_n289), .A4(new_n291), .ZN(new_n331));
  AOI21_X1  g145(.A(G902), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n304), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n188), .B1(new_n324), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n283), .A2(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT16), .ZN(new_n338));
  OR3_X1    g152(.A1(new_n283), .A2(KEYINPUT16), .A3(G140), .ZN(new_n339));
  AOI21_X1  g153(.A(G146), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n338), .A2(G146), .A3(new_n339), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G237), .ZN(new_n344));
  AND4_X1   g158(.A1(G143), .A2(new_n344), .A3(new_n287), .A4(G214), .ZN(new_n345));
  NOR2_X1   g159(.A1(G237), .A2(G953), .ZN(new_n346));
  AOI21_X1  g160(.A(G143), .B1(new_n346), .B2(G214), .ZN(new_n347));
  OAI21_X1  g161(.A(G131), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT17), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n283), .A2(KEYINPUT16), .A3(G140), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(KEYINPUT16), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G146), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT74), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n344), .A2(new_n287), .A3(G214), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n268), .ZN(new_n357));
  INV_X1    g171(.A(G131), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n346), .A2(G143), .A3(G214), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n348), .A2(new_n349), .A3(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n343), .A2(new_n350), .A3(new_n355), .A4(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT88), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n345), .B2(new_n347), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n357), .A2(KEYINPUT88), .A3(new_n359), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT18), .A4(G131), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n336), .A2(new_n337), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT75), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n271), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(G146), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n345), .A2(new_n347), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT18), .A2(G131), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AND4_X1   g191(.A1(new_n374), .A2(new_n357), .A3(new_n376), .A4(new_n359), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n366), .B(new_n373), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(G113), .B(G122), .Z(new_n380));
  XOR2_X1   g194(.A(KEYINPUT90), .B(G104), .Z(new_n381));
  XOR2_X1   g195(.A(new_n380), .B(new_n381), .Z(new_n382));
  NAND3_X1  g196(.A1(new_n362), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n382), .B1(new_n362), .B2(new_n379), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n322), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G475), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT20), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n348), .A2(new_n360), .B1(new_n353), .B2(G146), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT19), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n369), .A2(new_n390), .A3(new_n370), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n367), .A2(KEYINPUT19), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n389), .B1(new_n393), .B2(G146), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n379), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n382), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n383), .ZN(new_n398));
  NOR2_X1   g212(.A1(G475), .A2(G902), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n388), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  AOI211_X1 g215(.A(KEYINPUT20), .B(new_n401), .C1(new_n397), .C2(new_n383), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n387), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n268), .A2(G128), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT13), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT91), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT91), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n407), .A2(new_n268), .A3(KEYINPUT13), .A4(G128), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n295), .A2(G143), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n405), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n406), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G134), .ZN(new_n412));
  XNOR2_X1  g226(.A(G116), .B(G122), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n198), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n211), .A2(G122), .ZN(new_n415));
  INV_X1    g229(.A(G122), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G116), .ZN(new_n417));
  OAI21_X1  g231(.A(G107), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n404), .A2(new_n409), .ZN(new_n419));
  INV_X1    g233(.A(G134), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n414), .A2(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n412), .A2(KEYINPUT92), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n412), .A2(new_n421), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT92), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n404), .A2(new_n409), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G134), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n404), .A2(new_n409), .A3(new_n420), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n427), .A2(new_n428), .B1(new_n198), .B2(new_n413), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n198), .B1(new_n417), .B2(KEYINPUT14), .ZN(new_n430));
  INV_X1    g244(.A(new_n413), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n430), .B1(new_n431), .B2(KEYINPUT14), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT70), .B(G217), .Z(new_n434));
  XOR2_X1   g248(.A(KEYINPUT9), .B(G234), .Z(new_n435));
  AND3_X1   g249(.A1(new_n434), .A2(new_n435), .A3(new_n287), .ZN(new_n436));
  AND4_X1   g250(.A1(new_n422), .A2(new_n425), .A3(new_n433), .A4(new_n436), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n423), .A2(new_n424), .B1(new_n432), .B2(new_n429), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n438), .B2(new_n422), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n322), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G478), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI221_X1 g257(.A(new_n322), .B1(KEYINPUT15), .B2(new_n441), .C1(new_n437), .C2(new_n439), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n287), .A2(G952), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(G234), .B2(G237), .ZN(new_n447));
  AOI211_X1 g261(.A(new_n322), .B(new_n287), .C1(G234), .C2(G237), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(G898), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n403), .A2(new_n445), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G221), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(new_n435), .B2(new_n322), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G140), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n287), .A2(G227), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n455), .B(new_n456), .Z(new_n457));
  OAI211_X1 g271(.A(new_n282), .B(new_n255), .C1(new_n260), .C2(new_n261), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT10), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n297), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n271), .A2(G143), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n296), .A2(new_n461), .A3(new_n273), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n295), .B1(new_n461), .B2(KEYINPUT1), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(new_n279), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n203), .A3(new_n206), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n460), .A2(new_n207), .B1(new_n465), .B2(new_n459), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT11), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n420), .B2(G137), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n420), .A2(G137), .ZN(new_n469));
  INV_X1    g283(.A(G137), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT11), .A3(G134), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G131), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n468), .A2(new_n471), .A3(new_n358), .A4(new_n469), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT80), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n458), .A2(new_n466), .A3(new_n477), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n473), .A2(new_n474), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n458), .B2(new_n466), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n457), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n458), .A2(new_n466), .A3(new_n477), .ZN(new_n482));
  INV_X1    g296(.A(new_n457), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n274), .A2(new_n294), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n462), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n465), .B1(new_n207), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT81), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n487), .B1(new_n479), .B2(new_n488), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n486), .A2(new_n475), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n486), .B2(new_n475), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n482), .B(new_n483), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n481), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G469), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n322), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n322), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n482), .B1(new_n490), .B2(new_n491), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n457), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n458), .A2(new_n466), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n482), .B(new_n483), .C1(new_n500), .C2(new_n479), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(G469), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n495), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n451), .A2(new_n454), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n187), .B1(new_n334), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n188), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n305), .B1(new_n303), .B2(new_n323), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n328), .A2(new_n332), .A3(new_n304), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n502), .A2(new_n497), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n453), .B1(new_n511), .B2(new_n495), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n509), .A2(new_n512), .A3(KEYINPUT93), .A4(new_n451), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n346), .A2(G210), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT27), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(G101), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n470), .A2(G134), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n420), .A2(G137), .ZN(new_n519));
  OAI21_X1  g333(.A(G131), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n474), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n485), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n475), .A2(new_n282), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n263), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(KEYINPUT28), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(KEYINPUT28), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT65), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n475), .A2(new_n528), .A3(new_n282), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n475), .B2(new_n282), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n522), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n251), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n517), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n524), .A2(new_n517), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT68), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT68), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n524), .A2(new_n537), .A3(new_n517), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT30), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n536), .A2(new_n538), .B1(new_n541), .B2(new_n251), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT69), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT31), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n536), .A2(new_n538), .ZN(new_n545));
  INV_X1    g359(.A(new_n539), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n523), .A2(KEYINPUT65), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n475), .A2(new_n528), .A3(new_n282), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n547), .A2(new_n548), .B1(new_n485), .B2(new_n521), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n546), .B(new_n251), .C1(new_n549), .C2(KEYINPUT30), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n545), .A2(new_n543), .A3(KEYINPUT31), .A4(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n534), .B1(new_n544), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(G472), .A2(G902), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(KEYINPUT32), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT32), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n537), .B1(new_n524), .B2(new_n517), .ZN(new_n557));
  INV_X1    g371(.A(new_n538), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n550), .B(new_n543), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT31), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n533), .B1(new_n561), .B2(new_n551), .ZN(new_n562));
  INV_X1    g376(.A(new_n554), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n556), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G472), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n550), .A2(new_n524), .ZN(new_n566));
  INV_X1    g380(.A(new_n517), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT29), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n527), .A2(new_n532), .A3(new_n517), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n263), .B1(new_n522), .B2(new_n523), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n525), .B2(new_n526), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n567), .A2(new_n569), .ZN(new_n574));
  AOI21_X1  g388(.A(G902), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n565), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n555), .A2(new_n564), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT22), .B(G137), .ZN(new_n579));
  INV_X1    g393(.A(G234), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n452), .A2(new_n580), .A3(G953), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n579), .B(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G110), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT72), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n209), .A2(new_n210), .A3(new_n295), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT23), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n217), .A2(G128), .A3(new_n218), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(KEYINPUT72), .A3(KEYINPUT23), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n295), .B1(new_n209), .B2(new_n210), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT73), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(KEYINPUT73), .B(new_n295), .C1(new_n209), .C2(new_n210), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n587), .A2(new_n589), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n295), .A2(KEYINPUT23), .A3(G119), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n583), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n338), .A2(new_n339), .A3(new_n342), .A4(G146), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n353), .B2(G146), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n342), .B1(new_n353), .B2(G146), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n588), .B1(new_n216), .B2(G128), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT24), .B(G110), .ZN(new_n601));
  OAI22_X1  g415(.A1(new_n598), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n354), .A2(new_n371), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT72), .B1(new_n588), .B2(KEYINPUT23), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n583), .B(new_n595), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n600), .A2(new_n601), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n582), .B1(new_n603), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n608), .ZN(new_n611));
  INV_X1    g425(.A(new_n604), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n595), .B1(new_n605), .B2(new_n606), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G110), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n600), .A2(new_n601), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n343), .B2(new_n355), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n582), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n613), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n610), .A2(new_n620), .A3(new_n322), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n621), .A2(KEYINPUT25), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT25), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n610), .A2(new_n620), .A3(new_n623), .A4(new_n322), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n434), .B1(new_n580), .B2(G902), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT71), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT76), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n621), .A2(KEYINPUT25), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT76), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n629), .A2(new_n630), .A3(new_n626), .A4(new_n624), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n610), .A2(new_n620), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n626), .A2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n628), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n505), .A2(new_n513), .A3(new_n578), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT94), .B(G101), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G3));
  NAND2_X1  g453(.A1(new_n561), .A2(new_n551), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n563), .B1(new_n640), .B2(new_n534), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n553), .A2(new_n322), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n641), .B1(new_n642), .B2(G472), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n503), .A2(new_n454), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  AOI211_X1 g459(.A(new_n506), .B(new_n450), .C1(new_n507), .C2(new_n508), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n441), .A2(G902), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT95), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n437), .B2(new_n439), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n649), .B(KEYINPUT33), .C1(new_n437), .C2(new_n439), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n440), .A2(new_n441), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n403), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n643), .A2(new_n645), .A3(new_n646), .A4(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT97), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  INV_X1    g476(.A(new_n445), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n403), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n643), .A2(new_n645), .A3(new_n646), .A4(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  OAI21_X1  g481(.A(G472), .B1(new_n562), .B2(G902), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n553), .A2(new_n554), .ZN(new_n669));
  OAI22_X1  g483(.A1(new_n603), .A2(new_n609), .B1(KEYINPUT36), .B2(new_n582), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n582), .A2(KEYINPUT36), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n613), .A2(new_n618), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n670), .A2(new_n672), .A3(new_n633), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT98), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n628), .A2(new_n631), .A3(new_n674), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n668), .A2(new_n669), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n505), .A2(new_n676), .A3(new_n513), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  NAND2_X1  g493(.A1(new_n507), .A2(new_n508), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n675), .A2(new_n188), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n664), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n447), .B1(new_n448), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n681), .A2(new_n578), .A3(new_n512), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  INV_X1    g501(.A(new_n542), .ZN(new_n688));
  INV_X1    g502(.A(new_n524), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n567), .B1(new_n689), .B2(new_n572), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n691), .B2(G902), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n555), .A2(new_n564), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n403), .A2(new_n445), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n693), .A2(new_n506), .A3(new_n675), .A4(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n684), .B(KEYINPUT39), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n512), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT100), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n680), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n695), .A2(new_n698), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n703), .B(KEYINPUT101), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  INV_X1    g519(.A(new_n684), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n403), .B(new_n706), .C1(new_n654), .C2(new_n655), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n681), .A2(new_n578), .A3(new_n512), .A4(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT102), .B(G146), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G48));
  NOR3_X1   g525(.A1(new_n334), .A2(new_n450), .A3(new_n656), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n494), .B1(new_n493), .B2(new_n322), .ZN(new_n713));
  AOI211_X1 g527(.A(G469), .B(G902), .C1(new_n481), .C2(new_n492), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n714), .A3(new_n453), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n712), .A2(new_n578), .A3(new_n636), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NOR3_X1   g532(.A1(new_n334), .A2(new_n450), .A3(new_n682), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n578), .A3(new_n636), .A4(new_n715), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  AND3_X1   g535(.A1(new_n680), .A2(new_n715), .A3(new_n188), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n578), .A3(new_n451), .A4(new_n675), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  INV_X1    g538(.A(new_n715), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n694), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n573), .A2(new_n517), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n563), .B1(new_n640), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n642), .B2(G472), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n726), .A2(new_n729), .A3(new_n636), .A4(new_n646), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NAND4_X1  g545(.A1(new_n722), .A2(new_n729), .A3(new_n675), .A4(new_n708), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  NAND2_X1  g547(.A1(new_n564), .A2(KEYINPUT103), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n576), .B1(new_n641), .B2(KEYINPUT32), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n736), .B(new_n556), .C1(new_n562), .C2(new_n563), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n507), .A2(new_n188), .A3(new_n508), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n739), .A2(new_n644), .A3(new_n707), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n636), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT42), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n635), .B1(new_n735), .B2(new_n564), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n739), .A2(new_n644), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n742), .A2(KEYINPUT104), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT104), .B1(new_n742), .B2(new_n746), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  AND4_X1   g564(.A1(new_n578), .A2(new_n744), .A3(new_n636), .A4(new_n685), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n420), .ZN(G36));
  INV_X1    g566(.A(new_n739), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n668), .A2(new_n669), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n675), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n654), .A2(new_n655), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n758), .A2(KEYINPUT43), .A3(new_n403), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT43), .B1(new_n758), .B2(new_n403), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n757), .A2(KEYINPUT44), .A3(new_n761), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(KEYINPUT107), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(KEYINPUT107), .ZN(new_n765));
  OAI221_X1 g579(.A(new_n753), .B1(KEYINPUT44), .B2(new_n762), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n499), .A2(new_n501), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n494), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n501), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n496), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OR3_X1    g588(.A1(new_n774), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT105), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n714), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n454), .A3(new_n696), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n768), .A2(new_n769), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n778), .A2(KEYINPUT109), .A3(new_n454), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT109), .B1(new_n778), .B2(new_n454), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n783), .B(new_n784), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n787), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n783), .A2(new_n784), .ZN(new_n790));
  NAND2_X1  g604(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n789), .A2(new_n790), .A3(new_n785), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n578), .A2(new_n636), .A3(new_n707), .A4(new_n739), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  OR2_X1    g610(.A1(G952), .A2(G953), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n738), .A2(new_n636), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n759), .A2(new_n447), .A3(new_n760), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n725), .A2(new_n739), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT48), .Z(new_n802));
  XOR2_X1   g616(.A(new_n446), .B(KEYINPUT120), .Z(new_n803));
  AND2_X1   g617(.A1(new_n729), .A2(new_n636), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n799), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n803), .B1(new_n806), .B2(new_n722), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n693), .A2(new_n636), .A3(new_n447), .A4(new_n800), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n656), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT121), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT121), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n713), .A2(new_n714), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n453), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n788), .A2(new_n792), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n805), .A2(new_n739), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n701), .A2(new_n725), .A3(new_n188), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n806), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT50), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n806), .A2(KEYINPUT50), .A3(new_n818), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n808), .A2(new_n403), .A3(new_n655), .A4(new_n654), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n799), .A2(new_n675), .A3(new_n729), .A4(new_n800), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n811), .A2(new_n812), .B1(new_n817), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n817), .A2(KEYINPUT117), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n815), .A2(new_n835), .A3(new_n816), .ZN(new_n836));
  INV_X1    g650(.A(new_n830), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n838), .A2(KEYINPUT119), .A3(new_n831), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT119), .B1(new_n838), .B2(new_n831), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n833), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(KEYINPUT122), .B(new_n833), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n716), .A2(new_n720), .A3(new_n723), .A4(new_n730), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n742), .A3(new_n746), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n847), .B(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n628), .A2(new_n631), .A3(new_n674), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n454), .B(new_n706), .C1(new_n510), .C2(new_n714), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n852), .A3(KEYINPUT112), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n555), .A2(new_n564), .A3(new_n692), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n675), .B2(new_n851), .ZN(new_n856));
  AOI211_X1 g670(.A(new_n506), .B(new_n694), .C1(new_n507), .C2(new_n508), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n853), .A2(new_n854), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n686), .A2(new_n858), .A3(new_n709), .A4(new_n732), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n644), .B1(new_n735), .B2(new_n564), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n862), .B(new_n681), .C1(new_n685), .C2(new_n708), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(KEYINPUT52), .A3(new_n732), .A4(new_n858), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n403), .A2(new_n445), .A3(new_n684), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n578), .A2(new_n675), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n729), .A2(new_n675), .A3(new_n708), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n751), .B1(new_n869), .B2(new_n744), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n637), .A2(new_n677), .A3(new_n658), .A4(new_n665), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n849), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n865), .A2(KEYINPUT113), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n861), .A2(new_n877), .A3(new_n864), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n846), .A2(new_n871), .A3(new_n870), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n880), .A2(new_n748), .A3(new_n747), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n875), .B(KEYINPUT53), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n880), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n861), .A2(new_n877), .A3(new_n864), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n877), .B1(new_n861), .B2(new_n864), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n749), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT114), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n873), .B(new_n874), .C1(new_n882), .C2(new_n888), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n889), .A2(KEYINPUT116), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n886), .A2(KEYINPUT53), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n881), .A2(new_n887), .A3(new_n865), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(KEYINPUT54), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n889), .A2(KEYINPUT116), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n890), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n797), .B1(new_n845), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n758), .A2(new_n403), .ZN(new_n897));
  INV_X1    g711(.A(new_n813), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n897), .B1(KEYINPUT49), .B2(new_n898), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n899), .B(new_n701), .C1(KEYINPUT49), .C2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n635), .A2(new_n506), .A3(new_n453), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT111), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n693), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n896), .A2(new_n903), .ZN(G75));
  OAI21_X1  g718(.A(new_n873), .B1(new_n882), .B2(new_n888), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(G902), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(G210), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n326), .A2(new_n327), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n325), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT55), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n908), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n908), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n287), .A2(G952), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G51));
  AND4_X1   g732(.A1(G902), .A2(new_n905), .A3(new_n773), .A4(new_n772), .ZN(new_n919));
  INV_X1    g733(.A(new_n493), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n889), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n496), .B(KEYINPUT124), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT57), .Z(new_n924));
  AOI21_X1  g738(.A(new_n920), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n919), .B1(new_n925), .B2(KEYINPUT125), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n927));
  INV_X1    g741(.A(new_n924), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n921), .B2(new_n889), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n929), .B2(new_n920), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n917), .B1(new_n926), .B2(new_n930), .ZN(G54));
  NAND4_X1  g745(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .A4(new_n398), .ZN(new_n932));
  INV_X1    g746(.A(new_n917), .ZN(new_n933));
  NAND2_X1  g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n383), .B(new_n397), .C1(new_n906), .C2(new_n934), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(G60));
  NAND2_X1  g750(.A1(new_n652), .A2(new_n653), .ZN(new_n937));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT59), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n895), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n922), .A2(new_n937), .A3(new_n939), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n917), .A3(new_n941), .ZN(G63));
  AND2_X1   g756(.A1(new_n670), .A2(new_n672), .ZN(new_n943));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n905), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n933), .B1(new_n948), .B2(KEYINPUT61), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n905), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(new_n945), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n947), .B(new_n950), .C1(new_n952), .C2(new_n632), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G66));
  INV_X1    g769(.A(G224), .ZN(new_n956));
  OAI21_X1  g770(.A(G953), .B1(new_n449), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n846), .A2(new_n871), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(G953), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n909), .B1(G898), .B2(new_n287), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G69));
  XNOR2_X1  g775(.A(new_n541), .B(KEYINPUT127), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(new_n393), .Z(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(G900), .B(G953), .C1(new_n964), .C2(G227), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(G227), .B2(new_n964), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n863), .A2(new_n732), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n704), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT62), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n739), .B(new_n697), .C1(new_n656), .C2(new_n682), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n743), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(new_n781), .A3(new_n795), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n963), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n780), .A2(new_n798), .A3(new_n857), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n967), .A2(new_n751), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n749), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n781), .A2(new_n795), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n979), .B2(new_n964), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n966), .B1(new_n974), .B2(new_n980), .ZN(G72));
  NAND2_X1  g795(.A1(new_n566), .A2(new_n517), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n972), .A2(new_n781), .A3(new_n795), .A4(new_n958), .ZN(new_n983));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  AOI21_X1  g799(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n781), .A2(new_n795), .A3(new_n958), .A4(new_n977), .ZN(new_n987));
  AOI211_X1 g801(.A(new_n517), .B(new_n566), .C1(new_n987), .C2(new_n985), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n688), .A2(new_n568), .ZN(new_n989));
  AND4_X1   g803(.A1(new_n891), .A2(new_n892), .A3(new_n985), .A4(new_n989), .ZN(new_n990));
  NOR4_X1   g804(.A1(new_n986), .A2(new_n988), .A3(new_n917), .A4(new_n990), .ZN(G57));
endmodule


