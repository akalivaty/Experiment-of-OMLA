//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT64), .Z(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n209), .B1(new_n211), .B2(new_n214), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  INV_X1    g0047(.A(G68), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n247), .A2(G77), .B1(G20), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n249), .B1(new_n202), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(new_n255), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT11), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT73), .B1(new_n262), .B2(new_n248), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT12), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n262), .A2(new_n255), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n260), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G68), .A3(new_n266), .ZN(new_n267));
  AND4_X1   g0067(.A1(new_n256), .A2(new_n259), .A3(new_n264), .A4(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT67), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G226), .A2(G1698), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n230), .B2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n246), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n274), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G97), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n271), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(new_n271), .A3(G274), .ZN(new_n288));
  INV_X1    g0088(.A(G238), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n271), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT13), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT13), .B1(new_n284), .B2(new_n292), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G179), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT14), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n296), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(KEYINPUT74), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n297), .A2(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(new_n298), .A3(new_n301), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n269), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n296), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n284), .A2(KEYINPUT13), .A3(new_n292), .ZN(new_n307));
  OAI21_X1  g0107(.A(G200), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n295), .A2(G190), .A3(new_n296), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n268), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G58), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT8), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT8), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G58), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n250), .B1(G20), .B2(G77), .ZN(new_n316));
  INV_X1    g0116(.A(G20), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G33), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n255), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT70), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n253), .A2(new_n254), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n261), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n266), .A2(G77), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n265), .A2(KEYINPUT70), .A3(G77), .A4(new_n266), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G77), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n262), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n321), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G244), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n288), .B1(new_n332), .B2(new_n291), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n274), .A2(new_n281), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n289), .A2(G1698), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(G232), .B2(G1698), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT69), .A2(G107), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT69), .A2(G107), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n271), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n333), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G190), .ZN(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n331), .B(new_n344), .C1(new_n345), .C2(new_n343), .ZN(new_n346));
  INV_X1    g0146(.A(G179), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT71), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT71), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n343), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n338), .A2(new_n342), .ZN(new_n353));
  INV_X1    g0153(.A(new_n333), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n320), .A2(new_n255), .B1(new_n329), .B2(new_n262), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n355), .A2(new_n300), .B1(new_n356), .B2(new_n328), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n305), .A2(new_n310), .A3(new_n346), .A4(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT72), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT10), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n360), .A2(KEYINPUT10), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n315), .A2(new_n247), .B1(G150), .B2(new_n250), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n203), .A2(G20), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n323), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n266), .A2(G50), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n324), .A2(new_n366), .B1(G50), .B2(new_n261), .ZN(new_n367));
  OR3_X1    g0167(.A1(new_n365), .A2(new_n367), .A3(KEYINPUT9), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT9), .B1(new_n365), .B2(new_n367), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n334), .A2(G77), .ZN(new_n371));
  XOR2_X1   g0171(.A(KEYINPUT68), .B(G223), .Z(new_n372));
  NAND4_X1  g0172(.A1(new_n372), .A2(new_n274), .A3(new_n281), .A4(G1698), .ZN(new_n373));
  INV_X1    g0173(.A(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G222), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n371), .B(new_n373), .C1(new_n334), .C2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n271), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G226), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n288), .B1(new_n379), .B2(new_n291), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n370), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n380), .B1(new_n376), .B2(new_n377), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(new_n345), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n361), .B(new_n362), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n386), .ZN(new_n388));
  AOI22_X1  g0188(.A1(G190), .A2(new_n385), .B1(new_n368), .B2(new_n369), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n360), .A4(KEYINPUT10), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n382), .A2(G179), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n365), .A2(new_n367), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n385), .B2(G169), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n387), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n315), .A2(new_n266), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n324), .A2(new_n396), .B1(new_n261), .B2(new_n315), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n311), .A2(new_n248), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n398), .A2(new_n201), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(G20), .B1(G159), .B2(new_n250), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  NOR4_X1   g0201(.A1(new_n272), .A2(new_n273), .A3(new_n401), .A4(G20), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT67), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n279), .B1(new_n278), .B2(new_n280), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n317), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n402), .B1(new_n405), .B2(new_n401), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n400), .B1(new_n406), .B2(new_n248), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n272), .A2(new_n273), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT7), .B1(new_n410), .B2(new_n317), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n411), .B2(new_n402), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n400), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n255), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n397), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n271), .A2(G232), .A3(new_n290), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n288), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT75), .ZN(new_n419));
  OR2_X1    g0219(.A1(G223), .A2(G1698), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n379), .A2(G1698), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(new_n272), .C2(new_n273), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G87), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n377), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT75), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n288), .A2(new_n417), .A3(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n419), .A2(new_n425), .A3(new_n427), .A4(new_n347), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n271), .B1(new_n422), .B2(new_n423), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n300), .B1(new_n429), .B2(new_n418), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT76), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n428), .A2(KEYINPUT76), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT18), .B1(new_n416), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n428), .A2(KEYINPUT76), .A3(new_n430), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT76), .B1(new_n428), .B2(new_n430), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n397), .ZN(new_n440));
  INV_X1    g0240(.A(new_n402), .ZN(new_n441));
  AOI21_X1  g0241(.A(G20), .B1(new_n274), .B2(new_n281), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(KEYINPUT7), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G68), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT16), .B1(new_n444), .B2(new_n400), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n440), .B1(new_n445), .B2(new_n414), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n439), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n345), .B1(new_n429), .B2(new_n418), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n419), .A2(new_n427), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n425), .A2(new_n383), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n440), .C1(new_n445), .C2(new_n414), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT17), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n409), .A2(new_n415), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(KEYINPUT17), .A3(new_n440), .A4(new_n452), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n436), .A2(new_n448), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n359), .A2(new_n395), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT23), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n341), .B2(G20), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n317), .A2(G107), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n461), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(new_n318), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT81), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT69), .B(G107), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT23), .B1(new_n468), .B2(new_n317), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT81), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n461), .A2(new_n463), .B1(new_n247), .B2(G116), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n278), .A2(new_n280), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(new_n317), .A3(G87), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT22), .ZN(new_n476));
  OR3_X1    g0276(.A1(new_n216), .A2(KEYINPUT22), .A3(G20), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n334), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT80), .B(KEYINPUT24), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n473), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n473), .B2(new_n478), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n255), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G13), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n463), .ZN(new_n486));
  XNOR2_X1  g0286(.A(new_n486), .B(KEYINPUT25), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n260), .A2(G33), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n261), .A2(new_n488), .A3(new_n254), .A4(new_n253), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(G107), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n260), .A2(G45), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n285), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G264), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n496), .A2(new_n377), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT82), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n374), .A2(G250), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n410), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G294), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n246), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n219), .A2(new_n374), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n474), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n474), .A2(KEYINPUT82), .A3(G250), .A4(new_n374), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n498), .B1(new_n507), .B2(new_n377), .ZN(new_n508));
  INV_X1    g0308(.A(G274), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n210), .B2(new_n270), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n496), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(new_n383), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(G200), .B1(new_n508), .B2(new_n511), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT83), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n511), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n498), .B(new_n516), .C1(new_n507), .C2(new_n377), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n517), .A2(KEYINPUT83), .A3(G200), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n483), .B(new_n491), .C1(new_n515), .C2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(G169), .B1(new_n508), .B2(new_n511), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n347), .B2(new_n517), .ZN(new_n521));
  INV_X1    g0321(.A(new_n472), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n470), .B1(new_n469), .B2(new_n471), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n478), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n479), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n473), .A2(new_n478), .A3(new_n480), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n323), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n491), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n521), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n519), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n519), .B2(new_n529), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT79), .ZN(new_n535));
  OAI21_X1  g0335(.A(G303), .B1(new_n403), .B2(new_n404), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n219), .A2(new_n374), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n497), .A2(G1698), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n538), .C1(new_n272), .C2(new_n273), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n271), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n286), .A2(G1), .ZN(new_n541));
  INV_X1    g0341(.A(new_n495), .ZN(new_n542));
  NOR2_X1   g0342(.A1(KEYINPUT5), .A2(G41), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n271), .ZN(new_n545));
  INV_X1    g0345(.A(G270), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n511), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n535), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G303), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n274), .B2(new_n281), .ZN(new_n550));
  INV_X1    g0350(.A(new_n539), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n377), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n494), .A2(new_n495), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(new_n541), .B1(new_n210), .B2(new_n270), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(G270), .B1(new_n510), .B2(new_n496), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n555), .A3(KEYINPUT79), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G283), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n557), .B(new_n317), .C1(G33), .C2(new_n218), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n465), .A2(G20), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n255), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT20), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n558), .A2(KEYINPUT20), .A3(new_n255), .A4(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n261), .A2(G116), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n490), .B2(G116), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n300), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n548), .A2(KEYINPUT21), .A3(new_n556), .A4(new_n567), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n540), .A2(new_n547), .A3(new_n347), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n548), .A2(new_n556), .A3(new_n567), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n552), .A2(new_n555), .A3(KEYINPUT79), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT79), .B1(new_n552), .B2(new_n555), .ZN(new_n577));
  OAI21_X1  g0377(.A(G190), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n570), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n548), .A2(G200), .A3(new_n556), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n572), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n319), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n261), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n489), .A2(new_n319), .ZN(new_n585));
  NAND3_X1  g0385(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n317), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G87), .A2(G97), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n587), .B1(new_n468), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n317), .B(G68), .C1(new_n272), .C2(new_n273), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n318), .B2(new_n218), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AOI211_X1 g0394(.A(new_n584), .B(new_n585), .C1(new_n594), .C2(new_n255), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n289), .A2(new_n374), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n332), .A2(G1698), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(new_n272), .C2(new_n273), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n246), .A2(new_n465), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n271), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n271), .A2(G274), .A3(new_n541), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n217), .B1(new_n260), .B2(G45), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n271), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n300), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n510), .A2(new_n541), .B1(new_n271), .B2(new_n603), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G238), .A2(G1698), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n332), .B2(G1698), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n599), .B1(new_n609), .B2(new_n474), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n607), .B(new_n347), .C1(new_n610), .C2(new_n271), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n601), .B2(new_n605), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n607), .B(G190), .C1(new_n610), .C2(new_n271), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n341), .A2(new_n588), .B1(new_n317), .B2(new_n586), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n591), .A2(new_n593), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n255), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n584), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n490), .A2(G87), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n595), .A2(new_n612), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT78), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n618), .A2(new_n619), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n606), .B(new_n611), .C1(new_n624), .C2(new_n585), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n584), .B1(new_n594), .B2(new_n255), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(new_n620), .A3(new_n613), .A4(new_n614), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT78), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n544), .A2(G257), .A3(new_n271), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n511), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n274), .A2(new_n281), .A3(G250), .A4(G1698), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT4), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n634), .A2(new_n332), .A3(G1698), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n274), .A2(new_n281), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n374), .A2(G244), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n410), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n633), .A2(new_n636), .A3(new_n557), .A4(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n632), .B1(new_n639), .B2(new_n377), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n300), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n261), .A2(G97), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n490), .B2(G97), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT6), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n645), .A2(new_n218), .A3(G107), .ZN(new_n646));
  XNOR2_X1  g0446(.A(G97), .B(G107), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  OAI22_X1  g0448(.A1(new_n648), .A2(new_n317), .B1(new_n329), .B2(new_n251), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n443), .B2(new_n468), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n644), .B1(new_n650), .B2(new_n323), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT77), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n640), .A2(new_n652), .A3(new_n347), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(new_n640), .B2(new_n347), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n642), .B(new_n651), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n650), .A2(new_n323), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n641), .A2(G200), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n640), .A2(G190), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n644), .A4(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n630), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  NOR4_X1   g0460(.A1(new_n460), .A2(new_n534), .A3(new_n582), .A4(new_n660), .ZN(G372));
  INV_X1    g0461(.A(new_n394), .ZN(new_n662));
  INV_X1    g0462(.A(new_n305), .ZN(new_n663));
  INV_X1    g0463(.A(new_n358), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n310), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT85), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n457), .A2(new_n455), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n439), .A2(new_n446), .A3(new_n447), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n447), .B1(new_n439), .B2(new_n446), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n387), .A2(new_n390), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n662), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n529), .A2(new_n575), .A3(new_n572), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n527), .A2(new_n528), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n513), .A2(new_n514), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT83), .B1(new_n517), .B2(G200), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(new_n512), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n622), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n655), .A2(new_n659), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n677), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n622), .A2(KEYINPUT78), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n628), .B1(new_n625), .B2(new_n627), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT26), .B1(new_n687), .B2(new_n655), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n653), .A2(new_n654), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n642), .A2(new_n651), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT26), .ZN(new_n691));
  INV_X1    g0491(.A(new_n622), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n688), .A2(new_n625), .A3(new_n693), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n684), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n459), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n676), .A2(new_n696), .ZN(G369));
  NAND2_X1  g0497(.A1(new_n485), .A2(new_n317), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT86), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(G343), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(G343), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n529), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n705), .B1(new_n527), .B2(new_n528), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n707), .B1(new_n533), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n572), .A2(new_n575), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n706), .A2(new_n579), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n582), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n529), .A2(new_n705), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n705), .B1(new_n572), .B2(new_n575), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n717), .B1(new_n533), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n207), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n468), .A2(G116), .A3(new_n589), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(G1), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n214), .B2(new_n723), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n695), .A2(new_n706), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT87), .B1(new_n728), .B2(KEYINPUT29), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n630), .A2(new_n689), .A3(new_n691), .A4(new_n690), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT26), .B1(new_n655), .B2(new_n622), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n625), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT88), .ZN(new_n733));
  AND4_X1   g0533(.A1(new_n519), .A2(new_n655), .A3(new_n659), .A4(new_n692), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n732), .A2(new_n733), .B1(new_n734), .B2(new_n677), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n730), .A2(new_n731), .A3(KEYINPUT88), .A4(new_n625), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n705), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n695), .A2(new_n706), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT87), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT29), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n729), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n572), .A2(new_n581), .A3(new_n575), .A4(new_n706), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n660), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n531), .B2(new_n532), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n540), .A2(new_n547), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n601), .A2(new_n605), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(G179), .A3(new_n508), .A4(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n747), .B1(new_n750), .B2(new_n641), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n508), .A2(new_n749), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n752), .A2(KEYINPUT30), .A3(new_n569), .A4(new_n640), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n347), .B1(new_n601), .B2(new_n605), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n508), .B2(new_n511), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n755), .A2(new_n641), .A3(new_n548), .A4(new_n556), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n751), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT31), .B1(new_n757), .B2(new_n705), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n746), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G330), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n743), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n727), .B1(new_n763), .B2(G1), .ZN(G364));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n254), .B1(G20), .B2(new_n300), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n721), .A2(new_n474), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n213), .B2(new_n286), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(KEYINPUT90), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n772), .A2(KEYINPUT90), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n773), .B(new_n774), .C1(G45), .C2(new_n244), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n335), .A2(G355), .A3(new_n207), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G116), .B2(new_n207), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n769), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n317), .A2(new_n347), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G190), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G200), .ZN(new_n781));
  NOR4_X1   g0581(.A1(new_n317), .A2(new_n345), .A3(G179), .A4(G190), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n781), .A2(G322), .B1(G283), .B2(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n383), .A2(G179), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n317), .ZN(new_n785));
  INV_X1    g0585(.A(G326), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n780), .A2(new_n345), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n783), .B1(new_n502), .B2(new_n785), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n779), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n790), .A2(new_n345), .A3(G190), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT33), .B(G317), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(G311), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n317), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT91), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT91), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G329), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n334), .B(new_n794), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NOR4_X1   g0601(.A1(new_n317), .A2(new_n383), .A3(new_n345), .A4(G179), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT92), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(KEYINPUT92), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n789), .B(new_n801), .C1(G303), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  OAI21_X1  g0609(.A(KEYINPUT32), .B1(new_n799), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n216), .B2(new_n806), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G68), .A2(new_n791), .B1(new_n793), .B2(G77), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n785), .A2(new_n218), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G58), .B2(new_n781), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n787), .A2(G50), .B1(G107), .B2(new_n782), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n812), .A2(new_n814), .A3(new_n335), .A4(new_n815), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n799), .A2(KEYINPUT32), .A3(new_n809), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n811), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n768), .B1(new_n808), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n484), .A2(G20), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G45), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G1), .ZN(new_n822));
  OR3_X1    g0622(.A1(new_n722), .A2(new_n822), .A3(KEYINPUT89), .ZN(new_n823));
  OAI21_X1  g0623(.A(KEYINPUT89), .B1(new_n722), .B2(new_n822), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n778), .A2(new_n819), .A3(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT93), .Z(new_n828));
  INV_X1    g0628(.A(new_n767), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n713), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n713), .A2(G330), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n714), .A2(new_n825), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT94), .Z(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G396));
  INV_X1    g0635(.A(KEYINPUT96), .ZN(new_n836));
  INV_X1    g0636(.A(new_n351), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n350), .B1(new_n343), .B2(new_n347), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n357), .B(new_n706), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n356), .A2(new_n328), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n705), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n346), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n836), .B(new_n839), .C1(new_n664), .C2(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n352), .A2(new_n357), .B1(new_n346), .B2(new_n841), .ZN(new_n844));
  INV_X1    g0644(.A(new_n839), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT96), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n706), .B(new_n847), .C1(new_n684), .C2(new_n694), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n847), .B(KEYINPUT97), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n848), .B1(new_n850), .B2(new_n728), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n826), .B1(new_n851), .B2(new_n762), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n762), .B2(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(new_n791), .ZN(new_n854));
  INV_X1    g0654(.A(G283), .ZN(new_n855));
  INV_X1    g0655(.A(new_n793), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n854), .A2(new_n855), .B1(new_n856), .B2(new_n465), .ZN(new_n857));
  INV_X1    g0657(.A(new_n799), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n335), .B(new_n857), .C1(new_n858), .C2(G311), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n807), .A2(G107), .ZN(new_n860));
  INV_X1    g0660(.A(new_n782), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n788), .A2(new_n549), .B1(new_n216), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n813), .B(new_n862), .C1(G294), .C2(new_n781), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G150), .A2(new_n791), .B1(new_n793), .B2(G159), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n781), .A2(G143), .ZN(new_n866));
  INV_X1    g0666(.A(G137), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n865), .B(new_n866), .C1(new_n867), .C2(new_n788), .ZN(new_n868));
  XNOR2_X1  g0668(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n868), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n474), .B1(new_n861), .B2(new_n248), .ZN(new_n871));
  INV_X1    g0671(.A(new_n785), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(G58), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(G132), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n873), .B1(new_n799), .B2(new_n874), .C1(new_n806), .C2(new_n202), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n864), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n768), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n768), .A2(new_n765), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n825), .B1(new_n329), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n877), .B(new_n879), .C1(new_n847), .C2(new_n766), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n853), .A2(new_n880), .ZN(G384));
  INV_X1    g0681(.A(new_n648), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n465), .B(new_n211), .C1(new_n882), .C2(KEYINPUT35), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(KEYINPUT35), .B2(new_n882), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT36), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n214), .A2(new_n329), .A3(new_n398), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n202), .B2(G68), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n484), .A2(G1), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT98), .Z(new_n890));
  NAND4_X1  g0690(.A1(new_n729), .A2(new_n738), .A3(new_n459), .A4(new_n742), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n891), .A2(new_n676), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n663), .A2(new_n706), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT100), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT16), .B1(new_n412), .B2(new_n400), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n440), .B1(new_n414), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n701), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n458), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n897), .A2(new_n433), .A3(new_n434), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n453), .A3(new_n899), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n439), .A2(new_n446), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n446), .A2(new_n898), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .A4(new_n453), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n901), .A2(KEYINPUT38), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n901), .B2(new_n909), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n895), .B(KEYINPUT39), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n901), .A2(KEYINPUT38), .A3(new_n909), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n905), .A2(new_n906), .A3(new_n453), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n916));
  INV_X1    g0716(.A(new_n906), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n908), .A2(new_n916), .B1(new_n458), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n913), .B(new_n914), .C1(new_n918), .C2(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT38), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n899), .B1(new_n673), .B2(new_n668), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n904), .A2(new_n908), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n913), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n895), .B1(new_n925), .B2(KEYINPUT39), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n894), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n673), .A2(new_n898), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n297), .A2(new_n298), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n299), .A2(new_n301), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n303), .B(new_n310), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n268), .A2(new_n706), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT99), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n305), .B(new_n310), .C1(new_n268), .C2(new_n706), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT99), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n931), .A2(new_n936), .A3(new_n932), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n839), .B2(new_n848), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n928), .B1(new_n940), .B2(new_n925), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n927), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n892), .B(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n761), .A2(new_n938), .A3(new_n847), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n910), .A2(new_n911), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n847), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n746), .B2(new_n760), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n913), .B1(new_n918), .B2(KEYINPUT38), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n949), .A2(new_n950), .A3(KEYINPUT40), .A4(new_n938), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n947), .A2(new_n459), .A3(new_n951), .A4(new_n761), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(G330), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n947), .A2(new_n951), .B1(new_n459), .B2(new_n761), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n943), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n260), .B2(new_n820), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n943), .A2(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n890), .B1(new_n957), .B2(new_n958), .ZN(G367));
  NOR2_X1   g0759(.A1(new_n785), .A2(new_n248), .ZN(new_n960));
  INV_X1    g0760(.A(new_n781), .ZN(new_n961));
  INV_X1    g0761(.A(G150), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n961), .A2(new_n962), .B1(new_n329), .B2(new_n861), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n960), .B(new_n963), .C1(G143), .C2(new_n787), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n807), .A2(G58), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n858), .A2(G137), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n854), .A2(new_n809), .B1(new_n856), .B2(new_n202), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n334), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT106), .B1(new_n807), .B2(G116), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT46), .Z(new_n971));
  OAI22_X1  g0771(.A1(new_n861), .A2(new_n218), .B1(new_n785), .B2(new_n341), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n410), .B1(new_n854), .B2(new_n502), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(G283), .C2(new_n793), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n781), .A2(G303), .B1(new_n787), .B2(G311), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT105), .Z(new_n976));
  INV_X1    g0776(.A(G317), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n974), .B(new_n976), .C1(new_n977), .C2(new_n799), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n969), .B1(new_n971), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT47), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n768), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n236), .A2(new_n770), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n768), .B(new_n767), .C1(new_n721), .C2(new_n583), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n825), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n705), .A2(new_n621), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n625), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT101), .ZN(new_n987));
  INV_X1    g0787(.A(new_n985), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n986), .B(new_n987), .C1(new_n622), .C2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n987), .B2(new_n986), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n981), .B(new_n984), .C1(new_n991), .C2(new_n829), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n822), .B(KEYINPUT104), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n651), .A2(new_n705), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n683), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n655), .B2(new_n706), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n719), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT45), .Z(new_n999));
  NOR2_X1   g0799(.A1(new_n719), .A2(new_n997), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT44), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n716), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(new_n716), .A3(new_n1001), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n718), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n709), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT103), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n533), .B2(new_n718), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n534), .A2(new_n1005), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n1007), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n714), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n714), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1003), .A2(new_n763), .A3(new_n1004), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n763), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n722), .B(KEYINPUT41), .Z(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n994), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1010), .A2(new_n997), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n659), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n655), .B1(new_n1022), .B2(new_n529), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1021), .A2(KEYINPUT42), .B1(new_n706), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(KEYINPUT42), .B2(new_n1021), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1025), .A2(new_n1028), .A3(new_n1026), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n715), .A2(new_n997), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(KEYINPUT102), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1033), .B(KEYINPUT102), .Z(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n992), .B1(new_n1020), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT107), .Z(G387));
  NOR2_X1   g0838(.A1(new_n763), .A2(new_n1015), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n714), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1042), .A2(new_n743), .A3(new_n762), .A4(new_n1012), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n722), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n1012), .A3(new_n994), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT108), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n709), .A2(new_n767), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n724), .ZN(new_n1049));
  AOI211_X1 g0849(.A(G45), .B(new_n1049), .C1(G68), .C2(G77), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(KEYINPUT109), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n315), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n1052), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1053));
  OAI21_X1  g0853(.A(KEYINPUT50), .B1(new_n1052), .B2(G50), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1050), .A2(KEYINPUT109), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n770), .B1(new_n286), .B2(new_n233), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1049), .A2(new_n335), .A3(new_n207), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(G107), .C2(new_n207), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n825), .B1(new_n1059), .B2(new_n769), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n785), .A2(new_n319), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n961), .A2(new_n202), .B1(new_n788), .B2(new_n809), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(G97), .C2(new_n782), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n474), .B1(new_n856), .B2(new_n248), .C1(new_n1052), .C2(new_n854), .ZN(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT110), .B(G150), .Z(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n858), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n807), .A2(G77), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n1063), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n807), .A2(G294), .B1(G283), .B2(new_n872), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G303), .A2(new_n793), .B1(new_n791), .B2(G311), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n787), .A2(G322), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n977), .C2(new_n961), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1069), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT111), .Z(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1070), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT49), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n410), .B1(new_n465), .B2(new_n861), .C1(new_n799), .C2(new_n786), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n1078), .B2(KEYINPUT49), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1068), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n768), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1048), .B(new_n1060), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1045), .A2(new_n1047), .A3(new_n1084), .ZN(G393));
  INV_X1    g0885(.A(new_n1004), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1043), .B1(new_n1086), .B2(new_n1002), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1016), .A2(new_n1087), .A3(new_n722), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n241), .A2(new_n771), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n769), .B1(new_n218), .B2(new_n207), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n826), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n861), .A2(new_n216), .B1(new_n785), .B2(new_n329), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n474), .B1(new_n856), .B2(new_n1052), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(G50), .C2(new_n791), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n781), .A2(G159), .B1(new_n787), .B2(G150), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT51), .Z(new_n1096));
  NAND2_X1  g0896(.A1(new_n807), .A2(G68), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n858), .A2(G143), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n781), .A2(G311), .B1(new_n787), .B2(G317), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1101));
  XNOR2_X1  g0901(.A(new_n1100), .B(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n807), .A2(G283), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n858), .A2(G322), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n854), .A2(new_n549), .B1(new_n856), .B2(new_n502), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n335), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n872), .A2(G116), .B1(G107), .B2(new_n782), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1099), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1091), .B1(new_n1109), .B2(new_n768), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n997), .B2(new_n829), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1088), .B(new_n1111), .C1(new_n1112), .C2(new_n993), .ZN(G390));
  NAND2_X1  g0913(.A1(new_n949), .A2(G330), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n939), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n949), .A2(G330), .A3(new_n938), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1115), .A2(new_n1116), .B1(new_n839), .B2(new_n848), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n939), .B1(new_n849), .B2(new_n762), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n845), .B1(new_n737), .B2(new_n847), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1118), .A2(new_n1119), .A3(new_n1116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT113), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT113), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1118), .A2(new_n1119), .A3(new_n1122), .A4(new_n1116), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1117), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n761), .A2(new_n459), .A3(G330), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n891), .A2(new_n676), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1116), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n848), .A2(new_n839), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n894), .B1(new_n1130), .B2(new_n938), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1131), .A2(new_n920), .A3(new_n926), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n950), .A2(new_n893), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n732), .A2(new_n733), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n734), .A2(new_n677), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n736), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n706), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n839), .B1(new_n1137), .B2(new_n948), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1133), .B1(new_n1138), .B2(new_n938), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1129), .B1(new_n1132), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n893), .B(new_n950), .C1(new_n1119), .C2(new_n939), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT100), .B1(new_n946), .B2(new_n914), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n919), .A3(new_n912), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1141), .B(new_n1116), .C1(new_n1143), .C2(new_n1131), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n723), .B1(new_n1128), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1145), .B2(new_n1128), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1140), .A2(new_n1144), .A3(new_n994), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n807), .A2(new_n1065), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT53), .Z(new_n1150));
  AOI22_X1  g0950(.A1(new_n872), .A2(G159), .B1(G50), .B2(new_n782), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n781), .A2(G132), .B1(new_n787), .B2(G128), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n335), .B1(new_n854), .B2(new_n867), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT114), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(new_n856), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1153), .B(new_n1157), .C1(G125), .C2(new_n858), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1158), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n799), .A2(new_n502), .B1(new_n248), .B2(new_n861), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT116), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n468), .A2(new_n791), .B1(new_n793), .B2(G97), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n855), .B2(new_n788), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT115), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n334), .B1(new_n329), .B2(new_n785), .C1(new_n961), .C2(new_n465), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n807), .B2(G87), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1161), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1083), .B1(new_n1159), .B2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n825), .B(new_n1168), .C1(new_n1052), .C2(new_n878), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n1143), .B2(new_n766), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1147), .A2(new_n1148), .A3(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(KEYINPUT120), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n761), .A2(new_n847), .A3(new_n938), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT40), .B1(new_n1173), .B2(new_n925), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n916), .A2(new_n908), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n458), .A2(new_n917), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT38), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT40), .B1(new_n910), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(G330), .B1(new_n1178), .B2(new_n945), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1172), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n392), .A2(new_n898), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n395), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n387), .A2(new_n390), .A3(new_n394), .A4(new_n1181), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1183), .A2(new_n1186), .A3(new_n1184), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n947), .A2(KEYINPUT120), .A3(new_n951), .A4(G330), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1180), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT118), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1183), .A2(new_n1186), .A3(new_n1184), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1186), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1188), .A2(KEYINPUT118), .A3(new_n1189), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n947), .A2(G330), .A3(new_n951), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1192), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n942), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1199), .A2(new_n927), .A3(new_n941), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT121), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1203), .A2(new_n1204), .A3(new_n1192), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n1203), .B2(new_n1192), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1202), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT122), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(KEYINPUT122), .B(new_n1202), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1127), .B1(new_n1145), .B2(new_n1124), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT123), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT123), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1214), .B(new_n1127), .C1(new_n1145), .C2(new_n1124), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT57), .B1(new_n1211), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT57), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1203), .A2(new_n1192), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1202), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1216), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n722), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1217), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1196), .A2(new_n1197), .A3(new_n765), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n878), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n826), .B1(G50), .B2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n474), .A2(G41), .ZN(new_n1227));
  AOI211_X1 g1027(.A(G50), .B(new_n1227), .C1(new_n246), .C2(new_n285), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1227), .B1(new_n856), .B2(new_n319), .C1(new_n218), .C2(new_n854), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G283), .B2(new_n858), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n861), .A2(new_n311), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n960), .B(new_n1231), .C1(G116), .C2(new_n787), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n781), .A2(G107), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT117), .Z(new_n1234));
  NAND4_X1  g1034(.A1(new_n1230), .A2(new_n1232), .A3(new_n1067), .A4(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT58), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1228), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n854), .A2(new_n874), .B1(new_n856), .B2(new_n867), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G125), .B2(new_n787), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n872), .A2(G150), .B1(new_n781), .B2(G128), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n806), .C2(new_n1156), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n858), .A2(G124), .ZN(new_n1243));
  AOI211_X1 g1043(.A(G33), .B(G41), .C1(new_n782), .C2(G159), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1237), .B1(new_n1236), .B2(new_n1235), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1226), .B1(new_n1247), .B2(new_n768), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1224), .A2(new_n1248), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT119), .Z(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1211), .B2(new_n994), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1223), .A2(new_n1251), .ZN(G375));
  INV_X1    g1052(.A(new_n1127), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1124), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n1128), .A3(new_n1019), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT124), .Z(new_n1256));
  OAI21_X1  g1056(.A(new_n826), .B1(G68), .B2(new_n1225), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n961), .A2(new_n855), .B1(new_n788), .B2(new_n502), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1061), .B(new_n1258), .C1(G77), .C2(new_n782), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n807), .A2(G97), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n858), .A2(G303), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n854), .A2(new_n465), .B1(new_n856), .B2(new_n341), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(new_n335), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .A4(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n474), .B1(new_n856), .B2(new_n962), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1231), .B(new_n1265), .C1(new_n791), .C2(new_n1155), .ZN(new_n1266));
  INV_X1    g1066(.A(G128), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n799), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n872), .A2(G50), .B1(new_n781), .B2(G137), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n1269), .B1(new_n874), .B2(new_n788), .C1(new_n806), .C2(new_n809), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1264), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1257), .B1(new_n1271), .B2(new_n768), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n938), .B2(new_n766), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1256), .B(new_n1273), .C1(new_n993), .C2(new_n1124), .ZN(G381));
  NAND4_X1  g1074(.A1(new_n1045), .A2(new_n1047), .A3(new_n834), .A4(new_n1084), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G384), .A2(G378), .A3(G390), .A4(new_n1275), .ZN(new_n1276));
  OR4_X1    g1076(.A1(G387), .A2(G375), .A3(new_n1276), .A4(G381), .ZN(G407));
  INV_X1    g1077(.A(G378), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n703), .A2(new_n704), .A3(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G407), .B(G213), .C1(G375), .C2(new_n1281), .ZN(G409));
  XOR2_X1   g1082(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1283));
  OAI211_X1 g1083(.A(G378), .B(new_n1251), .C1(new_n1217), .C2(new_n1222), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1219), .A2(KEYINPUT121), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1203), .A2(new_n1192), .A3(new_n1204), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT122), .B1(new_n1287), .B2(new_n1202), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1210), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1019), .B(new_n1216), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n993), .B1(new_n1202), .B2(new_n1219), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1224), .B2(new_n1248), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1278), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1284), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1279), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  OAI221_X1 g1097(.A(new_n1273), .B1(new_n1124), .B2(new_n993), .C1(G384), .C2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1128), .A2(KEYINPUT60), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1254), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1253), .A2(KEYINPUT60), .A3(new_n1124), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1301), .A2(new_n722), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1298), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT125), .B1(new_n853), .B2(new_n880), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1283), .B1(new_n1296), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1280), .A2(G2897), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1310), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1047), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1084), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1319));
  OAI21_X1  g1119(.A(G396), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1275), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(G390), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT107), .B1(new_n1320), .B2(new_n1275), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1322), .B1(G390), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1037), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1322), .B(new_n1037), .C1(G390), .C2(new_n1323), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1280), .B1(new_n1284), .B2(new_n1294), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1308), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(KEYINPUT63), .A3(new_n1330), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1309), .A2(new_n1317), .A3(new_n1328), .A4(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1329), .A2(new_n1333), .A3(new_n1330), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT61), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1335), .B1(new_n1329), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1333), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1334), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1326), .A2(KEYINPUT127), .A3(new_n1327), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT127), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1332), .B1(new_n1339), .B2(new_n1342), .ZN(G405));
  AOI21_X1  g1143(.A(G378), .B1(new_n1223), .B2(new_n1251), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1284), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1308), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(G375), .A2(new_n1278), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(new_n1284), .A3(new_n1330), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1342), .A2(new_n1346), .A3(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1342), .B1(new_n1348), .B2(new_n1346), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1349), .A2(new_n1350), .ZN(G402));
endmodule


