//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G71gat), .ZN(new_n204));
  INV_X1    g003(.A(G99gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G227gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(G183gat), .A3(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT24), .ZN(new_n211));
  NOR2_X1   g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(G169gat), .A3(G176gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n215), .A2(new_n217), .B1(KEYINPUT23), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n213), .B1(new_n219), .B2(KEYINPUT66), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n215), .A2(new_n217), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n220), .A2(new_n225), .A3(KEYINPUT25), .A4(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n228));
  INV_X1    g027(.A(new_n212), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT24), .A3(new_n210), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n230), .A2(new_n226), .A3(new_n214), .A4(new_n209), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n228), .B1(new_n231), .B2(new_n224), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT26), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n214), .B1(new_n218), .B2(new_n234), .ZN(new_n235));
  NOR3_X1   g034(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n210), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g038(.A(KEYINPUT67), .B(new_n210), .C1(new_n235), .C2(new_n236), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT27), .B(G183gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT28), .ZN(new_n243));
  INV_X1    g042(.A(G190gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n243), .B1(new_n242), .B2(new_n244), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G113gat), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G120gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G127gat), .B(G134gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT1), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n253), .A2(G120gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n251), .A2(G113gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT69), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265));
  INV_X1    g064(.A(G127gat), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n266), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n256), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n264), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n265), .B1(new_n264), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n258), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n250), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n227), .A2(new_n232), .B1(new_n241), .B2(new_n248), .ZN(new_n274));
  INV_X1    g073(.A(new_n258), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n264), .A2(new_n269), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT70), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n264), .A2(new_n265), .A3(new_n269), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n207), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(KEYINPUT71), .B(new_n206), .C1(new_n281), .C2(KEYINPUT33), .ZN(new_n282));
  INV_X1    g081(.A(new_n207), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n250), .A2(new_n272), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n274), .A2(new_n279), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT32), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT33), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n274), .B(new_n272), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(new_n207), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT32), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n280), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(new_n283), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n291), .A2(new_n294), .A3(KEYINPUT71), .A4(new_n206), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n207), .A3(new_n280), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT34), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n288), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n297), .B1(new_n288), .B2(new_n295), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT89), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n297), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(new_n286), .B2(new_n289), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n294), .B1(new_n303), .B2(new_n206), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n282), .A2(new_n287), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT89), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n295), .A3(new_n297), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT85), .B(G22gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(G78gat), .B(G106gat), .ZN(new_n312));
  INV_X1    g111(.A(G50gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT22), .ZN(new_n319));
  NAND2_X1  g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320));
  INV_X1    g119(.A(G211gat), .ZN(new_n321));
  INV_X1    g120(.A(G218gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT22), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n320), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n326), .A2(new_n327), .A3(new_n318), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n326), .B2(new_n318), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n318), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT73), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n326), .A2(new_n327), .A3(new_n318), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(KEYINPUT74), .A3(new_n324), .ZN(new_n337));
  AND2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n339));
  NOR2_X1   g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G141gat), .B(G148gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n338), .A2(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n339), .A2(KEYINPUT77), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT2), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n344), .B1(new_n348), .B2(new_n342), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(KEYINPUT78), .B(new_n344), .C1(new_n348), .C2(new_n342), .ZN(new_n352));
  AOI211_X1 g151(.A(KEYINPUT3), .B(new_n343), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n332), .B(new_n337), .C1(new_n353), .C2(KEYINPUT29), .ZN(new_n354));
  INV_X1    g153(.A(G228gat), .ZN(new_n355));
  INV_X1    g154(.A(G233gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n343), .B1(new_n351), .B2(new_n352), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT3), .B1(new_n330), .B2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n354), .B(new_n357), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n360), .B2(new_n358), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n351), .A2(new_n352), .ZN(new_n364));
  INV_X1    g163(.A(new_n343), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n336), .B2(new_n324), .ZN(new_n367));
  OAI211_X1 g166(.A(KEYINPUT82), .B(new_n366), .C1(new_n367), .C2(KEYINPUT3), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n354), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n370));
  INV_X1    g169(.A(new_n357), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n370), .B1(new_n369), .B2(new_n371), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n361), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(KEYINPUT84), .B(new_n361), .C1(new_n372), .C2(new_n373), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n317), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n317), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n311), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n369), .A2(new_n371), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT83), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT84), .B1(new_n385), .B2(new_n361), .ZN(new_n386));
  INV_X1    g185(.A(new_n377), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n316), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n311), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n379), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n332), .A2(new_n337), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n250), .A2(new_n359), .B1(G226gat), .B2(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(G226gat), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n274), .A2(new_n394), .A3(new_n356), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n392), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n250), .A2(G226gat), .A3(G233gat), .ZN(new_n397));
  OAI22_X1  g196(.A1(new_n274), .A2(KEYINPUT29), .B1(new_n394), .B2(new_n356), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n391), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT30), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT76), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n396), .A2(KEYINPUT30), .A3(new_n399), .A4(new_n403), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT75), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n397), .A2(new_n398), .A3(new_n391), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n396), .A2(KEYINPUT75), .A3(new_n399), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n403), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n408), .A2(new_n407), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n409), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n310), .A2(new_n381), .A3(new_n390), .A4(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G1gat), .B(G29gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(G85gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT0), .B(G57gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n353), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n366), .A2(KEYINPUT3), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n272), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n358), .B(new_n258), .C1(new_n270), .C2(new_n271), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n427), .A2(KEYINPUT4), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(KEYINPUT4), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n423), .B(new_n426), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n431));
  NAND2_X1  g230(.A1(new_n272), .A2(new_n366), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n427), .ZN(new_n433));
  INV_X1    g232(.A(new_n423), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n427), .B(KEYINPUT4), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n437), .A2(new_n423), .A3(new_n426), .A4(new_n431), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n422), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n422), .A3(new_n438), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n436), .A2(new_n422), .A3(new_n438), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(new_n439), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(KEYINPUT86), .A3(new_n442), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n446), .A2(new_n449), .B1(new_n439), .B2(new_n441), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n202), .B1(new_n418), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n390), .A2(new_n381), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n439), .A2(new_n441), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n444), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n417), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(new_n202), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT72), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n288), .A2(new_n295), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n297), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n301), .A2(new_n288), .A3(new_n295), .A4(new_n458), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n453), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n451), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n411), .A2(new_n412), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT37), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n403), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n396), .A2(new_n470), .A3(new_n399), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n411), .A2(KEYINPUT87), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT37), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n468), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n474), .A2(new_n404), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT86), .B1(new_n448), .B2(new_n442), .ZN(new_n476));
  NOR4_X1   g275(.A1(new_n447), .A2(new_n439), .A3(new_n445), .A4(new_n441), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n475), .B(new_n454), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n468), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n467), .B1(new_n413), .B2(new_n414), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT38), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n446), .A2(new_n449), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n484), .A2(KEYINPUT88), .A3(new_n454), .A4(new_n475), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n437), .A2(KEYINPUT39), .A3(new_n426), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT39), .B1(new_n437), .B2(new_n426), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n434), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n433), .A2(KEYINPUT39), .A3(new_n423), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n422), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n493), .A2(new_n417), .A3(new_n439), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n452), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n486), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n452), .A2(new_n456), .ZN(new_n498));
  OR3_X1    g297(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT36), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n460), .A2(KEYINPUT36), .A3(new_n461), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n465), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G71gat), .B(G78gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT94), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507));
  INV_X1    g306(.A(G71gat), .ZN(new_n508));
  INV_X1    g307(.A(G78gat), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G64gat), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n511), .A2(G57gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(G57gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT95), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT96), .B(G57gat), .Z(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(new_n511), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n510), .B(new_n504), .C1(new_n519), .C2(new_n512), .ZN(new_n520));
  NAND2_X1  g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g321(.A(G106gat), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT8), .B1(new_n205), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n522), .B(new_n524), .C1(G85gat), .C2(G92gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(G99gat), .B(G106gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n517), .A2(new_n520), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n515), .A2(new_n516), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT95), .B1(new_n506), .B2(new_n514), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n520), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n527), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G230gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(new_n356), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G120gat), .B(G148gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(G176gat), .B(G204gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT10), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n533), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n531), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n545), .A2(KEYINPUT10), .A3(new_n527), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n536), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n542), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI211_X1 g348(.A(KEYINPUT98), .B(new_n536), .C1(new_n544), .C2(new_n546), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n537), .B(new_n541), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n536), .B1(new_n544), .B2(new_n546), .ZN(new_n552));
  INV_X1    g351(.A(new_n537), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n540), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G15gat), .B(G22gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT16), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(G1gat), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(G1gat), .B2(new_n557), .ZN(new_n560));
  INV_X1    g359(.A(G8gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G43gat), .B(G50gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT90), .B(G29gat), .ZN(new_n564));
  INV_X1    g363(.A(G36gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(G29gat), .A2(G36gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT14), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT15), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(KEYINPUT92), .ZN(new_n570));
  INV_X1    g369(.A(new_n568), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n564), .B2(new_n565), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT15), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n313), .A2(G43gat), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(KEYINPUT91), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n563), .B(new_n569), .C1(new_n574), .C2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n570), .A2(new_n571), .A3(new_n577), .A4(new_n573), .ZN(new_n579));
  INV_X1    g378(.A(new_n563), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(KEYINPUT17), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n578), .A2(KEYINPUT17), .A3(new_n581), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n562), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n562), .B(KEYINPUT93), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n583), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT18), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n587), .B(new_n583), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n589), .B(KEYINPUT13), .Z(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n586), .A2(new_n588), .A3(KEYINPUT18), .A4(new_n589), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G113gat), .B(G141gat), .ZN(new_n598));
  INV_X1    g397(.A(G197gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT11), .B(G169gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n592), .A2(new_n603), .A3(new_n595), .A4(new_n596), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n503), .A2(new_n556), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(G183gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n562), .B(KEYINPUT93), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n545), .A2(KEYINPUT21), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n611), .A3(new_n613), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n615), .B(new_n616), .C1(KEYINPUT21), .C2(new_n545), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n545), .A2(KEYINPUT21), .ZN(new_n620));
  INV_X1    g419(.A(new_n616), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(new_n614), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n619), .B1(new_n617), .B2(new_n622), .ZN(new_n625));
  XNOR2_X1  g424(.A(G127gat), .B(G155gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G211gat), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n617), .A2(new_n622), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n618), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n631), .B2(new_n623), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n610), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n627), .B1(new_n624), .B2(new_n625), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n623), .A3(new_n629), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n609), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n532), .B1(new_n584), .B2(new_n585), .ZN(new_n638));
  NAND3_X1  g437(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n639));
  XOR2_X1   g438(.A(G190gat), .B(G218gat), .Z(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(KEYINPUT97), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n583), .B2(new_n527), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n640), .A2(KEYINPUT97), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n643), .A2(new_n644), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n645), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n648), .B1(new_n645), .B2(new_n649), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n608), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n455), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g457(.A1(new_n654), .A2(new_n417), .ZN(new_n659));
  NAND2_X1  g458(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n558), .A2(new_n561), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n664), .B(new_n665), .C1(new_n561), .C2(new_n659), .ZN(G1325gat));
  INV_X1    g465(.A(G15gat), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n654), .A2(new_n667), .A3(new_n501), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n655), .A2(new_n310), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n667), .B2(new_n669), .ZN(G1326gat));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n453), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT43), .B(G22gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  INV_X1    g472(.A(new_n607), .ZN(new_n674));
  AOI211_X1 g473(.A(new_n555), .B(new_n674), .C1(new_n633), .C2(new_n636), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n503), .A2(new_n652), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n656), .A3(new_n564), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT45), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n675), .B(KEYINPUT99), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n498), .A2(new_n681), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n390), .A2(new_n381), .B1(new_n455), .B2(new_n417), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n501), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n465), .B1(new_n497), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(new_n652), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n502), .B1(new_n486), .B2(new_n496), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n652), .B1(new_n689), .B2(new_n464), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT44), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n680), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n455), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n679), .B1(new_n564), .B2(new_n694), .ZN(G1328gat));
  NOR3_X1   g494(.A1(new_n676), .A2(G36gat), .A3(new_n417), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT46), .ZN(new_n697));
  OAI21_X1  g496(.A(G36gat), .B1(new_n693), .B2(new_n417), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1329gat));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n700));
  INV_X1    g499(.A(new_n310), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n676), .A2(G43gat), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n501), .ZN(new_n703));
  INV_X1    g502(.A(new_n680), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n687), .B1(new_n503), .B2(new_n652), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n501), .B1(new_n683), .B2(KEYINPUT100), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n452), .A2(KEYINPUT100), .A3(new_n456), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n486), .A2(new_n496), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n464), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n652), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(KEYINPUT44), .A3(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n702), .B1(new_n713), .B2(G43gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n700), .B1(new_n714), .B2(KEYINPUT47), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716));
  INV_X1    g515(.A(G43gat), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n692), .B2(new_n703), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT101), .B(new_n716), .C1(new_n718), .C2(new_n702), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n692), .A2(KEYINPUT102), .A3(new_n703), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(G43gat), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n702), .A2(new_n716), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n724), .A2(KEYINPUT103), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT103), .B1(new_n724), .B2(new_n725), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n720), .B1(new_n726), .B2(new_n727), .ZN(G1330gat));
  NAND3_X1  g527(.A1(new_n692), .A2(G50gat), .A3(new_n452), .ZN(new_n729));
  NAND2_X1  g528(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n313), .B1(new_n676), .B2(new_n453), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n732), .B(new_n733), .Z(G1331gat));
  NAND4_X1  g533(.A1(new_n686), .A2(new_n653), .A3(new_n555), .A4(new_n674), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(new_n455), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT105), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(new_n518), .ZN(G1332gat));
  AOI211_X1 g537(.A(new_n417), .B(new_n735), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1333gat));
  OAI21_X1  g540(.A(new_n508), .B1(new_n735), .B2(new_n701), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n735), .A2(new_n508), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n743), .A2(KEYINPUT106), .A3(new_n703), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT106), .B1(new_n743), .B2(new_n703), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n735), .A2(new_n453), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n509), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n637), .A2(new_n674), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n556), .B(new_n750), .C1(new_n688), .C2(new_n691), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n656), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(KEYINPUT107), .A3(new_n656), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(G85gat), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n686), .A2(KEYINPUT108), .A3(new_n652), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n710), .B2(new_n711), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n634), .A2(new_n635), .A3(new_n609), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n609), .B1(new_n634), .B2(new_n635), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n607), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n757), .A2(new_n759), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n757), .A2(new_n759), .A3(KEYINPUT51), .A4(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n455), .A2(G85gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n555), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n756), .A2(new_n770), .ZN(G1336gat));
  NOR2_X1   g570(.A1(new_n417), .A2(G92gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n768), .A2(new_n555), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  INV_X1    g573(.A(new_n417), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n751), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(G92gat), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n773), .B(new_n774), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n772), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n556), .B(new_n779), .C1(new_n766), .C2(new_n767), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n777), .B1(new_n751), .B2(new_n775), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT52), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(G1337gat));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n205), .A3(new_n310), .A4(new_n555), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n751), .A2(new_n703), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(new_n205), .ZN(G1338gat));
  AOI21_X1  g585(.A(new_n523), .B1(new_n751), .B2(new_n452), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n452), .A2(new_n523), .A3(new_n555), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT109), .Z(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n766), .B2(new_n767), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n787), .A2(new_n791), .A3(KEYINPUT53), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT53), .B1(new_n787), .B2(new_n791), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1339gat));
  NAND3_X1  g593(.A1(new_n544), .A2(new_n536), .A3(new_n546), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n795), .B(KEYINPUT54), .C1(new_n549), .C2(new_n550), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n541), .B1(new_n552), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n551), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT110), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n798), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n799), .A2(new_n805), .A3(new_n551), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n801), .A2(new_n607), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n593), .A2(new_n594), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n589), .B1(new_n586), .B2(new_n588), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n602), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n606), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n555), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n652), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n801), .A2(new_n804), .A3(new_n806), .A4(new_n811), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n711), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n637), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n762), .A2(new_n711), .A3(new_n556), .A4(new_n674), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n455), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n452), .B1(new_n460), .B2(new_n461), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n417), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n253), .A3(new_n607), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n823));
  INV_X1    g622(.A(new_n418), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n818), .A2(KEYINPUT111), .A3(new_n824), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n607), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n823), .B1(new_n831), .B2(G113gat), .ZN(new_n832));
  AOI211_X1 g631(.A(KEYINPUT112), .B(new_n253), .C1(new_n830), .C2(new_n607), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n822), .B1(new_n832), .B2(new_n833), .ZN(G1340gat));
  OAI21_X1  g633(.A(G120gat), .B1(new_n829), .B2(new_n556), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n821), .A2(new_n251), .A3(new_n555), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1341gat));
  AOI21_X1  g636(.A(G127gat), .B1(new_n821), .B2(new_n762), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n637), .A2(new_n266), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n830), .B2(new_n839), .ZN(G1342gat));
  NOR3_X1   g639(.A1(new_n820), .A2(G134gat), .A3(new_n711), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT56), .ZN(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n829), .B2(new_n711), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1343gat));
  AOI21_X1  g643(.A(new_n453), .B1(new_n816), .B2(new_n817), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n656), .A3(new_n501), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n674), .A2(G141gat), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT114), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n850), .A2(new_n775), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n845), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n806), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n805), .B1(new_n799), .B2(new_n551), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n858), .A2(new_n652), .A3(new_n804), .A4(new_n811), .ZN(new_n859));
  XNOR2_X1  g658(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n802), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n607), .A2(new_n861), .A3(new_n551), .A4(new_n799), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n652), .B1(new_n862), .B2(new_n812), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n762), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n633), .A2(new_n636), .A3(new_n711), .A4(new_n674), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n555), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n452), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n703), .A2(new_n455), .A3(new_n775), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(G141gat), .B1(new_n871), .B2(new_n674), .ZN(new_n872));
  XNOR2_X1  g671(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n846), .A2(new_n775), .A3(new_n852), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  OAI22_X1  g676(.A1(new_n853), .A2(new_n874), .B1(new_n876), .B2(new_n877), .ZN(G1344gat));
  INV_X1    g677(.A(new_n850), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n556), .A2(G148gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n417), .A3(new_n880), .ZN(new_n881));
  MUX2_X1   g680(.A(new_n868), .B(new_n845), .S(KEYINPUT57), .Z(new_n882));
  NAND4_X1  g681(.A1(new_n882), .A2(KEYINPUT119), .A3(new_n555), .A4(new_n870), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n854), .B(new_n453), .C1(new_n816), .C2(new_n817), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n637), .B1(new_n815), .B2(new_n863), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n817), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n452), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n555), .B(new_n870), .C1(new_n884), .C2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n883), .A2(new_n890), .A3(G148gat), .ZN(new_n891));
  XOR2_X1   g690(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n892));
  AND2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n894), .B(G148gat), .C1(new_n871), .C2(new_n556), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n895), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n881), .B1(new_n893), .B2(new_n897), .ZN(G1345gat));
  INV_X1    g697(.A(G155gat), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n871), .A2(new_n899), .A3(new_n637), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n879), .A2(new_n762), .A3(new_n417), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n899), .ZN(G1346gat));
  INV_X1    g701(.A(G162gat), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n879), .A2(new_n903), .A3(new_n652), .A4(new_n417), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n871), .A2(new_n711), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT120), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n904), .B1(new_n906), .B2(new_n903), .ZN(G1347gat));
  AOI21_X1  g706(.A(new_n656), .B1(new_n816), .B2(new_n817), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n775), .A3(new_n819), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n909), .A2(KEYINPUT121), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(KEYINPUT121), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n674), .A2(G169gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n816), .A2(new_n817), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n656), .A2(new_n417), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT122), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n914), .A2(new_n453), .A3(new_n310), .A4(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n674), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT123), .ZN(G1348gat));
  INV_X1    g719(.A(G176gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n917), .A2(new_n921), .A3(new_n556), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n910), .A2(new_n911), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n555), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n922), .B1(new_n924), .B2(new_n921), .ZN(G1349gat));
  NOR2_X1   g724(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n926));
  INV_X1    g725(.A(new_n909), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n762), .A3(new_n242), .ZN(new_n928));
  OAI21_X1  g727(.A(G183gat), .B1(new_n917), .B2(new_n637), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n930), .B(new_n931), .Z(G1350gat));
  NAND3_X1  g731(.A1(new_n923), .A2(new_n244), .A3(new_n652), .ZN(new_n933));
  OAI21_X1  g732(.A(G190gat), .B1(new_n917), .B2(new_n711), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1351gat));
  AND2_X1   g735(.A1(new_n916), .A2(new_n501), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n882), .A2(new_n937), .ZN(new_n938));
  OR3_X1    g737(.A1(new_n938), .A2(KEYINPUT126), .A3(new_n674), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT126), .B1(new_n938), .B2(new_n674), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(G197gat), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n501), .A2(new_n775), .A3(new_n452), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n908), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(new_n599), .A3(new_n607), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n941), .A2(new_n947), .ZN(G1352gat));
  INV_X1    g747(.A(G204gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n949), .A3(new_n555), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n950), .A2(KEYINPUT127), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(KEYINPUT127), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n952), .B1(new_n951), .B2(new_n953), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n882), .A2(new_n555), .A3(new_n937), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n954), .A2(new_n955), .B1(new_n949), .B2(new_n956), .ZN(G1353gat));
  NAND3_X1  g756(.A1(new_n946), .A2(new_n321), .A3(new_n762), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n882), .A2(new_n762), .A3(new_n937), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1354gat));
  OAI21_X1  g761(.A(G218gat), .B1(new_n938), .B2(new_n711), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n322), .A3(new_n652), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


