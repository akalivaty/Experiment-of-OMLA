

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789;

  NOR2_X1 U372 ( .A1(n647), .A2(n646), .ZN(n652) );
  XNOR2_X1 U373 ( .A(G125), .B(G146), .ZN(n506) );
  NOR2_X1 U374 ( .A1(G953), .A2(G237), .ZN(n552) );
  INV_X1 U375 ( .A(G953), .ZN(n776) );
  NAND2_X2 U376 ( .A1(n663), .A2(n660), .ZN(n397) );
  NOR2_X2 U377 ( .A1(n417), .A2(n416), .ZN(n748) );
  XNOR2_X2 U378 ( .A(n449), .B(n650), .ZN(n483) );
  XNOR2_X2 U379 ( .A(n613), .B(n479), .ZN(n635) );
  NOR2_X2 U380 ( .A1(n740), .A2(G902), .ZN(n498) );
  XNOR2_X2 U381 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n424) );
  XNOR2_X2 U382 ( .A(KEYINPUT18), .B(KEYINPUT90), .ZN(n423) );
  INV_X1 U383 ( .A(G137), .ZN(n490) );
  NOR2_X1 U384 ( .A1(n390), .A2(n388), .ZN(n387) );
  NOR2_X1 U385 ( .A1(n372), .A2(n370), .ZN(n369) );
  NAND2_X1 U386 ( .A1(n440), .A2(n353), .ZN(n474) );
  NAND2_X1 U387 ( .A1(n452), .A2(n451), .ZN(n450) );
  XNOR2_X1 U388 ( .A(n458), .B(n457), .ZN(n789) );
  XNOR2_X1 U389 ( .A(n459), .B(KEYINPUT41), .ZN(n712) );
  XNOR2_X1 U390 ( .A(n478), .B(n477), .ZN(n713) );
  XNOR2_X1 U391 ( .A(n640), .B(KEYINPUT1), .ZN(n699) );
  NOR2_X1 U392 ( .A1(n585), .A2(n413), .ZN(n412) );
  XNOR2_X1 U393 ( .A(n456), .B(n512), .ZN(n617) );
  OR2_X1 U394 ( .A1(n746), .A2(G902), .ZN(n456) );
  XOR2_X1 U395 ( .A(G131), .B(G140), .Z(n510) );
  INV_X1 U396 ( .A(G146), .ZN(n491) );
  AND2_X2 U397 ( .A1(n775), .A2(n662), .ZN(n349) );
  BUF_X1 U398 ( .A(n635), .Z(n350) );
  BUF_X1 U399 ( .A(n421), .Z(n351) );
  XNOR2_X2 U400 ( .A(n618), .B(n462), .ZN(n641) );
  XNOR2_X1 U401 ( .A(n404), .B(n586), .ZN(n653) );
  XNOR2_X1 U402 ( .A(n648), .B(KEYINPUT38), .ZN(n716) );
  XNOR2_X1 U403 ( .A(n412), .B(n411), .ZN(n404) );
  INV_X1 U404 ( .A(KEYINPUT88), .ZN(n411) );
  INV_X1 U405 ( .A(n715), .ZN(n413) );
  NOR2_X1 U406 ( .A1(n752), .A2(G902), .ZN(n541) );
  XNOR2_X1 U407 ( .A(n496), .B(G469), .ZN(n497) );
  XNOR2_X1 U408 ( .A(n473), .B(n471), .ZN(n749) );
  XNOR2_X1 U409 ( .A(n515), .B(n472), .ZN(n471) );
  XNOR2_X1 U410 ( .A(n516), .B(KEYINPUT103), .ZN(n472) );
  XNOR2_X1 U411 ( .A(n406), .B(n354), .ZN(n405) );
  XNOR2_X1 U412 ( .A(n476), .B(KEYINPUT108), .ZN(n718) );
  NOR2_X1 U413 ( .A1(n602), .A2(n616), .ZN(n476) );
  INV_X1 U414 ( .A(n595), .ZN(n383) );
  XOR2_X1 U415 ( .A(n749), .B(KEYINPUT121), .Z(n750) );
  XOR2_X1 U416 ( .A(n746), .B(KEYINPUT59), .Z(n747) );
  NOR2_X1 U417 ( .A1(n683), .A2(n625), .ZN(n443) );
  NAND2_X1 U418 ( .A1(n360), .A2(n352), .ZN(n435) );
  INV_X1 U419 ( .A(KEYINPUT85), .ZN(n465) );
  INV_X1 U420 ( .A(G237), .ZN(n563) );
  INV_X1 U421 ( .A(KEYINPUT109), .ZN(n462) );
  XNOR2_X1 U422 ( .A(G113), .B(KEYINPUT73), .ZN(n556) );
  XNOR2_X1 U423 ( .A(G137), .B(G128), .ZN(n529) );
  XNOR2_X1 U424 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U425 ( .A(KEYINPUT95), .B(KEYINPUT74), .Z(n525) );
  NAND2_X1 U426 ( .A1(n581), .A2(G214), .ZN(n715) );
  INV_X1 U427 ( .A(n716), .ZN(n460) );
  INV_X1 U428 ( .A(n403), .ZN(n410) );
  INV_X1 U429 ( .A(KEYINPUT35), .ZN(n479) );
  NOR2_X1 U430 ( .A1(n622), .A2(n463), .ZN(n709) );
  AND2_X1 U431 ( .A1(n718), .A2(n702), .ZN(n484) );
  NAND2_X1 U432 ( .A1(n389), .A2(n394), .ZN(n388) );
  AND2_X1 U433 ( .A1(n398), .A2(n367), .ZN(n390) );
  NAND2_X1 U434 ( .A1(n371), .A2(n394), .ZN(n370) );
  AND2_X1 U435 ( .A1(n398), .A2(n366), .ZN(n372) );
  NAND2_X1 U436 ( .A1(n713), .A2(n718), .ZN(n459) );
  NAND2_X1 U437 ( .A1(n441), .A2(n444), .ZN(n378) );
  NAND2_X1 U438 ( .A1(n656), .A2(n445), .ZN(n444) );
  NAND2_X1 U439 ( .A1(n443), .A2(n442), .ZN(n441) );
  INV_X1 U440 ( .A(KEYINPUT46), .ZN(n434) );
  INV_X1 U441 ( .A(KEYINPUT10), .ZN(n505) );
  XNOR2_X1 U442 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n636) );
  NOR2_X1 U443 ( .A1(n606), .A2(n599), .ZN(n642) );
  XOR2_X1 U444 ( .A(KEYINPUT94), .B(n510), .Z(n769) );
  XNOR2_X1 U445 ( .A(G119), .B(G110), .ZN(n523) );
  XNOR2_X1 U446 ( .A(G116), .B(G107), .ZN(n516) );
  INV_X1 U447 ( .A(G134), .ZN(n489) );
  XNOR2_X1 U448 ( .A(G122), .B(KEYINPUT9), .ZN(n513) );
  XNOR2_X1 U449 ( .A(G104), .B(G122), .ZN(n501) );
  XOR2_X1 U450 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n502) );
  XOR2_X1 U451 ( .A(KEYINPUT102), .B(KEYINPUT12), .Z(n500) );
  XNOR2_X1 U452 ( .A(n379), .B(n475), .ZN(n482) );
  INV_X1 U453 ( .A(KEYINPUT48), .ZN(n475) );
  XNOR2_X1 U454 ( .A(n435), .B(KEYINPUT77), .ZN(n380) );
  NAND2_X1 U455 ( .A1(n705), .A2(n463), .ZN(n706) );
  XNOR2_X1 U456 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n608) );
  XNOR2_X1 U457 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n550) );
  INV_X1 U458 ( .A(G101), .ZN(n756) );
  XNOR2_X1 U459 ( .A(KEYINPUT16), .B(G122), .ZN(n576) );
  AND2_X1 U460 ( .A1(n474), .A2(n365), .ZN(n418) );
  OR2_X1 U461 ( .A1(n775), .A2(n364), .ZN(n414) );
  INV_X1 U462 ( .A(KEYINPUT114), .ZN(n477) );
  NAND2_X1 U463 ( .A1(n716), .A2(n715), .ZN(n478) );
  XNOR2_X1 U464 ( .A(n436), .B(KEYINPUT78), .ZN(n649) );
  NOR2_X1 U465 ( .A1(n619), .A2(n599), .ZN(n601) );
  BUF_X1 U466 ( .A(n606), .Z(n703) );
  XNOR2_X1 U467 ( .A(n520), .B(n521), .ZN(n616) );
  XNOR2_X1 U468 ( .A(n529), .B(n528), .ZN(n530) );
  INV_X1 U469 ( .A(KEYINPUT42), .ZN(n457) );
  INV_X1 U470 ( .A(KEYINPUT115), .ZN(n407) );
  NAND2_X1 U471 ( .A1(n383), .A2(n382), .ZN(n598) );
  AND2_X1 U472 ( .A1(n596), .A2(n607), .ZN(n382) );
  XNOR2_X1 U473 ( .A(n624), .B(n623), .ZN(n695) );
  BUF_X1 U474 ( .A(G143), .Z(n605) );
  NOR2_X2 U475 ( .A1(n655), .A2(n654), .ZN(n690) );
  XNOR2_X1 U476 ( .A(n469), .B(n468), .ZN(n694) );
  INV_X1 U477 ( .A(KEYINPUT107), .ZN(n468) );
  AND2_X1 U478 ( .A1(n617), .A2(n616), .ZN(n469) );
  AND2_X1 U479 ( .A1(n620), .A2(n621), .ZN(n683) );
  INV_X1 U480 ( .A(KEYINPUT122), .ZN(n392) );
  NAND2_X1 U481 ( .A1(n386), .A2(n750), .ZN(n385) );
  INV_X1 U482 ( .A(KEYINPUT60), .ZN(n374) );
  NAND2_X1 U483 ( .A1(n386), .A2(n747), .ZN(n368) );
  OR2_X1 U484 ( .A1(KEYINPUT47), .A2(n658), .ZN(n352) );
  AND2_X1 U485 ( .A1(n482), .A2(n361), .ZN(n353) );
  XOR2_X1 U486 ( .A(n511), .B(n510), .Z(n354) );
  XNOR2_X1 U487 ( .A(G472), .B(KEYINPUT76), .ZN(n355) );
  AND2_X1 U488 ( .A1(n697), .A2(n665), .ZN(n356) );
  AND2_X1 U489 ( .A1(n681), .A2(n628), .ZN(n357) );
  AND2_X1 U490 ( .A1(n378), .A2(n357), .ZN(n358) );
  AND2_X1 U491 ( .A1(n480), .A2(n698), .ZN(n359) );
  XOR2_X1 U492 ( .A(n466), .B(n465), .Z(n360) );
  AND2_X1 U493 ( .A1(n666), .A2(n665), .ZN(n361) );
  BUF_X1 U494 ( .A(n699), .Z(n438) );
  XOR2_X1 U495 ( .A(KEYINPUT89), .B(KEYINPUT33), .Z(n362) );
  XOR2_X1 U496 ( .A(n651), .B(KEYINPUT113), .Z(n363) );
  NAND2_X1 U497 ( .A1(n661), .A2(KEYINPUT66), .ZN(n364) );
  OR2_X1 U498 ( .A1(n661), .A2(KEYINPUT66), .ZN(n365) );
  NOR2_X1 U499 ( .A1(n747), .A2(n373), .ZN(n366) );
  NOR2_X1 U500 ( .A1(n750), .A2(n391), .ZN(n367) );
  INV_X1 U501 ( .A(KEYINPUT66), .ZN(n662) );
  AND2_X1 U502 ( .A1(n671), .A2(G953), .ZN(n755) );
  INV_X1 U503 ( .A(n755), .ZN(n394) );
  NAND2_X1 U504 ( .A1(n369), .A2(n368), .ZN(n375) );
  NAND2_X1 U505 ( .A1(n747), .A2(n373), .ZN(n371) );
  INV_X1 U506 ( .A(G475), .ZN(n373) );
  XNOR2_X1 U507 ( .A(n375), .B(n374), .ZN(G60) );
  AND2_X1 U508 ( .A1(n378), .A2(n681), .ZN(n629) );
  NAND2_X1 U509 ( .A1(n376), .A2(n358), .ZN(n455) );
  NAND2_X1 U510 ( .A1(n377), .A2(n615), .ZN(n376) );
  XNOR2_X1 U511 ( .A(n635), .B(n614), .ZN(n377) );
  NAND2_X1 U512 ( .A1(n384), .A2(n627), .ZN(n681) );
  NAND2_X1 U513 ( .A1(n482), .A2(n356), .ZN(n659) );
  NAND2_X1 U514 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U515 ( .A1(n429), .A2(n428), .ZN(n381) );
  NOR2_X1 U516 ( .A1(n595), .A2(n480), .ZN(n384) );
  NAND2_X1 U517 ( .A1(n387), .A2(n385), .ZN(n393) );
  INV_X1 U518 ( .A(n398), .ZN(n386) );
  NAND2_X1 U519 ( .A1(n750), .A2(n391), .ZN(n389) );
  INV_X1 U520 ( .A(G478), .ZN(n391) );
  XNOR2_X1 U521 ( .A(n393), .B(n392), .ZN(G63) );
  XNOR2_X2 U522 ( .A(n485), .B(KEYINPUT22), .ZN(n595) );
  XNOR2_X1 U523 ( .A(n560), .B(n559), .ZN(n668) );
  NAND2_X1 U524 ( .A1(n359), .A2(n699), .ZN(n481) );
  XNOR2_X2 U525 ( .A(n395), .B(n396), .ZN(n421) );
  NOR2_X2 U526 ( .A1(n653), .A2(n591), .ZN(n395) );
  XOR2_X1 U527 ( .A(n592), .B(KEYINPUT0), .Z(n396) );
  NAND2_X1 U528 ( .A1(n789), .A2(n434), .ZN(n432) );
  NAND2_X1 U529 ( .A1(n431), .A2(n786), .ZN(n429) );
  NOR2_X1 U530 ( .A1(n734), .A2(n439), .ZN(n735) );
  NOR2_X1 U531 ( .A1(n417), .A2(n416), .ZN(n398) );
  INV_X1 U532 ( .A(n731), .ZN(n399) );
  BUF_X1 U533 ( .A(n618), .Z(n400) );
  XNOR2_X1 U534 ( .A(n397), .B(n637), .ZN(n401) );
  BUF_X1 U535 ( .A(n675), .Z(n402) );
  XNOR2_X1 U536 ( .A(n397), .B(n637), .ZN(n420) );
  INV_X1 U537 ( .A(n506), .ZN(n570) );
  XNOR2_X1 U538 ( .A(n770), .B(n527), .ZN(n531) );
  BUF_X1 U539 ( .A(n653), .Z(n654) );
  XNOR2_X1 U540 ( .A(n583), .B(n582), .ZN(n585) );
  OR2_X1 U541 ( .A1(n638), .A2(n404), .ZN(n403) );
  XNOR2_X1 U542 ( .A(n405), .B(n770), .ZN(n746) );
  XNOR2_X2 U543 ( .A(n509), .B(KEYINPUT71), .ZN(n770) );
  XNOR2_X1 U544 ( .A(n504), .B(n503), .ZN(n406) );
  XNOR2_X2 U545 ( .A(n408), .B(n407), .ZN(n786) );
  NAND2_X1 U546 ( .A1(n409), .A2(n438), .ZN(n408) );
  XNOR2_X1 U547 ( .A(n410), .B(KEYINPUT36), .ZN(n409) );
  NAND2_X2 U548 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X2 U549 ( .A(n659), .B(KEYINPUT87), .ZN(n775) );
  OR2_X2 U550 ( .A1(n420), .A2(n364), .ZN(n415) );
  NAND2_X1 U551 ( .A1(n419), .A2(n418), .ZN(n417) );
  NAND2_X1 U552 ( .A1(n349), .A2(n401), .ZN(n419) );
  NAND2_X1 U553 ( .A1(n421), .A2(n723), .ZN(n609) );
  NAND2_X1 U554 ( .A1(n421), .A2(n484), .ZN(n485) );
  NAND2_X1 U555 ( .A1(n351), .A2(n709), .ZN(n624) );
  AND2_X1 U556 ( .A1(n351), .A2(n702), .ZN(n620) );
  XNOR2_X1 U557 ( .A(n422), .B(n571), .ZN(n573) );
  XNOR2_X1 U558 ( .A(n424), .B(n423), .ZN(n422) );
  NAND2_X1 U559 ( .A1(n425), .A2(n630), .ZN(n464) );
  NAND2_X1 U560 ( .A1(n425), .A2(n632), .ZN(n633) );
  XNOR2_X1 U561 ( .A(n425), .B(G119), .ZN(G21) );
  XNOR2_X2 U562 ( .A(n598), .B(n597), .ZN(n425) );
  NAND2_X1 U563 ( .A1(n430), .A2(n426), .ZN(n428) );
  NOR2_X1 U564 ( .A1(n788), .A2(n427), .ZN(n426) );
  INV_X1 U565 ( .A(n786), .ZN(n427) );
  NOR2_X1 U566 ( .A1(n789), .A2(n434), .ZN(n430) );
  NAND2_X1 U567 ( .A1(n433), .A2(n432), .ZN(n431) );
  NAND2_X1 U568 ( .A1(n788), .A2(n434), .ZN(n433) );
  XNOR2_X1 U569 ( .A(n447), .B(n600), .ZN(n446) );
  NAND2_X1 U570 ( .A1(n641), .A2(n715), .ZN(n447) );
  INV_X2 U571 ( .A(G143), .ZN(n488) );
  NAND2_X1 U572 ( .A1(n446), .A2(n601), .ZN(n436) );
  XNOR2_X1 U573 ( .A(n437), .B(n757), .ZN(n675) );
  XNOR2_X1 U574 ( .A(n574), .B(n575), .ZN(n437) );
  INV_X1 U575 ( .A(n474), .ZN(n439) );
  INV_X1 U576 ( .A(n730), .ZN(n440) );
  INV_X1 U577 ( .A(n695), .ZN(n442) );
  INV_X1 U578 ( .A(n625), .ZN(n445) );
  XNOR2_X2 U579 ( .A(n448), .B(n363), .ZN(n788) );
  NAND2_X1 U580 ( .A1(n483), .A2(n692), .ZN(n448) );
  NOR2_X2 U581 ( .A1(n649), .A2(n460), .ZN(n449) );
  XNOR2_X2 U582 ( .A(n450), .B(n636), .ZN(n663) );
  NAND2_X1 U583 ( .A1(n455), .A2(n454), .ZN(n451) );
  NAND2_X1 U584 ( .A1(n453), .A2(KEYINPUT44), .ZN(n452) );
  NAND2_X1 U585 ( .A1(n634), .A2(n350), .ZN(n453) );
  NAND2_X1 U586 ( .A1(n464), .A2(n629), .ZN(n454) );
  NAND2_X1 U587 ( .A1(n712), .A2(n652), .ZN(n458) );
  XNOR2_X2 U588 ( .A(n461), .B(n490), .ZN(n774) );
  XNOR2_X1 U589 ( .A(n461), .B(n519), .ZN(n473) );
  XNOR2_X2 U590 ( .A(n571), .B(n489), .ZN(n461) );
  XNOR2_X1 U591 ( .A(n618), .B(KEYINPUT6), .ZN(n607) );
  INV_X1 U592 ( .A(n400), .ZN(n463) );
  XNOR2_X2 U593 ( .A(n561), .B(n355), .ZN(n618) );
  NAND2_X1 U594 ( .A1(n467), .A2(n657), .ZN(n466) );
  NAND2_X1 U595 ( .A1(n658), .A2(KEYINPUT47), .ZN(n467) );
  NAND2_X1 U596 ( .A1(n714), .A2(n690), .ZN(n658) );
  NOR2_X1 U597 ( .A1(n692), .A2(n694), .ZN(n656) );
  XNOR2_X2 U598 ( .A(n470), .B(KEYINPUT106), .ZN(n692) );
  NOR2_X1 U599 ( .A1(n617), .A2(n616), .ZN(n470) );
  INV_X1 U600 ( .A(n350), .ZN(n787) );
  NAND2_X1 U601 ( .A1(n698), .A2(n699), .ZN(n622) );
  INV_X1 U602 ( .A(n607), .ZN(n480) );
  XNOR2_X2 U603 ( .A(n481), .B(n362), .ZN(n723) );
  NAND2_X1 U604 ( .A1(n483), .A2(n694), .ZN(n697) );
  BUF_X1 U605 ( .A(n748), .Z(n751) );
  XNOR2_X1 U606 ( .A(n560), .B(n577), .ZN(n494) );
  XNOR2_X2 U607 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n768) );
  XNOR2_X2 U608 ( .A(n488), .B(G128), .ZN(n571) );
  INV_X1 U609 ( .A(KEYINPUT69), .ZN(n614) );
  INV_X1 U610 ( .A(KEYINPUT24), .ZN(n528) );
  XNOR2_X1 U611 ( .A(n573), .B(n572), .ZN(n574) );
  INV_X1 U612 ( .A(KEYINPUT30), .ZN(n600) );
  XNOR2_X1 U613 ( .A(n643), .B(KEYINPUT111), .ZN(n644) );
  XNOR2_X1 U614 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U615 ( .A(n495), .B(n494), .ZN(n740) );
  XNOR2_X1 U616 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U617 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n623) );
  XOR2_X1 U618 ( .A(n769), .B(KEYINPUT80), .Z(n487) );
  NAND2_X1 U619 ( .A1(G227), .A2(n776), .ZN(n486) );
  XNOR2_X1 U620 ( .A(n487), .B(n486), .ZN(n495) );
  XNOR2_X1 U621 ( .A(n768), .B(n756), .ZN(n572) );
  XNOR2_X1 U622 ( .A(n572), .B(n491), .ZN(n492) );
  XNOR2_X2 U623 ( .A(n774), .B(n492), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G110), .B(G107), .ZN(n493) );
  XNOR2_X1 U625 ( .A(n493), .B(G104), .ZN(n577) );
  INV_X1 U626 ( .A(KEYINPUT72), .ZN(n496) );
  XNOR2_X2 U627 ( .A(n498), .B(n497), .ZN(n640) );
  XNOR2_X1 U628 ( .A(KEYINPUT13), .B(G475), .ZN(n512) );
  NAND2_X1 U629 ( .A1(G214), .A2(n552), .ZN(n499) );
  XNOR2_X1 U630 ( .A(n500), .B(n499), .ZN(n504) );
  XNOR2_X1 U631 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U632 ( .A1(n570), .A2(KEYINPUT10), .ZN(n508) );
  NAND2_X1 U633 ( .A1(n506), .A2(n505), .ZN(n507) );
  NAND2_X1 U634 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U635 ( .A(n605), .B(G113), .ZN(n511) );
  XNOR2_X1 U636 ( .A(KEYINPUT105), .B(G478), .ZN(n521) );
  XOR2_X1 U637 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n514) );
  XNOR2_X1 U638 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U639 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n518) );
  NAND2_X1 U640 ( .A1(G234), .A2(n776), .ZN(n517) );
  XNOR2_X1 U641 ( .A(n518), .B(n517), .ZN(n522) );
  NAND2_X1 U642 ( .A1(G217), .A2(n522), .ZN(n519) );
  NOR2_X1 U643 ( .A1(G902), .A2(n749), .ZN(n520) );
  NAND2_X1 U644 ( .A1(G221), .A2(n522), .ZN(n533) );
  XOR2_X1 U645 ( .A(KEYINPUT23), .B(G140), .Z(n524) );
  XNOR2_X1 U646 ( .A(n524), .B(n523), .ZN(n526) );
  XNOR2_X1 U647 ( .A(n533), .B(n532), .ZN(n752) );
  XOR2_X1 U648 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n539) );
  XOR2_X1 U649 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n537) );
  XNOR2_X1 U650 ( .A(G902), .B(KEYINPUT91), .ZN(n535) );
  INV_X1 U651 ( .A(KEYINPUT15), .ZN(n534) );
  XNOR2_X1 U652 ( .A(n535), .B(n534), .ZN(n580) );
  NAND2_X1 U653 ( .A1(G234), .A2(n580), .ZN(n536) );
  XNOR2_X1 U654 ( .A(n537), .B(n536), .ZN(n547) );
  AND2_X1 U655 ( .A1(n547), .A2(G217), .ZN(n538) );
  XNOR2_X1 U656 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X2 U657 ( .A(n541), .B(n540), .ZN(n606) );
  NAND2_X1 U658 ( .A1(G234), .A2(G237), .ZN(n542) );
  XNOR2_X1 U659 ( .A(n542), .B(KEYINPUT14), .ZN(n544) );
  NAND2_X1 U660 ( .A1(G902), .A2(n544), .ZN(n587) );
  NOR2_X1 U661 ( .A1(G900), .A2(n587), .ZN(n543) );
  NAND2_X1 U662 ( .A1(n543), .A2(G953), .ZN(n546) );
  NAND2_X1 U663 ( .A1(G952), .A2(n544), .ZN(n545) );
  XNOR2_X1 U664 ( .A(KEYINPUT93), .B(n545), .ZN(n727) );
  NAND2_X1 U665 ( .A1(n727), .A2(n776), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n546), .A2(n590), .ZN(n549) );
  AND2_X1 U667 ( .A1(n547), .A2(G221), .ZN(n548) );
  XNOR2_X1 U668 ( .A(n548), .B(KEYINPUT21), .ZN(n702) );
  NAND2_X1 U669 ( .A1(n549), .A2(n702), .ZN(n599) );
  XOR2_X1 U670 ( .A(G131), .B(KEYINPUT5), .Z(n551) );
  XNOR2_X1 U671 ( .A(n551), .B(n550), .ZN(n554) );
  NAND2_X1 U672 ( .A1(n552), .A2(G210), .ZN(n553) );
  XNOR2_X1 U673 ( .A(n554), .B(n553), .ZN(n558) );
  XNOR2_X1 U674 ( .A(G119), .B(G116), .ZN(n555) );
  XNOR2_X1 U675 ( .A(n555), .B(KEYINPUT3), .ZN(n557) );
  XNOR2_X1 U676 ( .A(n557), .B(n556), .ZN(n578) );
  XNOR2_X1 U677 ( .A(n558), .B(n578), .ZN(n559) );
  INV_X1 U678 ( .A(G902), .ZN(n564) );
  NAND2_X1 U679 ( .A1(n668), .A2(n564), .ZN(n561) );
  AND2_X1 U680 ( .A1(n642), .A2(n480), .ZN(n562) );
  NAND2_X1 U681 ( .A1(n692), .A2(n562), .ZN(n638) );
  INV_X1 U682 ( .A(n638), .ZN(n565) );
  NAND2_X1 U683 ( .A1(n564), .A2(n563), .ZN(n581) );
  NAND2_X1 U684 ( .A1(n565), .A2(n715), .ZN(n566) );
  NOR2_X1 U685 ( .A1(n438), .A2(n566), .ZN(n567) );
  XNOR2_X1 U686 ( .A(n567), .B(KEYINPUT43), .ZN(n584) );
  NAND2_X1 U687 ( .A1(n776), .A2(G224), .ZN(n568) );
  XNOR2_X1 U688 ( .A(n568), .B(KEYINPUT81), .ZN(n569) );
  XNOR2_X1 U689 ( .A(n570), .B(n569), .ZN(n575) );
  XNOR2_X1 U690 ( .A(n577), .B(n576), .ZN(n579) );
  XNOR2_X1 U691 ( .A(n579), .B(n578), .ZN(n757) );
  INV_X1 U692 ( .A(n580), .ZN(n660) );
  NOR2_X1 U693 ( .A1(n675), .A2(n660), .ZN(n583) );
  AND2_X1 U694 ( .A1(n581), .A2(G210), .ZN(n582) );
  BUF_X1 U695 ( .A(n585), .Z(n648) );
  INV_X1 U696 ( .A(n648), .ZN(n604) );
  OR2_X1 U697 ( .A1(n584), .A2(n604), .ZN(n665) );
  XNOR2_X1 U698 ( .A(n665), .B(G140), .ZN(G42) );
  XNOR2_X1 U699 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n586) );
  INV_X1 U700 ( .A(n587), .ZN(n588) );
  NOR2_X1 U701 ( .A1(G898), .A2(n776), .ZN(n758) );
  NAND2_X1 U702 ( .A1(n588), .A2(n758), .ZN(n589) );
  AND2_X1 U703 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U704 ( .A(KEYINPUT68), .ZN(n592) );
  INV_X1 U705 ( .A(n617), .ZN(n602) );
  INV_X1 U706 ( .A(n438), .ZN(n639) );
  NOR2_X1 U707 ( .A1(n703), .A2(n641), .ZN(n593) );
  NAND2_X1 U708 ( .A1(n639), .A2(n593), .ZN(n594) );
  OR2_X1 U709 ( .A1(n595), .A2(n594), .ZN(n630) );
  XNOR2_X1 U710 ( .A(n630), .B(G110), .ZN(G12) );
  INV_X1 U711 ( .A(n703), .ZN(n626) );
  AND2_X1 U712 ( .A1(n438), .A2(n626), .ZN(n596) );
  XNOR2_X1 U713 ( .A(KEYINPUT82), .B(KEYINPUT32), .ZN(n597) );
  NAND2_X1 U714 ( .A1(n606), .A2(n640), .ZN(n619) );
  NAND2_X1 U715 ( .A1(n602), .A2(n616), .ZN(n610) );
  NOR2_X1 U716 ( .A1(n649), .A2(n610), .ZN(n603) );
  NAND2_X1 U717 ( .A1(n604), .A2(n603), .ZN(n657) );
  XNOR2_X1 U718 ( .A(n657), .B(n605), .ZN(G45) );
  INV_X1 U719 ( .A(KEYINPUT44), .ZN(n615) );
  AND2_X1 U720 ( .A1(n702), .A2(n606), .ZN(n698) );
  XNOR2_X1 U721 ( .A(n609), .B(n608), .ZN(n612) );
  INV_X1 U722 ( .A(n610), .ZN(n611) );
  NAND2_X1 U723 ( .A1(n612), .A2(n611), .ZN(n613) );
  INV_X1 U724 ( .A(KEYINPUT67), .ZN(n628) );
  NOR2_X1 U725 ( .A1(n619), .A2(n400), .ZN(n621) );
  NOR2_X1 U726 ( .A1(KEYINPUT44), .A2(n628), .ZN(n625) );
  NOR2_X1 U727 ( .A1(n438), .A2(n626), .ZN(n627) );
  INV_X1 U728 ( .A(n630), .ZN(n631) );
  NOR2_X1 U729 ( .A1(n631), .A2(KEYINPUT69), .ZN(n632) );
  NAND2_X1 U730 ( .A1(n633), .A2(n628), .ZN(n634) );
  INV_X1 U731 ( .A(KEYINPUT86), .ZN(n637) );
  XOR2_X1 U732 ( .A(n640), .B(KEYINPUT110), .Z(n647) );
  NAND2_X1 U733 ( .A1(n642), .A2(n641), .ZN(n645) );
  XOR2_X1 U734 ( .A(KEYINPUT28), .B(KEYINPUT112), .Z(n643) );
  INV_X1 U735 ( .A(KEYINPUT39), .ZN(n650) );
  INV_X1 U736 ( .A(KEYINPUT40), .ZN(n651) );
  INV_X1 U737 ( .A(n652), .ZN(n655) );
  INV_X1 U738 ( .A(n656), .ZN(n714) );
  NAND2_X1 U739 ( .A1(n660), .A2(KEYINPUT2), .ZN(n661) );
  INV_X1 U740 ( .A(n663), .ZN(n730) );
  NAND2_X1 U741 ( .A1(KEYINPUT2), .A2(n697), .ZN(n664) );
  XNOR2_X1 U742 ( .A(KEYINPUT83), .B(n664), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n748), .A2(G472), .ZN(n670) );
  XNOR2_X1 U744 ( .A(KEYINPUT116), .B(KEYINPUT62), .ZN(n667) );
  XNOR2_X1 U745 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n670), .B(n669), .ZN(n672) );
  INV_X1 U747 ( .A(G952), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n672), .A2(n394), .ZN(n673) );
  XNOR2_X1 U749 ( .A(n673), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U750 ( .A1(n748), .A2(G210), .ZN(n677) );
  XNOR2_X1 U751 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n674) );
  XNOR2_X1 U752 ( .A(n402), .B(n674), .ZN(n676) );
  XNOR2_X1 U753 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U754 ( .A1(n678), .A2(n394), .ZN(n680) );
  INV_X1 U755 ( .A(KEYINPUT56), .ZN(n679) );
  XNOR2_X1 U756 ( .A(n680), .B(n679), .ZN(G51) );
  XNOR2_X1 U757 ( .A(G101), .B(n681), .ZN(G3) );
  NAND2_X1 U758 ( .A1(n692), .A2(n683), .ZN(n682) );
  XNOR2_X1 U759 ( .A(n682), .B(G104), .ZN(G6) );
  XOR2_X1 U760 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n685) );
  NAND2_X1 U761 ( .A1(n683), .A2(n694), .ZN(n684) );
  XNOR2_X1 U762 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U763 ( .A(G107), .B(n686), .ZN(G9) );
  XOR2_X1 U764 ( .A(KEYINPUT29), .B(KEYINPUT117), .Z(n688) );
  NAND2_X1 U765 ( .A1(n690), .A2(n694), .ZN(n687) );
  XNOR2_X1 U766 ( .A(n688), .B(n687), .ZN(n689) );
  XOR2_X1 U767 ( .A(G128), .B(n689), .Z(G30) );
  NAND2_X1 U768 ( .A1(n690), .A2(n692), .ZN(n691) );
  XNOR2_X1 U769 ( .A(n691), .B(G146), .ZN(G48) );
  NAND2_X1 U770 ( .A1(n695), .A2(n692), .ZN(n693) );
  XNOR2_X1 U771 ( .A(n693), .B(G113), .ZN(G15) );
  NAND2_X1 U772 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U773 ( .A(n696), .B(G116), .ZN(G18) );
  XNOR2_X1 U774 ( .A(G134), .B(n697), .ZN(G36) );
  NAND2_X1 U775 ( .A1(n712), .A2(n723), .ZN(n738) );
  XNOR2_X1 U776 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n701) );
  NOR2_X1 U777 ( .A1(n438), .A2(n698), .ZN(n700) );
  XNOR2_X1 U778 ( .A(n701), .B(n700), .ZN(n707) );
  NOR2_X1 U779 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U780 ( .A(KEYINPUT49), .B(n704), .ZN(n705) );
  NOR2_X1 U781 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U782 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U783 ( .A(KEYINPUT51), .B(n710), .ZN(n711) );
  NAND2_X1 U784 ( .A1(n712), .A2(n711), .ZN(n725) );
  NAND2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n721) );
  NOR2_X1 U786 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U787 ( .A(KEYINPUT119), .B(n717), .ZN(n719) );
  NAND2_X1 U788 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U789 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U791 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U792 ( .A(n726), .B(KEYINPUT52), .ZN(n728) );
  NAND2_X1 U793 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U794 ( .A1(n729), .A2(n776), .ZN(n736) );
  INV_X1 U795 ( .A(n775), .ZN(n731) );
  NOR2_X1 U796 ( .A1(n731), .A2(n730), .ZN(n733) );
  XNOR2_X1 U797 ( .A(KEYINPUT84), .B(KEYINPUT2), .ZN(n732) );
  NOR2_X1 U798 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U799 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U800 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U801 ( .A(KEYINPUT53), .B(n739), .Z(G75) );
  NAND2_X1 U802 ( .A1(n751), .A2(G469), .ZN(n744) );
  XOR2_X1 U803 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n742) );
  XNOR2_X1 U804 ( .A(n740), .B(KEYINPUT120), .ZN(n741) );
  XNOR2_X1 U805 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U806 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U807 ( .A1(n755), .A2(n745), .ZN(G54) );
  NAND2_X1 U808 ( .A1(n751), .A2(G217), .ZN(n753) );
  XNOR2_X1 U809 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U810 ( .A1(n755), .A2(n754), .ZN(G66) );
  XNOR2_X1 U811 ( .A(n757), .B(n756), .ZN(n759) );
  NOR2_X1 U812 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U813 ( .A(KEYINPUT124), .B(n760), .ZN(n767) );
  NAND2_X1 U814 ( .A1(n440), .A2(n776), .ZN(n765) );
  XOR2_X1 U815 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n762) );
  NAND2_X1 U816 ( .A1(G224), .A2(G953), .ZN(n761) );
  XNOR2_X1 U817 ( .A(n762), .B(n761), .ZN(n763) );
  NAND2_X1 U818 ( .A1(n763), .A2(G898), .ZN(n764) );
  NAND2_X1 U819 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U820 ( .A(n767), .B(n766), .ZN(G69) );
  XNOR2_X1 U821 ( .A(n769), .B(n768), .ZN(n772) );
  XNOR2_X1 U822 ( .A(n770), .B(KEYINPUT125), .ZN(n771) );
  XNOR2_X1 U823 ( .A(n772), .B(n771), .ZN(n773) );
  XNOR2_X1 U824 ( .A(n774), .B(n773), .ZN(n779) );
  XOR2_X1 U825 ( .A(n779), .B(n399), .Z(n777) );
  NAND2_X1 U826 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U827 ( .A(n778), .B(KEYINPUT126), .ZN(n784) );
  XNOR2_X1 U828 ( .A(G227), .B(n779), .ZN(n780) );
  NAND2_X1 U829 ( .A1(n780), .A2(G900), .ZN(n781) );
  XOR2_X1 U830 ( .A(KEYINPUT127), .B(n781), .Z(n782) );
  NAND2_X1 U831 ( .A1(n782), .A2(G953), .ZN(n783) );
  NAND2_X1 U832 ( .A1(n784), .A2(n783), .ZN(G72) );
  XOR2_X1 U833 ( .A(G125), .B(KEYINPUT37), .Z(n785) );
  XNOR2_X1 U834 ( .A(n786), .B(n785), .ZN(G27) );
  XOR2_X1 U835 ( .A(n787), .B(G122), .Z(G24) );
  XOR2_X1 U836 ( .A(n788), .B(G131), .Z(G33) );
  XOR2_X1 U837 ( .A(G137), .B(n789), .Z(G39) );
endmodule

