//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n532, new_n533, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT66), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT67), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  XNOR2_X1  g028(.A(G325), .B(KEYINPUT68), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  INV_X1    g030(.A(G2105), .ZN(new_n456));
  AND2_X1   g031(.A1(new_n456), .A2(G2104), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G101), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(new_n456), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n459), .A2(new_n460), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(G160));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G112), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n466), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n466), .A2(new_n456), .ZN(new_n480));
  AOI211_X1 g055(.A(new_n476), .B(new_n479), .C1(G124), .C2(new_n480), .ZN(G162));
  OR2_X1    g056(.A1(G102), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G114), .C2(new_n456), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n462), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n480), .A2(G126), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n477), .A2(KEYINPUT4), .A3(G138), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n484), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  INV_X1    g066(.A(G543), .ZN(new_n492));
  OR2_X1    g067(.A1(KEYINPUT6), .A2(G651), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT6), .A2(G651), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G50), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n493), .A2(new_n494), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(new_n492), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g077(.A(KEYINPUT71), .B(G88), .Z(new_n503));
  OAI21_X1  g078(.A(new_n496), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n504), .A2(new_n507), .ZN(G166));
  NAND3_X1  g083(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n495), .A2(G51), .ZN(new_n510));
  NAND3_X1  g085(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT7), .ZN(new_n512));
  INV_X1    g087(.A(G89), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n502), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n509), .B(new_n510), .C1(new_n514), .C2(KEYINPUT72), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n514), .A2(KEYINPUT72), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(G168));
  NAND2_X1  g092(.A1(new_n495), .A2(G52), .ZN(new_n518));
  INV_X1    g093(.A(G90), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n502), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n506), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n520), .A2(new_n522), .ZN(G171));
  NAND2_X1  g098(.A1(new_n495), .A2(G43), .ZN(new_n524));
  INV_X1    g099(.A(G81), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n502), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n506), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G860), .ZN(G153));
  NAND4_X1  g105(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g106(.A1(G1), .A2(G3), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT8), .ZN(new_n533));
  NAND4_X1  g108(.A1(G319), .A2(G483), .A3(G661), .A4(new_n533), .ZN(G188));
  AND2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  NOR3_X1   g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT73), .B1(new_n499), .B2(new_n500), .ZN(new_n539));
  OAI21_X1  g114(.A(G65), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(G78), .A2(G543), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(KEYINPUT74), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n543));
  INV_X1    g118(.A(G65), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n537), .B1(new_n535), .B2(new_n536), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n500), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n541), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n542), .A2(new_n549), .A3(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n495), .A2(G53), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n495), .A2(new_n553), .A3(G53), .ZN(new_n554));
  INV_X1    g129(.A(new_n502), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n552), .A2(new_n554), .B1(G91), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n550), .A2(KEYINPUT75), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT75), .B1(new_n550), .B2(new_n556), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n557), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND2_X1  g137(.A1(new_n495), .A2(G49), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT76), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n501), .A2(G74), .ZN(new_n565));
  AOI22_X1  g140(.A1(G87), .A2(new_n555), .B1(new_n565), .B2(G651), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(G288));
  AND2_X1   g142(.A1(new_n555), .A2(G86), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(new_n501), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(G48), .B2(new_n495), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n570), .A2(new_n571), .A3(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(G72), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G60), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n506), .B1(new_n580), .B2(KEYINPUT78), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n581), .B1(KEYINPUT78), .B2(new_n580), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n555), .A2(G85), .B1(G47), .B2(new_n495), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n555), .A2(KEYINPUT10), .A3(G92), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n587));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n502), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n545), .B2(new_n546), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT79), .Z(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n495), .A2(G54), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n585), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n585), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT80), .Z(new_n602));
  INV_X1    g177(.A(G299), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(G868), .B2(new_n603), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(G868), .B2(new_n603), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n529), .ZN(G323));
  XOR2_X1   g185(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n611));
  XNOR2_X1  g186(.A(G323), .B(new_n611), .ZN(G282));
  NAND2_X1  g187(.A1(new_n461), .A2(new_n457), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT82), .B(G2100), .Z(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT83), .Z(new_n618));
  NAND2_X1  g193(.A1(new_n477), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n480), .A2(G123), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n456), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G2096), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n618), .B(new_n625), .C1(new_n616), .C2(new_n615), .ZN(G156));
  INV_X1    g201(.A(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n632), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT84), .B(G2100), .Z(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n646), .B2(KEYINPUT18), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n624), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT20), .Z(new_n664));
  OR2_X1    g239(.A1(new_n658), .A2(new_n659), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(new_n660), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n666), .A2(KEYINPUT86), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(KEYINPUT86), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(new_n662), .ZN(new_n669));
  OAI221_X1 g244(.A(new_n664), .B1(new_n665), .B2(new_n662), .C1(new_n667), .C2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1991), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G229));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G303), .B2(G16), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT90), .B(G1971), .Z(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT32), .B(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(new_n685));
  MUX2_X1   g260(.A(G6), .B(G305), .S(G16), .Z(new_n686));
  OAI21_X1  g261(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n678), .A2(G23), .ZN(new_n688));
  INV_X1    g263(.A(G288), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(new_n678), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT33), .ZN(new_n691));
  INV_X1    g266(.A(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n687), .B(new_n693), .C1(new_n685), .C2(new_n686), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT34), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n477), .A2(G131), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n480), .A2(G119), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n456), .A2(G107), .ZN(new_n700));
  OAI21_X1  g275(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n698), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G25), .B(new_n702), .S(G29), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n678), .A2(G24), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT87), .Z(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G290), .B2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G1986), .Z(new_n710));
  NOR4_X1   g285(.A1(new_n696), .A2(new_n697), .A3(new_n706), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT36), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n678), .A2(G20), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT23), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n603), .B2(new_n678), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1956), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G35), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G162), .B2(new_n717), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT29), .Z(new_n720));
  INV_X1    g295(.A(G2090), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G4), .A2(G16), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n598), .B2(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G1348), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n720), .A2(new_n721), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n717), .A2(G32), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n457), .A2(G105), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT94), .Z(new_n730));
  INV_X1    g305(.A(G141), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n462), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n480), .A2(G129), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(KEYINPUT26), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(KEYINPUT26), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n728), .B1(new_n738), .B2(new_n717), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G1341), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n529), .A2(new_n678), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n678), .B2(G19), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n741), .B1(new_n742), .B2(new_n744), .C1(G1348), .C2(new_n724), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n717), .B1(new_n746), .B2(G34), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(KEYINPUT93), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(KEYINPUT93), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n746), .B2(G34), .ZN(new_n750));
  AOI22_X1  g325(.A1(G160), .A2(G29), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2084), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n727), .A2(new_n745), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n678), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n678), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(G164), .A2(G29), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G27), .B2(G29), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n717), .A2(G33), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n456), .A2(G103), .A3(G2104), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT92), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT25), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n477), .A2(G139), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n765), .B(new_n766), .C1(new_n456), .C2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G2072), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n759), .A2(new_n760), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n761), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n678), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n678), .ZN(new_n775));
  INV_X1    g350(.A(G1961), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n744), .A2(new_n742), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT31), .B(G11), .Z(new_n779));
  NOR2_X1   g354(.A1(new_n623), .A2(new_n717), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT30), .B(G28), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n779), .B(new_n780), .C1(new_n717), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n777), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n717), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT91), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n477), .A2(G140), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n480), .A2(G128), .ZN(new_n788));
  OR2_X1    g363(.A1(G104), .A2(G2105), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n789), .B(G2104), .C1(G116), .C2(new_n456), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n786), .B1(new_n792), .B2(new_n717), .ZN(new_n793));
  INV_X1    g368(.A(G2067), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n770), .B2(G2072), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n773), .A2(new_n783), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n753), .A2(new_n757), .A3(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n712), .A2(new_n716), .A3(new_n798), .ZN(G311));
  OR3_X1    g374(.A1(new_n712), .A2(new_n716), .A3(new_n798), .ZN(G150));
  NAND2_X1  g375(.A1(new_n598), .A2(G559), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT38), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n495), .A2(G55), .ZN(new_n803));
  INV_X1    g378(.A(G93), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n502), .B2(new_n804), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n506), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n529), .A2(new_n808), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n528), .A2(new_n526), .B1(new_n805), .B2(new_n807), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n802), .B(new_n811), .Z(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  INV_X1    g388(.A(G860), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n808), .A2(new_n814), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT96), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(G145));
  XNOR2_X1  g396(.A(G162), .B(new_n623), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G160), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n490), .B(new_n791), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n768), .ZN(new_n825));
  INV_X1    g400(.A(new_n738), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n702), .B(KEYINPUT97), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n614), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n480), .A2(G130), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n456), .A2(G118), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G142), .B2(new_n477), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n829), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n827), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n827), .A2(new_n835), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n823), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G37), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n836), .A2(KEYINPUT98), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n838), .A2(new_n823), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n836), .A2(KEYINPUT98), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n841), .A2(KEYINPUT99), .A3(new_n845), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g426(.A(G290), .B(G288), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT102), .ZN(new_n853));
  XNOR2_X1  g428(.A(G305), .B(G166), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n854), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT42), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n550), .A2(new_n556), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT75), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n550), .A2(KEYINPUT75), .A3(new_n556), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n864), .A3(new_n598), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT100), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n863), .A2(new_n867), .A3(new_n864), .A4(new_n598), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n866), .A2(new_n868), .B1(new_n603), .B2(new_n597), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n597), .B1(new_n557), .B2(new_n558), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT101), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n872), .B(new_n597), .C1(new_n557), .C2(new_n558), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n867), .B1(G299), .B2(new_n598), .ZN(new_n874));
  INV_X1    g449(.A(new_n868), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n871), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(new_n866), .B2(new_n868), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n876), .A2(new_n877), .B1(new_n878), .B2(new_n870), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n608), .B(new_n811), .Z(new_n880));
  MUX2_X1   g455(.A(new_n869), .B(new_n879), .S(new_n880), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n860), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G868), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(G868), .B2(new_n808), .ZN(G331));
  XNOR2_X1  g459(.A(G331), .B(KEYINPUT103), .ZN(G295));
  OR2_X1    g460(.A1(new_n521), .A2(new_n506), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n555), .A2(G90), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n886), .A2(KEYINPUT104), .A3(new_n518), .A4(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n520), .B2(new_n522), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n811), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n890), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n810), .A3(new_n809), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n892), .A2(G168), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G168), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n869), .A2(new_n897), .A3(KEYINPUT106), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n900));
  INV_X1    g475(.A(new_n896), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(G168), .A3(new_n894), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n899), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n879), .B2(new_n903), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n871), .A2(new_n873), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n866), .A2(new_n868), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT41), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n909), .A2(KEYINPUT41), .A3(new_n870), .ZN(new_n911));
  OAI211_X1 g486(.A(KEYINPUT105), .B(new_n897), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n905), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n859), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(KEYINPUT43), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n908), .A2(new_n897), .A3(new_n878), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n900), .B1(new_n903), .B2(new_n877), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n859), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(G37), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n840), .B1(new_n913), .B2(new_n859), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g499(.A(KEYINPUT107), .B(new_n840), .C1(new_n913), .C2(new_n859), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n920), .B2(new_n914), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n925), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n930), .B2(new_n916), .ZN(new_n931));
  MUX2_X1   g506(.A(new_n928), .B(new_n931), .S(KEYINPUT44), .Z(G397));
  NAND2_X1  g507(.A1(G160), .A2(G40), .ZN(new_n933));
  INV_X1    g508(.A(G1384), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n490), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G8), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT113), .ZN(new_n939));
  OR2_X1    g514(.A1(G305), .A2(G1981), .ZN(new_n940));
  INV_X1    g515(.A(new_n576), .ZN(new_n941));
  OAI21_X1  g516(.A(G1981), .B1(new_n941), .B2(new_n568), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT115), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(KEYINPUT116), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT49), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n939), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n940), .A2(new_n942), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n944), .B1(KEYINPUT116), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n692), .A3(new_n689), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n939), .B1(new_n951), .B2(new_n940), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n939), .B1(G1976), .B2(new_n689), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n954), .B(new_n953), .C1(G1976), .C2(new_n689), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n956), .A2(KEYINPUT114), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(KEYINPUT114), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(G40), .B(G160), .C1(new_n935), .C2(KEYINPUT50), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n935), .A2(KEYINPUT50), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT112), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n935), .A2(new_n963), .A3(KEYINPUT50), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n960), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n721), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n935), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n933), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT108), .B(G1384), .Z(new_n970));
  NAND3_X1  g545(.A1(new_n490), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1971), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n937), .B1(new_n966), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G303), .A2(G8), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT55), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n975), .A2(new_n978), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT63), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G2084), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n965), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n490), .A2(KEYINPUT45), .A3(new_n934), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n968), .A2(new_n969), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n756), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(G8), .A3(G168), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT118), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n959), .A2(new_n979), .A3(new_n982), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n952), .B1(new_n991), .B2(KEYINPUT63), .ZN(new_n992));
  INV_X1    g567(.A(new_n979), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n968), .A2(new_n969), .A3(new_n760), .A4(new_n971), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n760), .A2(KEYINPUT53), .ZN(new_n997));
  OAI221_X1 g572(.A(new_n996), .B1(new_n997), .B2(new_n986), .C1(new_n965), .C2(G1961), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G171), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G168), .A2(new_n937), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1000), .B1(new_n1002), .B2(KEYINPUT122), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(G8), .B(new_n1004), .C1(new_n988), .C2(G286), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n965), .A2(new_n983), .B1(new_n986), .B2(new_n756), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1002), .B(new_n1003), .C1(new_n1006), .C2(new_n937), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT121), .B1(new_n988), .B2(new_n1001), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1006), .A2(new_n1009), .A3(new_n1002), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1005), .B(new_n1007), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n999), .B1(new_n1011), .B2(KEYINPUT62), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT62), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n1007), .A4(new_n1005), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n982), .A2(new_n979), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1012), .A2(new_n1015), .B1(new_n1016), .B2(new_n990), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n861), .B(KEYINPUT57), .Z(new_n1018));
  INV_X1    g593(.A(G1956), .ZN(new_n1019));
  INV_X1    g594(.A(new_n961), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(new_n960), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT56), .B(G2072), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n968), .A2(new_n969), .A3(new_n971), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1018), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n965), .ZN(new_n1026));
  INV_X1    g601(.A(G1348), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1026), .A2(new_n1027), .B1(new_n794), .B2(new_n936), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1025), .B1(new_n1028), .B2(new_n597), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1021), .A2(new_n1018), .A3(new_n1023), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT61), .B1(new_n1024), .B2(KEYINPUT120), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1032), .B1(new_n1024), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1996), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n968), .A2(new_n969), .A3(new_n1036), .A4(new_n971), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT58), .B(G1341), .Z(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n933), .B2(new_n935), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n529), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1035), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1025), .A2(KEYINPUT61), .A3(new_n1030), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n936), .A2(new_n794), .ZN(new_n1049));
  OAI211_X1 g624(.A(KEYINPUT60), .B(new_n1049), .C1(new_n965), .C2(G1348), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1050), .A2(new_n598), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1028), .A2(KEYINPUT60), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n598), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1048), .B(new_n1051), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1031), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1011), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1026), .A2(KEYINPUT123), .A3(new_n776), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n965), .B2(G1961), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n490), .A2(new_n970), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT45), .B1(new_n1061), .B2(KEYINPUT109), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(KEYINPUT109), .B2(new_n1061), .ZN(new_n1063));
  INV_X1    g638(.A(G40), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n464), .A2(new_n1064), .A3(new_n997), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n971), .A2(new_n469), .A3(new_n1065), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1063), .A2(new_n1066), .B1(new_n994), .B2(new_n995), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1060), .A2(G301), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n999), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1060), .A2(KEYINPUT124), .A3(new_n1067), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT124), .B1(new_n1060), .B2(new_n1067), .ZN(new_n1073));
  OAI21_X1  g648(.A(G171), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1069), .B1(new_n998), .B2(G301), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1017), .B1(new_n1056), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1020), .A2(new_n960), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n974), .B1(new_n1079), .B2(G2090), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n978), .B1(new_n1080), .B2(G8), .ZN(new_n1081));
  XOR2_X1   g656(.A(new_n1081), .B(KEYINPUT117), .Z(new_n1082));
  AOI21_X1  g657(.A(new_n993), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n959), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n992), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n702), .A2(new_n705), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n702), .A2(new_n705), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n933), .B(new_n1063), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1063), .A2(new_n933), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n826), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(new_n1036), .ZN(new_n1091));
  XOR2_X1   g666(.A(new_n1091), .B(KEYINPUT111), .Z(new_n1092));
  NAND2_X1  g667(.A1(new_n1089), .A2(new_n1036), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT110), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n738), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n791), .B(G2067), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1089), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1092), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(G290), .B(G1986), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1088), .B(new_n1098), .C1(new_n1089), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1085), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(G290), .A2(G1986), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1089), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT48), .Z(new_n1104));
  NOR3_X1   g679(.A1(new_n1098), .A2(new_n1088), .A3(new_n1104), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1094), .A2(KEYINPUT46), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n1107), .B(KEYINPUT125), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1094), .A2(KEYINPUT46), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT47), .Z(new_n1111));
  OAI22_X1  g686(.A1(new_n1098), .A2(new_n1086), .B1(G2067), .B2(new_n791), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n1105), .B(new_n1111), .C1(new_n1089), .C2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1101), .A2(new_n1113), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n1116));
  INV_X1    g690(.A(G227), .ZN(new_n1117));
  NAND2_X1  g691(.A1(new_n1117), .A2(G319), .ZN(new_n1118));
  XOR2_X1   g692(.A(new_n1118), .B(KEYINPUT126), .Z(new_n1119));
  INV_X1    g693(.A(new_n1119), .ZN(new_n1120));
  NAND3_X1  g694(.A1(new_n676), .A2(new_n641), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g695(.A(new_n1121), .B1(new_n848), .B2(new_n849), .ZN(new_n1122));
  AND3_X1   g696(.A1(new_n928), .A2(new_n1116), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g697(.A(new_n1116), .B1(new_n928), .B2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g698(.A1(new_n1123), .A2(new_n1124), .ZN(G308));
  NAND2_X1  g699(.A1(new_n928), .A2(new_n1122), .ZN(new_n1126));
  NAND2_X1  g700(.A1(new_n1126), .A2(KEYINPUT127), .ZN(new_n1127));
  NAND3_X1  g701(.A1(new_n928), .A2(new_n1116), .A3(new_n1122), .ZN(new_n1128));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1128), .ZN(G225));
endmodule


