//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n191), .B1(KEYINPUT0), .B2(G128), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n188), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT0), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT65), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n189), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT66), .B1(new_n193), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n190), .B1(new_n188), .B2(new_n192), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(new_n189), .A3(new_n201), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(G137), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT67), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n216), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n218), .A2(new_n210), .A3(new_n211), .A4(new_n213), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n203), .A2(new_n207), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT68), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n203), .A2(new_n223), .A3(new_n207), .A4(new_n220), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n196), .A2(G146), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n194), .A2(G143), .ZN(new_n227));
  OAI211_X1 g041(.A(G128), .B(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n210), .A2(new_n213), .A3(new_n215), .A4(new_n211), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n209), .A2(G137), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n212), .A2(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(G131), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n195), .B(new_n197), .C1(KEYINPUT1), .C2(new_n200), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n228), .A2(new_n229), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n222), .A2(new_n224), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT2), .A2(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT2), .A2(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT69), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT2), .A3(G113), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n238), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G116), .B(G119), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n243), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n217), .A2(KEYINPUT70), .A3(new_n219), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT70), .B1(new_n217), .B2(new_n219), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n204), .A2(new_n205), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n228), .A2(new_n233), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n229), .A2(new_n232), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT71), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n234), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT30), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n237), .A2(new_n247), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n257), .ZN(new_n261));
  INV_X1    g075(.A(new_n249), .ZN(new_n262));
  INV_X1    g076(.A(new_n250), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n217), .A2(KEYINPUT70), .A3(new_n219), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n261), .A2(new_n246), .A3(new_n265), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT72), .B(KEYINPUT27), .Z(new_n267));
  NOR2_X1   g081(.A1(G237), .A2(G953), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G101), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n260), .A2(new_n266), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT31), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n260), .A2(new_n275), .A3(new_n266), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n234), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n221), .B2(KEYINPUT68), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n246), .B1(new_n279), .B2(new_n224), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n266), .B1(new_n280), .B2(KEYINPUT73), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n282));
  AOI211_X1 g096(.A(new_n282), .B(new_n246), .C1(new_n279), .C2(new_n224), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT28), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n265), .A2(new_n234), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n247), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n265), .A2(KEYINPUT74), .A3(new_n234), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT28), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n272), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n187), .B1(new_n277), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n294), .A2(G472), .A3(G902), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n277), .B2(new_n292), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n300));
  INV_X1    g114(.A(new_n266), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n235), .A2(new_n236), .B1(new_n258), .B2(KEYINPUT30), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(new_n247), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n300), .B1(new_n303), .B2(new_n272), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT28), .B1(new_n287), .B2(new_n288), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n235), .A2(new_n247), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n282), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n280), .A2(KEYINPUT73), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(new_n266), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n305), .B1(new_n309), .B2(KEYINPUT28), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n304), .B1(new_n310), .B2(new_n272), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT76), .B(G902), .Z(new_n312));
  OAI21_X1  g126(.A(new_n247), .B1(new_n251), .B2(new_n257), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n266), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(KEYINPUT75), .B(new_n247), .C1(new_n251), .C2(new_n257), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(KEYINPUT28), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n291), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n272), .A2(KEYINPUT29), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n312), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G472), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n274), .B(new_n276), .C1(new_n310), .C2(new_n272), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(KEYINPUT77), .A3(new_n296), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n295), .A2(new_n299), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G110), .B(G140), .ZN(new_n325));
  INV_X1    g139(.A(G953), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(G227), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n325), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  INV_X1    g143(.A(G107), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G104), .ZN(new_n331));
  INV_X1    g145(.A(G104), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G107), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n331), .B2(KEYINPUT3), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT85), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n332), .A2(G107), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT85), .B(KEYINPUT3), .C1(new_n332), .C2(G107), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n334), .B1(new_n341), .B2(new_n329), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT10), .B1(new_n342), .B2(new_n252), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n330), .A2(G104), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n338), .B2(new_n337), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT85), .B1(new_n331), .B2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g160(.A(new_n340), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n345), .B(new_n329), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n334), .ZN(new_n349));
  AND4_X1   g163(.A1(KEYINPUT10), .A2(new_n252), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G101), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT4), .A3(new_n348), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n339), .A2(new_n340), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n329), .B1(new_n355), .B2(new_n345), .ZN(new_n356));
  XOR2_X1   g170(.A(KEYINPUT86), .B(KEYINPUT4), .Z(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT87), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n360));
  NOR4_X1   g174(.A1(new_n341), .A2(new_n360), .A3(new_n329), .A4(new_n357), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n263), .B(new_n354), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n248), .A2(new_n249), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n351), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n351), .B2(new_n362), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n328), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n252), .A2(new_n348), .A3(new_n349), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n348), .A2(new_n349), .B1(new_n233), .B2(new_n228), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT12), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n371), .B1(new_n217), .B2(new_n219), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n368), .B2(new_n369), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(KEYINPUT88), .B(new_n373), .C1(new_n368), .C2(new_n369), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n372), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n351), .A2(new_n362), .A3(new_n364), .ZN(new_n379));
  INV_X1    g193(.A(new_n328), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n367), .A2(new_n381), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT89), .B(G469), .Z(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n312), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n378), .A2(new_n379), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n328), .B(KEYINPUT84), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n366), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n379), .A3(new_n380), .ZN(new_n390));
  AOI21_X1  g204(.A(G902), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G469), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n385), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G221), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT9), .B(G234), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G902), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G478), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT15), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G116), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n330), .B1(new_n404), .B2(KEYINPUT14), .ZN(new_n405));
  INV_X1    g219(.A(G116), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G122), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n408), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT95), .B1(new_n196), .B2(G128), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT95), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n200), .A3(G143), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n196), .A2(G128), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n414), .A2(new_n209), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n209), .B1(new_n414), .B2(new_n415), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n409), .B(new_n410), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT13), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n196), .A2(KEYINPUT13), .A3(G128), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n414), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G134), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n414), .A2(new_n209), .A3(new_n415), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n408), .A2(G107), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n404), .A2(new_n407), .A3(new_n330), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n418), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G217), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n395), .A2(new_n430), .A3(G953), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n418), .A2(new_n428), .A3(new_n431), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n402), .B1(new_n435), .B2(new_n312), .ZN(new_n436));
  INV_X1    g250(.A(new_n312), .ZN(new_n437));
  AOI211_X1 g251(.A(new_n437), .B(new_n401), .C1(new_n433), .C2(new_n434), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(KEYINPUT90), .A2(G143), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(KEYINPUT90), .A2(G143), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n441), .A2(new_n442), .B1(new_n268), .B2(G214), .ZN(new_n443));
  INV_X1    g257(.A(G237), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n326), .A3(G214), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(new_n440), .ZN(new_n446));
  OAI21_X1  g260(.A(G131), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT17), .ZN(new_n448));
  INV_X1    g262(.A(new_n442), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n445), .B1(new_n449), .B2(new_n440), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n441), .A2(G214), .A3(new_n268), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(new_n215), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n447), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G125), .B(G140), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT16), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT16), .ZN(new_n456));
  INV_X1    g270(.A(G140), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(G125), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT79), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT79), .A4(G125), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n194), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n455), .A2(G146), .A3(new_n460), .A4(new_n461), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n215), .B1(new_n450), .B2(new_n451), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT17), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n453), .A2(new_n463), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G113), .B(G122), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(new_n332), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n454), .B(new_n194), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT18), .A2(G131), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n450), .A2(new_n451), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT18), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n470), .B(new_n472), .C1(new_n447), .C2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n467), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n469), .B1(new_n467), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n397), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT94), .B(G475), .Z(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n457), .A2(G125), .ZN(new_n483));
  INV_X1    g297(.A(G125), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G140), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n483), .A2(new_n485), .A3(KEYINPUT19), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT19), .B1(new_n483), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n194), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n443), .A2(new_n446), .A3(G131), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n464), .B(new_n488), .C1(new_n489), .C2(new_n465), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n474), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n469), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n491), .B1(new_n490), .B2(new_n474), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n475), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT92), .ZN(new_n497));
  NOR2_X1   g311(.A1(G475), .A2(G902), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT92), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n475), .B(new_n499), .C1(new_n494), .C2(new_n495), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT20), .ZN(new_n502));
  NOR3_X1   g316(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n496), .A2(KEYINPUT93), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT93), .B1(new_n496), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n482), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n393), .A2(new_n399), .A3(new_n439), .A4(new_n507), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n326), .B(new_n312), .C1(G234), .C2(G237), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT21), .B(G898), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G952), .ZN(new_n512));
  AOI211_X1 g326(.A(G953), .B(new_n512), .C1(G234), .C2(G237), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G214), .B1(G237), .B2(G902), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g332(.A(G119), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G116), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n518), .B(G113), .C1(KEYINPUT5), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n243), .A2(new_n244), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n348), .A2(new_n349), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n352), .A2(G101), .A3(new_n358), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n360), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n356), .A2(KEYINPUT87), .A3(new_n358), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT4), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n530), .B1(new_n352), .B2(G101), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n246), .B1(new_n531), .B2(new_n348), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n525), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(G110), .B(G122), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n517), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n525), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n359), .A2(new_n361), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n354), .A2(new_n247), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n534), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n250), .A2(G125), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(G125), .B2(new_n252), .ZN(new_n544));
  INV_X1    g358(.A(G224), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G953), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n544), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n539), .A2(new_n517), .A3(new_n540), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n542), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT7), .B1(new_n545), .B2(G953), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n544), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g365(.A(new_n534), .B(KEYINPUT8), .Z(new_n552));
  NAND2_X1  g366(.A1(new_n523), .A2(new_n524), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n536), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n533), .A2(new_n534), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G210), .B1(G237), .B2(G902), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n549), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n549), .B2(new_n557), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n515), .B(new_n516), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n508), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g376(.A(G119), .B(G128), .Z(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT24), .B(G110), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT78), .B1(new_n519), .B2(G128), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n566), .A2(KEYINPUT23), .B1(new_n519), .B2(G128), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(KEYINPUT23), .B2(new_n566), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n565), .B1(new_n568), .B2(G110), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n454), .A2(new_n194), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n464), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT22), .B(G137), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(KEYINPUT81), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n212), .A2(KEYINPUT22), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT22), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G137), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n574), .A2(new_n576), .A3(KEYINPUT81), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT82), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n576), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT81), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n572), .A2(KEYINPUT81), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT82), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G234), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n394), .A2(new_n586), .A3(G953), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n578), .A2(new_n587), .A3(new_n584), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n463), .A2(new_n464), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n563), .A2(new_n564), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n568), .B2(G110), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(KEYINPUT80), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT80), .B1(new_n592), .B2(new_n594), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n571), .B(new_n591), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n571), .ZN(new_n599));
  INV_X1    g413(.A(new_n597), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(new_n595), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT83), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n591), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n589), .A2(KEYINPUT83), .A3(new_n590), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n598), .B(new_n312), .C1(new_n601), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT25), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n571), .B1(new_n596), .B2(new_n597), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n604), .A3(new_n603), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n610), .A2(KEYINPUT25), .A3(new_n312), .A4(new_n598), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n430), .B1(new_n312), .B2(G234), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(G902), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n610), .A2(new_n615), .A3(new_n598), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n324), .A2(new_n562), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  AOI21_X1  g433(.A(new_n275), .B1(new_n303), .B2(new_n272), .ZN(new_n620));
  INV_X1    g434(.A(new_n276), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n284), .A2(new_n291), .ZN(new_n623));
  INV_X1    g437(.A(new_n272), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n437), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G472), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n293), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n365), .A2(new_n366), .A3(new_n328), .ZN(new_n629));
  INV_X1    g443(.A(new_n387), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n378), .B2(new_n379), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(G469), .B1(new_n632), .B2(G902), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n398), .B1(new_n633), .B2(new_n385), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n617), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT96), .B1(new_n628), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n312), .B1(new_n277), .B2(new_n292), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n637), .A2(G472), .B1(new_n322), .B2(new_n187), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT96), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n617), .A4(new_n634), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n502), .A2(new_n506), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n481), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n435), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n437), .A2(new_n400), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n434), .A2(KEYINPUT98), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n418), .A2(new_n428), .A3(new_n648), .A4(new_n431), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n429), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n418), .A2(new_n428), .A3(KEYINPUT97), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n432), .A3(new_n653), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n646), .A2(new_n650), .A3(new_n654), .A4(KEYINPUT33), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n431), .B1(new_n429), .B2(new_n651), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n643), .B1(new_n656), .B2(new_n653), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n646), .B1(new_n657), .B2(new_n650), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n644), .B(new_n645), .C1(new_n655), .C2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n435), .A2(new_n312), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n400), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n660), .B1(new_n659), .B2(new_n662), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n642), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n561), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n636), .A2(new_n640), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  NAND3_X1  g483(.A1(new_n497), .A2(new_n500), .A3(new_n503), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n502), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n481), .B1(new_n436), .B2(new_n438), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n561), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n636), .A2(new_n640), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT35), .B(G107), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G9));
  INV_X1    g491(.A(KEYINPUT36), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n605), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n601), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n615), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n614), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n508), .A2(new_n561), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n638), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n516), .B1(new_n559), .B2(new_n560), .ZN(new_n688));
  INV_X1    g502(.A(new_n673), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n513), .B1(new_n509), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n671), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n687), .B1(new_n688), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n516), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n549), .A2(new_n557), .ZN(new_n696));
  INV_X1    g510(.A(new_n558), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n549), .A2(new_n557), .A3(new_n558), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n695), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n691), .B(new_n673), .C1(new_n502), .C2(new_n670), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(KEYINPUT101), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n694), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n614), .A2(new_n681), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n399), .A3(new_n393), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n324), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  NAND2_X1  g522(.A1(new_n698), .A2(new_n699), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n507), .A2(new_n439), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n682), .A2(new_n712), .A3(new_n516), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n315), .A2(new_n316), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n397), .B1(new_n715), .B2(new_n272), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n303), .A2(new_n624), .ZN(new_n717));
  OAI21_X1  g531(.A(G472), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n295), .A2(new_n299), .A3(new_n323), .A4(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n691), .B(KEYINPUT39), .Z(new_n720));
  NAND2_X1  g534(.A1(new_n634), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n721), .A2(KEYINPUT40), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(KEYINPUT40), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n714), .A2(new_n719), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  OAI211_X1 g539(.A(new_n642), .B(new_n692), .C1(new_n663), .C2(new_n664), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n688), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n324), .A2(new_n727), .A3(new_n706), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  AOI21_X1  g543(.A(new_n437), .B1(new_n367), .B2(new_n381), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n385), .B(new_n399), .C1(new_n392), .C2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT103), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n382), .A2(new_n312), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(G469), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(KEYINPUT103), .A3(new_n399), .A4(new_n385), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n324), .A2(new_n737), .A3(new_n617), .A4(new_n666), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  NAND4_X1  g554(.A1(new_n324), .A2(new_n737), .A3(new_n617), .A4(new_n674), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  NOR2_X1   g556(.A1(new_n730), .A2(new_n392), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n437), .B(new_n383), .C1(new_n367), .C2(new_n381), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n398), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n700), .A3(KEYINPUT104), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT104), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n688), .B2(new_n731), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  AND4_X1   g563(.A1(new_n515), .A2(new_n704), .A3(new_n439), .A4(new_n507), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n324), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  AOI21_X1  g566(.A(new_n627), .B1(new_n322), .B2(new_n312), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n318), .A2(new_n624), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n274), .A3(new_n276), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(new_n187), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n614), .A2(new_n616), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n753), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n700), .A2(new_n712), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n758), .A2(new_n737), .A3(new_n515), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G122), .ZN(G24));
  NOR3_X1   g576(.A1(new_n753), .A2(new_n756), .A3(new_n682), .ZN(new_n763));
  INV_X1    g577(.A(new_n726), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n749), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  NAND3_X1  g580(.A1(new_n295), .A2(new_n321), .A3(new_n297), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n393), .A2(new_n399), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n698), .A2(new_n516), .A3(new_n699), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n767), .A2(new_n764), .A3(new_n617), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT42), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n726), .A2(new_n768), .A3(new_n769), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n324), .A3(new_n774), .A4(new_n617), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n215), .ZN(G33));
  NOR3_X1   g591(.A1(new_n768), .A2(new_n769), .A3(new_n693), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n324), .A2(new_n617), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  OAI21_X1  g594(.A(new_n507), .B1(new_n663), .B2(new_n664), .ZN(new_n781));
  XOR2_X1   g595(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  OAI221_X1 g598(.A(new_n507), .B1(KEYINPUT105), .B2(KEYINPUT43), .C1(new_n663), .C2(new_n664), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n784), .A2(new_n785), .A3(KEYINPUT106), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n638), .B2(new_n682), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n628), .A2(KEYINPUT107), .A3(new_n704), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n788), .A2(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT108), .B1(new_n793), .B2(KEYINPUT44), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n632), .A2(KEYINPUT45), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n629), .B2(new_n631), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(G469), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(G469), .A2(G902), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n799), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n385), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n769), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n399), .A3(new_n720), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n793), .B2(KEYINPUT44), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT108), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  INV_X1    g623(.A(new_n789), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT106), .B1(new_n784), .B2(new_n785), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n792), .A2(new_n791), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n808), .B(new_n809), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n794), .A2(new_n807), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  NOR4_X1   g630(.A1(new_n324), .A2(new_n617), .A3(new_n726), .A4(new_n769), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n399), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT47), .B1(new_n804), .B2(new_n399), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT109), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n822), .B(new_n817), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  INV_X1    g639(.A(new_n719), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n769), .A2(new_n731), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n617), .A2(new_n826), .A3(new_n513), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n659), .A2(new_n662), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT100), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n828), .A2(new_n642), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n514), .B1(new_n784), .B2(new_n785), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n749), .A3(new_n758), .ZN(new_n835));
  AND4_X1   g649(.A1(G952), .A2(new_n833), .A3(new_n326), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n827), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT116), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT48), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n767), .A2(new_n617), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n838), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n836), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n843), .A2(KEYINPUT118), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n711), .A2(new_n695), .A3(new_n745), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n834), .A2(new_n758), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n846), .B(KEYINPUT115), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n834), .A3(KEYINPUT50), .A4(new_n758), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n832), .A2(new_n642), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n850), .A2(new_n852), .B1(new_n828), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n818), .A2(new_n819), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n735), .A2(new_n385), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n399), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n849), .B2(new_n769), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n834), .A2(KEYINPUT114), .A3(new_n758), .A4(new_n805), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n838), .A2(new_n763), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n854), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n863), .A2(new_n864), .B1(new_n843), .B2(KEYINPUT118), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n854), .A2(KEYINPUT51), .A3(new_n861), .A4(new_n862), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n844), .B(new_n865), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n772), .A2(new_n775), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n439), .A2(new_n481), .A3(new_n692), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n502), .B2(new_n670), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n698), .A3(new_n516), .A4(new_n699), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n705), .A2(new_n873), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n773), .A2(new_n763), .B1(new_n324), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT111), .B1(new_n875), .B2(new_n779), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n637), .A2(G472), .B1(new_n187), .B2(new_n755), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n764), .A2(new_n770), .A3(new_n704), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n324), .A2(new_n874), .ZN(new_n879));
  AND4_X1   g693(.A1(KEYINPUT111), .A2(new_n779), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n870), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n738), .A2(new_n741), .A3(new_n751), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n761), .A2(new_n618), .A3(new_n684), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n507), .B1(new_n436), .B2(new_n438), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT110), .B1(new_n561), .B2(new_n884), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n561), .A2(new_n884), .A3(KEYINPUT110), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n636), .A2(new_n640), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n882), .A2(new_n883), .A3(new_n667), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n765), .A2(new_n707), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n768), .A2(new_n704), .A3(new_n691), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n719), .A2(new_n760), .A3(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n728), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT52), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n765), .A2(new_n707), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n728), .A2(new_n892), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n889), .A2(KEYINPUT53), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n733), .A2(new_n515), .A3(new_n736), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n759), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n902), .A2(new_n758), .B1(new_n683), .B2(new_n638), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n887), .A3(new_n618), .A4(new_n667), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n738), .A2(new_n741), .A3(new_n751), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n779), .A2(new_n878), .A3(new_n879), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT111), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n875), .A2(KEYINPUT111), .A3(new_n779), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n776), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT112), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n765), .A2(new_n707), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n765), .B2(new_n707), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n728), .A2(new_n892), .A3(KEYINPUT52), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT52), .B1(new_n890), .B2(new_n893), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT113), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n896), .A2(KEYINPUT112), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n765), .A2(new_n707), .A3(new_n913), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(KEYINPUT52), .A3(new_n921), .A4(new_n893), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT113), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n898), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n912), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n900), .B1(new_n925), .B2(KEYINPUT53), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT54), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n906), .A2(new_n911), .A3(KEYINPUT53), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n917), .A2(KEYINPUT113), .A3(new_n918), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n923), .B1(new_n922), .B2(new_n898), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n899), .A2(new_n906), .A3(new_n911), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT53), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT54), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  OAI22_X1  g750(.A1(new_n869), .A2(new_n936), .B1(G952), .B2(G953), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n856), .B(KEYINPUT49), .ZN(new_n938));
  NOR4_X1   g752(.A1(new_n938), .A2(new_n757), .A3(new_n695), .A4(new_n398), .ZN(new_n939));
  INV_X1    g753(.A(new_n781), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n939), .A2(new_n826), .A3(new_n711), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(new_n941), .ZN(G75));
  NAND2_X1  g756(.A1(new_n512), .A2(G953), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT120), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n932), .A2(new_n933), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n312), .B1(new_n931), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n697), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n542), .A2(new_n548), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n547), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  NOR2_X1   g765(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n952));
  AND2_X1   g766(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n944), .B1(new_n948), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT56), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n951), .B1(new_n947), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(G51));
  INV_X1    g772(.A(new_n944), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n799), .B(KEYINPUT57), .Z(new_n960));
  NAND3_X1  g774(.A1(new_n906), .A2(new_n911), .A3(KEYINPUT53), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n919), .B2(new_n924), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT53), .B1(new_n889), .B2(new_n899), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT54), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT121), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n931), .A2(new_n965), .A3(new_n934), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n965), .B1(new_n931), .B2(new_n934), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n960), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n382), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n946), .A2(G469), .A3(new_n795), .A4(new_n797), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n959), .B1(new_n970), .B2(new_n971), .ZN(G54));
  NAND3_X1  g786(.A1(new_n946), .A2(KEYINPUT58), .A3(G475), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n497), .A2(new_n500), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n959), .B1(new_n975), .B2(new_n976), .ZN(G60));
  NAND2_X1  g791(.A1(new_n935), .A2(KEYINPUT121), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n966), .A3(new_n964), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n644), .B1(new_n655), .B2(new_n658), .ZN(new_n980));
  NAND2_X1  g794(.A1(G478), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT59), .Z(new_n982));
  NOR2_X1   g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n959), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  AOI22_X1  g798(.A1(new_n926), .A2(KEYINPUT54), .B1(new_n931), .B2(new_n934), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n980), .B1(new_n985), .B2(new_n982), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(G63));
  NAND2_X1  g801(.A1(G217), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT60), .Z(new_n989));
  OAI211_X1 g803(.A(new_n680), .B(new_n989), .C1(new_n962), .C2(new_n963), .ZN(new_n990));
  NOR2_X1   g804(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n959), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n989), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n931), .B2(new_n945), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n610), .A2(new_n598), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT122), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n990), .B(new_n992), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(G66));
  OAI21_X1  g813(.A(G953), .B1(new_n510), .B2(new_n545), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n906), .B2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n949), .B1(G898), .B2(new_n326), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT124), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1001), .B(new_n1003), .ZN(G69));
  AOI21_X1  g818(.A(new_n326), .B1(G227), .B2(G900), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n486), .A2(new_n487), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n302), .B(new_n1008), .Z(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT125), .Z(new_n1010));
  NOR2_X1   g824(.A1(new_n721), .A2(new_n769), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n665), .A2(new_n884), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1011), .A2(new_n324), .A3(new_n617), .A4(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n815), .A2(new_n824), .A3(new_n1013), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n920), .A2(new_n724), .A3(new_n728), .A4(new_n921), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT62), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1010), .B1(new_n1019), .B2(G953), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G900), .A2(G953), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n804), .A2(new_n399), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1022), .A2(new_n720), .A3(new_n760), .A4(new_n840), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n870), .A2(new_n1023), .A3(new_n779), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n920), .A2(new_n728), .A3(new_n921), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n815), .A3(new_n824), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1021), .B(new_n1009), .C1(new_n1027), .C2(G953), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1007), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1018), .A2(new_n1017), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n815), .A2(new_n824), .A3(new_n1013), .ZN(new_n1031));
  AOI21_X1  g845(.A(G953), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1010), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1028), .B(new_n1007), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1006), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1028), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(KEYINPUT126), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1038), .A2(new_n1005), .A3(new_n1034), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1036), .A2(new_n1039), .ZN(G72));
  INV_X1    g854(.A(new_n717), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n303), .A2(new_n624), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  AND4_X1   g858(.A1(new_n1041), .A2(new_n926), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1019), .A2(new_n906), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1041), .B1(new_n1046), .B2(new_n1044), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1044), .B1(new_n1027), .B2(new_n888), .ZN(new_n1048));
  XOR2_X1   g862(.A(new_n1042), .B(KEYINPUT127), .Z(new_n1049));
  AND2_X1   g863(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NOR4_X1   g864(.A1(new_n1045), .A2(new_n1047), .A3(new_n959), .A4(new_n1050), .ZN(G57));
endmodule


