//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G116), .A2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G50), .B2(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G107), .ZN(new_n216));
  INV_X1    g0016(.A(G264), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n207), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NOR2_X1   g0023(.A1(new_n207), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  NAND3_X1  g0026(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n202), .A2(G50), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT64), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n223), .B(new_n226), .C1(new_n227), .C2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n215), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT67), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT16), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT70), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n250), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT70), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n255), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT7), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n251), .A2(KEYINPUT78), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT78), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT3), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(KEYINPUT7), .B(new_n256), .C1(new_n266), .C2(new_n254), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n219), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G159), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G58), .A2(G68), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT79), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n202), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n272), .B1(new_n276), .B2(G20), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n249), .B1(new_n268), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT72), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT72), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n280), .A2(new_n284), .A3(new_n281), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n263), .A2(new_n265), .A3(KEYINPUT3), .ZN(new_n287));
  AOI21_X1  g0087(.A(G20), .B1(new_n287), .B2(new_n257), .ZN(new_n288));
  OAI21_X1  g0088(.A(G68), .B1(new_n288), .B2(new_n261), .ZN(new_n289));
  AOI211_X1 g0089(.A(KEYINPUT7), .B(G20), .C1(new_n287), .C2(new_n257), .ZN(new_n290));
  OAI211_X1 g0090(.A(KEYINPUT16), .B(new_n277), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n279), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  OAI211_X1 g0093(.A(G1), .B(G13), .C1(new_n251), .C2(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(G223), .A2(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G226), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G1698), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n287), .A2(new_n257), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G87), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G45), .ZN(new_n301));
  AOI21_X1  g0101(.A(G1), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G274), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT68), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT69), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G41), .A2(G45), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT69), .B1(new_n307), .B2(G1), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n294), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(new_n215), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n300), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(KEYINPUT80), .A2(G190), .ZN(new_n312));
  NAND2_X1  g0112(.A1(KEYINPUT80), .A2(G190), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT8), .B(G58), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G13), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n319), .A2(new_n256), .A3(G1), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G1), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n286), .B1(new_n322), .B2(G20), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n321), .B1(new_n324), .B2(new_n318), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n311), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n292), .A2(new_n316), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT17), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n291), .A2(new_n286), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n325), .B1(new_n332), .B2(new_n279), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n333), .A2(KEYINPUT17), .A3(new_n316), .A4(new_n328), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT70), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT70), .B1(new_n257), .B2(new_n258), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT7), .B1(new_n338), .B2(new_n256), .ZN(new_n339));
  INV_X1    g0139(.A(new_n267), .ZN(new_n340));
  OAI21_X1  g0140(.A(G68), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT16), .B1(new_n341), .B2(new_n277), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n291), .A2(new_n286), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n326), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n300), .A2(new_n304), .ZN(new_n346));
  INV_X1    g0146(.A(new_n310), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  NOR4_X1   g0149(.A1(new_n304), .A2(new_n300), .A3(new_n310), .A4(new_n349), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT18), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT18), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n348), .A2(new_n350), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n333), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n335), .B(KEYINPUT81), .C1(new_n352), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT81), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n355), .A2(new_n352), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n331), .A2(new_n334), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n309), .A2(new_n220), .ZN(new_n363));
  INV_X1    g0163(.A(G1698), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n296), .A2(new_n364), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n365), .B1(G232), .B2(new_n364), .C1(new_n336), .C2(new_n337), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G33), .A2(G97), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n281), .B1(G33), .B2(G41), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n304), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n362), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n294), .B1(new_n366), .B2(new_n367), .ZN(new_n373));
  NOR4_X1   g0173(.A1(new_n373), .A2(KEYINPUT13), .A3(new_n304), .A4(new_n363), .ZN(new_n374));
  OAI21_X1  g0174(.A(G169), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT14), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(KEYINPUT77), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  OAI221_X1 g0178(.A(G169), .B1(KEYINPUT77), .B2(new_n376), .C1(new_n372), .C2(new_n374), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n372), .A2(new_n374), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n376), .A2(KEYINPUT77), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n378), .A2(new_n379), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n384));
  INV_X1    g0184(.A(G77), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n256), .A2(G33), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n286), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g0188(.A(new_n388), .B(KEYINPUT11), .Z(new_n389));
  NAND2_X1  g0189(.A1(new_n320), .A2(new_n219), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT12), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n324), .B2(new_n219), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n383), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n323), .A2(G77), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n320), .A2(new_n385), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n317), .A2(new_n270), .B1(new_n256), .B2(new_n385), .ZN(new_n398));
  XNOR2_X1  g0198(.A(KEYINPUT15), .B(G87), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(new_n386), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n286), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n255), .A2(new_n259), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(G232), .A3(new_n364), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n338), .A2(G107), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n403), .A2(G238), .A3(G1698), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT74), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n403), .A2(new_n408), .A3(G232), .A4(new_n364), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n405), .A2(new_n406), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n369), .ZN(new_n411));
  INV_X1    g0211(.A(new_n309), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G244), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n411), .A2(new_n349), .A3(new_n371), .A4(new_n413), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n411), .A2(new_n371), .A3(new_n413), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n402), .B(new_n414), .C1(new_n415), .C2(G169), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(G190), .ZN(new_n417));
  INV_X1    g0217(.A(new_n402), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n327), .C2(new_n415), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n395), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n361), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT10), .ZN(new_n422));
  INV_X1    g0222(.A(G150), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n317), .A2(new_n386), .B1(new_n423), .B2(new_n270), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT73), .ZN(new_n425));
  OAI21_X1  g0225(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT73), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n427), .B1(new_n270), .B2(new_n423), .C1(new_n317), .C2(new_n386), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G50), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n429), .A2(new_n286), .B1(new_n430), .B2(new_n320), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n323), .A2(G50), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT9), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(G222), .A2(G1698), .ZN(new_n436));
  OR2_X1    g0236(.A1(KEYINPUT71), .A2(G223), .ZN(new_n437));
  NAND2_X1  g0237(.A1(KEYINPUT71), .A2(G223), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n364), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n403), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n440), .B(new_n369), .C1(G77), .C2(new_n403), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n412), .A2(G226), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(G190), .A3(new_n442), .A4(new_n371), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n431), .A2(KEYINPUT9), .A3(new_n432), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n435), .A2(KEYINPUT76), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n441), .A2(new_n442), .A3(new_n371), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G200), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT75), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(KEYINPUT75), .A3(G200), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n435), .A2(new_n443), .A3(new_n444), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n422), .B(new_n445), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n452), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(new_n450), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n455), .C1(KEYINPUT76), .C2(KEYINPUT10), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n446), .A2(G179), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n446), .A2(new_n345), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n433), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n380), .A2(G190), .ZN(new_n460));
  OAI21_X1  g0260(.A(G200), .B1(new_n372), .B2(new_n374), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n393), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n453), .A2(new_n456), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT82), .B1(new_n421), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NOR4_X1   g0266(.A1(new_n361), .A2(new_n420), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT21), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT86), .B(G303), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n255), .A2(new_n259), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G257), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n364), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n217), .A2(G1698), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n287), .A2(new_n257), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n294), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g0277(.A(KEYINPUT5), .B(G41), .Z(new_n478));
  NOR2_X1   g0278(.A1(new_n301), .A2(G1), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(G270), .B(new_n294), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G274), .A3(new_n479), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(G169), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G116), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n280), .A2(new_n281), .B1(G20), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n256), .C1(G33), .C2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n487), .A2(KEYINPUT20), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT20), .B1(new_n487), .B2(new_n490), .ZN(new_n492));
  INV_X1    g0292(.A(new_n320), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n491), .A2(new_n492), .B1(G116), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n322), .A2(G33), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n493), .A2(new_n283), .A3(new_n285), .A4(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n486), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n470), .B1(new_n485), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n477), .A2(new_n484), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n315), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n498), .C1(new_n327), .C2(new_n500), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n472), .A2(new_n476), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n369), .ZN(new_n504));
  INV_X1    g0304(.A(new_n484), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(G179), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT21), .B(G169), .C1(new_n477), .C2(new_n484), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(KEYINPUT87), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT87), .ZN(new_n510));
  AOI211_X1 g0310(.A(new_n510), .B(new_n498), .C1(new_n506), .C2(new_n507), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n499), .B(new_n502), .C1(new_n509), .C2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT85), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n479), .A2(G274), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n294), .A2(new_n480), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n514), .B1(new_n515), .B2(new_n211), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G238), .A2(G1698), .ZN(new_n518));
  INV_X1    g0318(.A(G244), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(G1698), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(new_n287), .A3(new_n257), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n486), .B1(new_n263), .B2(new_n265), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n513), .B(new_n517), .C1(new_n524), .C2(new_n294), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n294), .B1(new_n521), .B2(new_n523), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT85), .B1(new_n526), .B2(new_n516), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n287), .A2(new_n256), .A3(G68), .A4(new_n257), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n256), .B1(new_n367), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(G87), .B2(new_n205), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n386), .B2(new_n489), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n286), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n399), .A2(new_n320), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g0337(.A1(new_n496), .A2(new_n399), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n528), .A2(new_n349), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n525), .A2(new_n345), .A3(new_n527), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n535), .B(new_n536), .C1(new_n210), .C2(new_n496), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n528), .B2(G190), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n525), .A2(G200), .A3(new_n527), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n512), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n211), .A2(new_n364), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n473), .A2(G1698), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n287), .A2(new_n257), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n263), .A2(new_n265), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G294), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n369), .B1(new_n479), .B2(new_n482), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n553), .A2(new_n369), .B1(G264), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n483), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n327), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G190), .B2(new_n556), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n256), .B2(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n216), .A2(KEYINPUT23), .A3(G20), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n522), .A2(new_n256), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n256), .A2(G87), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n287), .A2(new_n565), .A3(new_n257), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n563), .B1(new_n255), .B2(new_n259), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n562), .B(new_n566), .C1(new_n567), .C2(KEYINPUT22), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT88), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n564), .B1(new_n338), .B2(new_n563), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n571), .A2(KEYINPUT88), .A3(new_n562), .A4(new_n566), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n572), .A3(KEYINPUT24), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n568), .A2(new_n569), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n286), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n320), .A2(new_n216), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n577), .B(KEYINPUT25), .ZN(new_n578));
  INV_X1    g0378(.A(new_n496), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(G107), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n558), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(new_n580), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n555), .A2(G179), .A3(new_n483), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n345), .B1(new_n555), .B2(new_n483), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT89), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n556), .A2(G169), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT89), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n583), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n581), .B1(new_n582), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n496), .A2(new_n489), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n320), .A2(new_n489), .ZN(new_n594));
  XOR2_X1   g0394(.A(new_n594), .B(KEYINPUT83), .Z(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n216), .B1(new_n262), .B2(new_n267), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n270), .A2(new_n385), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT6), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n489), .A2(new_n216), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n204), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n216), .A2(KEYINPUT6), .A3(G97), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(new_n256), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n597), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n286), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n593), .B(new_n596), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n287), .A2(G244), .A3(new_n364), .A4(new_n257), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT4), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(KEYINPUT4), .B(new_n364), .C1(new_n336), .C2(new_n337), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(new_n519), .ZN(new_n612));
  OAI211_X1 g0412(.A(G250), .B(G1698), .C1(new_n336), .C2(new_n337), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n488), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n369), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n483), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n554), .B2(G257), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n345), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n607), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n615), .A2(new_n349), .A3(new_n617), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n615), .A2(G190), .A3(new_n617), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n607), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT84), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n615), .A2(KEYINPUT84), .A3(new_n617), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(G200), .A3(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n620), .A2(new_n621), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n469), .A2(new_n547), .A3(new_n591), .A4(new_n629), .ZN(G372));
  INV_X1    g0430(.A(new_n459), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT93), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n355), .B2(new_n352), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n353), .B1(new_n333), .B2(new_n354), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n344), .A2(new_n351), .A3(KEYINPUT18), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(KEYINPUT93), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n395), .ZN(new_n637));
  INV_X1    g0437(.A(new_n416), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n462), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n633), .B(new_n636), .C1(new_n639), .C2(new_n359), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n453), .A2(new_n456), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n631), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n607), .A2(new_n619), .A3(new_n621), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT90), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n526), .A2(new_n646), .ZN(new_n647));
  AOI211_X1 g0447(.A(KEYINPUT90), .B(new_n294), .C1(new_n521), .C2(new_n523), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n517), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n345), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(G200), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n539), .A2(new_n650), .B1(new_n543), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n644), .A2(new_n645), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT26), .B1(new_n546), .B2(new_n643), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n539), .A2(new_n650), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(G107), .B1(new_n339), .B2(new_n340), .ZN(new_n657));
  INV_X1    g0457(.A(new_n598), .ZN(new_n658));
  INV_X1    g0458(.A(new_n604), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AOI211_X1 g0460(.A(new_n592), .B(new_n595), .C1(new_n660), .C2(new_n286), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n628), .A2(new_n622), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n558), .A2(new_n576), .A3(new_n580), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(new_n643), .A4(new_n652), .ZN(new_n664));
  INV_X1    g0464(.A(new_n485), .ZN(new_n665));
  INV_X1    g0465(.A(new_n498), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT21), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT91), .B1(new_n667), .B2(new_n508), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT91), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n506), .A2(new_n507), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n669), .B(new_n499), .C1(new_n670), .C2(new_n498), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n584), .A2(new_n585), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n576), .B2(new_n580), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT92), .B1(new_n664), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n652), .A2(new_n663), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT92), .ZN(new_n679));
  INV_X1    g0479(.A(new_n673), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n582), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n671), .A3(new_n668), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n678), .A2(new_n629), .A3(new_n679), .A4(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n656), .B1(new_n676), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n642), .B1(new_n468), .B2(new_n684), .ZN(G369));
  NOR2_X1   g0485(.A1(new_n319), .A2(G20), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OR3_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .A3(G1), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT27), .B1(new_n687), .B2(G1), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G343), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT94), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n666), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT95), .Z(new_n695));
  NOR2_X1   g0495(.A1(new_n509), .A2(new_n511), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n667), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(new_n697), .A3(new_n502), .ZN(new_n698));
  INV_X1    g0498(.A(new_n672), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n695), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT96), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT96), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G330), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n582), .ZN(new_n704));
  INV_X1    g0504(.A(new_n693), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n591), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n590), .A2(new_n582), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n693), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n705), .B1(new_n696), .B2(new_n667), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n708), .A2(new_n712), .A3(new_n581), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n681), .A2(new_n693), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n224), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G41), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n229), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n719), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT97), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n684), .B2(new_n693), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n697), .A2(new_n707), .ZN(new_n728));
  INV_X1    g0528(.A(new_n627), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT84), .B1(new_n615), .B2(new_n617), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n729), .A2(new_n730), .A3(new_n327), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n592), .B1(new_n660), .B2(new_n286), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n622), .A3(new_n596), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n643), .B(KEYINPUT100), .C1(new_n731), .C2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT100), .B1(new_n662), .B2(new_n643), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n678), .B(new_n728), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n645), .B1(new_n644), .B2(new_n652), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n546), .A2(new_n643), .A3(KEYINPUT26), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n539), .A2(new_n650), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(KEYINPUT29), .A3(new_n705), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n727), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n591), .A2(new_n629), .A3(new_n547), .A4(new_n705), .ZN(new_n745));
  INV_X1    g0545(.A(new_n618), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n506), .B1(new_n525), .B2(new_n527), .ZN(new_n747));
  NOR2_X1   g0547(.A1(KEYINPUT99), .A2(KEYINPUT30), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n294), .B1(new_n550), .B2(new_n552), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n748), .B(new_n749), .C1(G264), .C2(new_n554), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n746), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(KEYINPUT99), .A2(KEYINPUT30), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(G179), .B1(new_n615), .B2(new_n617), .ZN(new_n754));
  INV_X1    g0554(.A(new_n500), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n754), .A2(new_n755), .A3(new_n556), .A4(new_n649), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT99), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT30), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n746), .A2(new_n747), .A3(new_n759), .A4(new_n750), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n753), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n693), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT31), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT98), .B(KEYINPUT31), .Z(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n745), .B(new_n764), .C1(new_n762), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G330), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n744), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n725), .B1(new_n770), .B2(G1), .ZN(G364));
  AOI21_X1  g0571(.A(new_n322), .B1(new_n686), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n718), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n703), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(G330), .B1(new_n701), .B2(new_n702), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n700), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n281), .B1(G20), .B2(new_n345), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n256), .A2(new_n349), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n314), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n784), .A2(new_n327), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G190), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G50), .A2(new_n786), .B1(new_n788), .B2(G77), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n787), .A2(new_n314), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n789), .B1(new_n214), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT102), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G179), .A2(G200), .ZN(new_n794));
  INV_X1    g0594(.A(G190), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n794), .A2(G20), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G159), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT32), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(KEYINPUT32), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n256), .B1(new_n794), .B2(G190), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n489), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n785), .A2(G190), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n219), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n256), .A2(G179), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n806), .A2(G190), .A3(G200), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n210), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n806), .A2(new_n795), .A3(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n216), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n802), .A2(new_n805), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n793), .A2(new_n403), .A3(new_n799), .A4(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT103), .Z(new_n813));
  INV_X1    g0613(.A(new_n801), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n786), .A2(G326), .B1(G294), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n797), .A2(G329), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  INV_X1    g0617(.A(new_n788), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n815), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G322), .B2(new_n790), .ZN(new_n820));
  INV_X1    g0620(.A(new_n807), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G303), .ZN(new_n822));
  NOR2_X1   g0622(.A1(KEYINPUT33), .A2(G317), .ZN(new_n823));
  AND2_X1   g0623(.A1(KEYINPUT33), .A2(G317), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n803), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n820), .A2(new_n338), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n809), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(G283), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n783), .B1(new_n813), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n287), .A2(new_n257), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n224), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT101), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n247), .A2(G45), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(new_n230), .C2(G45), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n403), .A2(G355), .A3(new_n224), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n834), .B(new_n835), .C1(G116), .C2(new_n224), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n780), .A2(new_n783), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n829), .A2(new_n774), .A3(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n776), .A2(new_n777), .B1(new_n782), .B2(new_n839), .ZN(G396));
  INV_X1    g0640(.A(new_n656), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n643), .B1(new_n731), .B2(new_n733), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n677), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n679), .B1(new_n843), .B2(new_n682), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n664), .A2(KEYINPUT92), .A3(new_n675), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n693), .A2(new_n402), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n638), .B1(new_n419), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n416), .A2(new_n693), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n705), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n849), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n419), .A2(new_n847), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(new_n638), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n684), .B2(new_n693), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(G330), .A3(new_n767), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n851), .A2(new_n855), .A3(new_n768), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n775), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n783), .A2(new_n778), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n385), .ZN(new_n861));
  AOI22_X1  g0661(.A1(G150), .A2(new_n803), .B1(new_n788), .B2(G159), .ZN(new_n862));
  INV_X1    g0662(.A(G137), .ZN(new_n863));
  INV_X1    g0663(.A(new_n786), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(G143), .B2(new_n790), .ZN(new_n866));
  XOR2_X1   g0666(.A(KEYINPUT104), .B(KEYINPUT34), .Z(new_n867));
  XNOR2_X1  g0667(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(G132), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n809), .A2(new_n219), .B1(new_n869), .B2(new_n796), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n868), .A2(new_n830), .A3(new_n870), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n871), .B1(new_n430), .B2(new_n807), .C1(new_n214), .C2(new_n801), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n809), .A2(new_n210), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n786), .A2(G303), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n216), .B2(new_n807), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n873), .B(new_n875), .C1(G311), .C2(new_n797), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n803), .A2(G283), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n788), .A2(G116), .B1(G97), .B2(new_n814), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n403), .B1(G294), .B2(new_n790), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n783), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n861), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n850), .A2(new_n779), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n774), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n859), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT105), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(G384));
  OR2_X1    g0690(.A1(new_n289), .A2(new_n290), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT16), .B1(new_n891), .B2(new_n277), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n326), .B1(new_n892), .B2(new_n343), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n690), .B(new_n893), .C1(new_n358), .C2(new_n359), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n344), .B1(new_n351), .B2(new_n690), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n896), .A3(new_n329), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n893), .B1(new_n351), .B2(new_n690), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n898), .A2(new_n329), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n899), .B2(new_n896), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n894), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT39), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n895), .A2(new_n896), .A3(new_n329), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n896), .B1(new_n895), .B2(new_n329), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n335), .A2(new_n633), .A3(new_n636), .ZN(new_n909));
  INV_X1    g0709(.A(new_n690), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n333), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n904), .B(new_n905), .C1(new_n912), .C2(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n903), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n383), .A2(new_n394), .A3(new_n705), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n894), .A2(new_n900), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n905), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n394), .A2(new_n693), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n383), .A2(new_n394), .B1(new_n462), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n684), .A2(new_n854), .A3(new_n693), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n920), .B(new_n923), .C1(new_n924), .C2(new_n849), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n634), .A2(KEYINPUT93), .A3(new_n635), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT93), .B1(new_n634), .B2(new_n635), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n910), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n916), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n727), .B(new_n743), .C1(new_n465), .C2(new_n467), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n642), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n762), .A2(new_n766), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n761), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n745), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n935), .A2(new_n923), .A3(new_n850), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT40), .B1(new_n936), .B2(new_n920), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n905), .B1(new_n912), .B2(KEYINPUT38), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT107), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT107), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n940), .B(new_n905), .C1(new_n912), .C2(KEYINPUT38), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n935), .A2(new_n923), .A3(KEYINPUT40), .A4(new_n850), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n937), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n469), .A3(new_n935), .ZN(new_n946));
  OAI211_X1 g0746(.A(G330), .B(new_n935), .C1(new_n465), .C2(new_n467), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n943), .B1(new_n939), .B2(new_n941), .ZN(new_n949));
  INV_X1    g0749(.A(G330), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n949), .A2(new_n950), .A3(new_n937), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n946), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n932), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n322), .B2(new_n686), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n229), .A2(G77), .A3(new_n275), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(G50), .B2(new_n219), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(G1), .A3(new_n319), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT35), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n227), .B1(new_n603), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n959), .B(G116), .C1(new_n958), .C2(new_n603), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT106), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT36), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n954), .A2(new_n957), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT108), .ZN(G367));
  INV_X1    g0764(.A(KEYINPUT44), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n735), .A2(new_n736), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n607), .A2(new_n693), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n966), .A2(new_n967), .B1(new_n644), .B2(new_n693), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n965), .B1(new_n969), .B2(new_n715), .ZN(new_n970));
  INV_X1    g0770(.A(new_n715), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(new_n971), .A3(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n969), .A2(KEYINPUT45), .A3(new_n715), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n968), .B2(new_n971), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n703), .A2(new_n710), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT110), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n970), .A2(new_n972), .B1(new_n974), .B2(new_n976), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(KEYINPUT111), .A3(new_n711), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT111), .B1(new_n982), .B2(new_n711), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n713), .B1(new_n710), .B2(new_n712), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n703), .B(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n770), .B(new_n988), .C1(new_n980), .C2(KEYINPUT110), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n770), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n718), .B(KEYINPUT41), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n773), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n966), .A2(new_n708), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n705), .B1(new_n993), .B2(new_n644), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n966), .A2(new_n713), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(KEYINPUT42), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n995), .A2(KEYINPUT42), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n693), .A2(new_n542), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n655), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n652), .B2(new_n999), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n998), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT109), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(KEYINPUT109), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n1003), .C2(new_n998), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n711), .A2(new_n968), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1008), .B(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1001), .A2(new_n780), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n832), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n837), .B1(new_n224), .B2(new_n399), .C1(new_n1013), .C2(new_n239), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n809), .A2(new_n385), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n803), .A2(G159), .B1(new_n821), .B2(G58), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n423), .B2(new_n791), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(G137), .C2(new_n797), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n786), .A2(G143), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n801), .A2(new_n219), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n788), .B2(G50), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n403), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n864), .A2(new_n817), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G283), .A2(new_n788), .B1(new_n790), .B2(new_n471), .ZN(new_n1024));
  INV_X1    g0824(.A(G294), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n830), .C1(new_n1025), .C2(new_n804), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n807), .A2(new_n486), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT46), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n801), .A2(new_n216), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n797), .A2(G317), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n827), .A2(G97), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1022), .B1(new_n1023), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT47), .Z(new_n1035));
  OAI211_X1 g0835(.A(new_n774), .B(new_n1014), .C1(new_n1035), .C2(new_n882), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n992), .A2(new_n1011), .B1(new_n1012), .B2(new_n1036), .ZN(G387));
  NAND2_X1  g0837(.A1(new_n988), .A2(new_n773), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT112), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n988), .A2(new_n770), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n988), .A2(new_n770), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n718), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n710), .A2(new_n780), .ZN(new_n1043));
  AOI21_X1  g0843(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n318), .A2(new_n430), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n720), .B(new_n1044), .C1(new_n1045), .C2(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(KEYINPUT50), .B2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n832), .B1(new_n236), .B2(new_n301), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n338), .A2(new_n717), .A3(new_n720), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n216), .B2(new_n717), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n837), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n774), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT113), .Z(new_n1054));
  NAND2_X1  g0854(.A1(new_n786), .A2(G159), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n803), .A2(new_n318), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n821), .A2(G77), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1032), .A4(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n818), .A2(new_n219), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n791), .A2(new_n430), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n796), .A2(new_n423), .ZN(new_n1061));
  NOR4_X1   g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n801), .A2(new_n399), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1062), .A2(new_n257), .A3(new_n287), .A4(new_n1063), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT114), .Z(new_n1065));
  AOI22_X1  g0865(.A1(G317), .A2(new_n790), .B1(new_n788), .B2(new_n471), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT115), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n817), .B2(new_n804), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G322), .B2(new_n786), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT48), .Z(new_n1070));
  INV_X1    g0870(.A(G283), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n801), .C1(new_n1025), .C2(new_n807), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT49), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n827), .A2(G116), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n797), .A2(G326), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1074), .A2(new_n830), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1065), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1043), .B(new_n1054), .C1(new_n1077), .C2(new_n882), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1039), .A2(new_n1042), .A3(new_n1078), .ZN(G393));
  INV_X1    g0879(.A(KEYINPUT116), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n984), .B2(new_n985), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT111), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n978), .B2(new_n979), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(KEYINPUT116), .A3(new_n983), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1081), .A2(new_n1084), .A3(new_n980), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1041), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n986), .A2(new_n989), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n1087), .A3(new_n718), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1081), .A2(new_n1084), .A3(new_n773), .A4(new_n980), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n968), .A2(new_n780), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT117), .Z(new_n1091));
  AOI22_X1  g0891(.A1(G311), .A2(new_n790), .B1(new_n786), .B2(G317), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT52), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n810), .B(new_n1093), .C1(new_n471), .C2(new_n803), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n821), .A2(G283), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n814), .A2(G116), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n818), .A2(new_n1025), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n403), .B(new_n1097), .C1(G322), .C2(new_n797), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G150), .A2(new_n786), .B1(new_n790), .B2(G159), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT51), .Z(new_n1101));
  NAND2_X1  g0901(.A1(new_n803), .A2(G50), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n830), .B(new_n873), .C1(G143), .C2(new_n797), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n801), .A2(new_n385), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n807), .A2(new_n219), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(new_n318), .C2(new_n788), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n882), .B1(new_n1099), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n837), .B1(new_n489), .B2(new_n224), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n244), .B2(new_n832), .ZN(new_n1110));
  OR4_X1    g0910(.A1(new_n775), .A2(new_n1091), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1089), .A2(KEYINPUT118), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT118), .B1(new_n1089), .B2(new_n1111), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1088), .B1(new_n1112), .B2(new_n1113), .ZN(G390));
  INV_X1    g0914(.A(new_n914), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n923), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n851), .B2(new_n852), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1117), .B2(new_n915), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n922), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n693), .B(new_n848), .C1(new_n737), .C2(new_n741), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n849), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n915), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n942), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n935), .A2(new_n923), .A3(G330), .A4(new_n850), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n767), .A2(new_n923), .A3(G330), .A4(new_n850), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1118), .A2(new_n1128), .A3(new_n1123), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n773), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n775), .B1(new_n1115), .B2(new_n778), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n860), .A2(new_n317), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n814), .A2(G159), .B1(new_n797), .B2(G125), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT54), .B(G143), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1133), .B(new_n403), .C1(new_n818), .C2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n807), .A2(new_n423), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n790), .A2(G132), .B1(new_n827), .B2(G50), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(new_n863), .C2(new_n804), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1135), .B(new_n1139), .C1(G128), .C2(new_n786), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n790), .A2(G116), .B1(new_n827), .B2(G68), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1141), .B1(new_n216), .B2(new_n804), .C1(new_n1025), .C2(new_n796), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n338), .B1(new_n818), .B2(new_n489), .C1(new_n1071), .C2(new_n864), .ZN(new_n1143));
  NOR4_X1   g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n808), .A4(new_n1104), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n783), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1131), .A2(new_n1132), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1130), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1118), .A2(new_n1128), .A3(new_n1123), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1125), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n851), .A2(new_n852), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1116), .B1(new_n768), .B2(new_n854), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1125), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n935), .A2(G330), .A3(new_n850), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n1116), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1155), .A2(new_n1128), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1120), .A2(new_n849), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1151), .A2(new_n1153), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n947), .A2(new_n930), .A3(new_n642), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n719), .B1(new_n1150), .B2(new_n1160), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1147), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(G378));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n908), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n926), .A2(new_n927), .A3(new_n359), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n911), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n918), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n940), .B1(new_n1171), .B2(new_n905), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n941), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n944), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n937), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(G330), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n929), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n453), .A2(new_n456), .A3(new_n459), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT119), .Z(new_n1181));
  AOI21_X1  g0981(.A(new_n910), .B1(new_n431), .B2(new_n432), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1179), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1178), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n916), .A2(new_n925), .A3(new_n928), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n945), .A3(G330), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1177), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1190), .B1(new_n1177), .B2(new_n1192), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT121), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1159), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n947), .A2(new_n930), .A3(KEYINPUT121), .A4(new_n642), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1150), .B2(new_n1160), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1166), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n929), .A2(new_n1176), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n951), .A2(new_n1191), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1189), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1177), .A2(new_n1192), .A3(new_n1190), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1160), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1209), .A3(KEYINPUT57), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1201), .A2(new_n718), .A3(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1185), .A2(new_n1188), .A3(new_n778), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n830), .B1(new_n214), .B2(new_n809), .C1(new_n791), .C2(new_n216), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1020), .B(new_n1213), .C1(G116), .C2(new_n786), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n803), .A2(G97), .B1(G283), .B2(new_n797), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1215), .A2(new_n293), .A3(new_n1057), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(new_n399), .C2(new_n818), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT58), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n804), .A2(new_n869), .B1(new_n807), .B2(new_n1134), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G150), .B2(new_n814), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G125), .A2(new_n786), .B1(new_n788), .B2(G137), .ZN(new_n1221));
  INV_X1    g1021(.A(G128), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1220), .B(new_n1221), .C1(new_n1222), .C2(new_n791), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT59), .Z(new_n1224));
  OAI21_X1  g1024(.A(new_n293), .B1(new_n809), .B2(new_n271), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G124), .B2(new_n797), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n251), .A3(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n293), .B1(new_n265), .B2(new_n253), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n430), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1218), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n783), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n860), .A2(new_n430), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1212), .A2(new_n774), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT120), .Z(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1206), .B2(new_n773), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1211), .A2(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1236), .A2(KEYINPUT122), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(KEYINPUT122), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(G375));
  INV_X1    g1039(.A(new_n1158), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1063), .B1(new_n791), .B2(new_n1071), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT124), .Z(new_n1242));
  AOI211_X1 g1042(.A(new_n1015), .B(new_n1242), .C1(G294), .C2(new_n786), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n821), .A2(G97), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n403), .B1(G303), .B2(new_n797), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G107), .A2(new_n788), .B1(new_n803), .B2(G116), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n796), .A2(new_n1222), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n791), .A2(new_n863), .B1(new_n271), .B2(new_n807), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(G132), .C2(new_n786), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n809), .A2(new_n214), .B1(new_n801), .B2(new_n430), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n830), .B(new_n1251), .C1(G150), .C2(new_n788), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1250), .B(new_n1252), .C1(new_n804), .C2(new_n1134), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n882), .B1(new_n1247), .B2(new_n1253), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n775), .B(new_n1254), .C1(new_n219), .C2(new_n860), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1116), .A2(new_n778), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT123), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1240), .A2(new_n773), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n991), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1260), .B2(new_n1160), .ZN(G381));
  NAND3_X1  g1061(.A1(new_n1237), .A2(new_n1164), .A3(new_n1238), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(G384), .A2(G381), .ZN(new_n1264));
  OR2_X1    g1064(.A1(G390), .A2(G387), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1265), .A2(G396), .A3(G393), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .ZN(G407));
  OAI211_X1 g1067(.A(G407), .B(G213), .C1(G343), .C2(new_n1262), .ZN(G409));
  NAND2_X1  g1068(.A1(new_n1236), .A2(G378), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT125), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT125), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1204), .A2(new_n1271), .A3(new_n1205), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1272), .A3(new_n773), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1206), .A2(new_n1209), .A3(new_n991), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1233), .B(KEYINPUT120), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1273), .A2(new_n1164), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(G343), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(G213), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1259), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1158), .A2(new_n1159), .A3(KEYINPUT60), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1162), .A3(new_n718), .A4(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1258), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n889), .B2(new_n888), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G384), .A2(new_n1258), .A3(new_n1283), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1269), .A2(new_n1279), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT62), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1277), .A2(G213), .A3(G2897), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1291), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1164), .B1(new_n1211), .B2(new_n1235), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1292), .B(new_n1295), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT62), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1269), .A2(new_n1279), .A3(new_n1287), .A4(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1289), .A2(new_n1290), .A3(new_n1298), .A4(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G390), .B(G387), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(G393), .B(G396), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G390), .A2(G387), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1265), .A2(new_n1305), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1298), .A2(new_n1290), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1311), .A2(new_n1289), .A3(KEYINPUT126), .A4(new_n1300), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1303), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1298), .A2(KEYINPUT63), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT61), .B1(new_n1315), .B2(new_n1288), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1314), .B(new_n1316), .C1(new_n1317), .C2(new_n1288), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1313), .A2(new_n1318), .ZN(G405));
  AOI21_X1  g1119(.A(new_n1293), .B1(new_n1262), .B2(new_n1269), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1262), .A2(new_n1269), .A3(new_n1293), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1314), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1262), .A2(new_n1269), .A3(new_n1293), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1324), .A2(new_n1320), .A3(new_n1310), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1323), .A2(new_n1325), .ZN(G402));
endmodule


