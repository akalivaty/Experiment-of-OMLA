//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT38), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT29), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n212));
  AOI21_X1  g011(.A(G183gat), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g017(.A(KEYINPUT25), .B(new_n210), .C1(new_n213), .C2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT23), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT65), .A4(KEYINPUT23), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n210), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n216), .B(new_n217), .C1(G183gat), .C2(G190gat), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n224), .A2(new_n210), .A3(KEYINPUT66), .A4(new_n225), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n232));
  AOI21_X1  g031(.A(new_n222), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n212), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT28), .ZN(new_n235));
  NOR2_X1   g034(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n234), .B(new_n235), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT67), .B(G190gat), .Z(new_n240));
  INV_X1    g039(.A(new_n236), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(KEYINPUT68), .A3(new_n237), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(new_n238), .B2(new_n236), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n240), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n214), .B(new_n239), .C1(new_n245), .C2(new_n235), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n209), .A2(KEYINPUT26), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n209), .A2(KEYINPUT26), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n247), .A2(new_n205), .A3(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n204), .B1(new_n233), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n233), .B2(new_n250), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT74), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT74), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n257), .B(new_n254), .C1(new_n233), .C2(new_n250), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G197gat), .B(G204gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT22), .ZN(new_n261));
  INV_X1    g060(.A(G211gat), .ZN(new_n262));
  INV_X1    g061(.A(G218gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n260), .A3(new_n264), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n255), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n271), .B(KEYINPUT37), .C1(new_n270), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n270), .ZN(new_n274));
  INV_X1    g073(.A(new_n270), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n253), .A2(new_n256), .A3(new_n275), .A4(new_n258), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT37), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G8gat), .B(G36gat), .Z(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(G64gat), .ZN(new_n281));
  INV_X1    g080(.A(G92gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  AND4_X1   g082(.A1(new_n203), .A2(new_n273), .A3(new_n279), .A4(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n285));
  AND2_X1   g084(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n287));
  OAI21_X1  g086(.A(G141gat), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G141gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G148gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n288), .A2(new_n290), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G155gat), .B(G162gat), .ZN(new_n296));
  INV_X1    g095(.A(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G141gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n296), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT3), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302));
  INV_X1    g101(.A(new_n291), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(new_n292), .ZN(new_n304));
  XNOR2_X1  g103(.A(G141gat), .B(G148gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(KEYINPUT2), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n297), .A2(G141gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT76), .B(G148gat), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(G141gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n291), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n302), .B(new_n306), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n314));
  INV_X1    g113(.A(G134gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G127gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n314), .B(new_n318), .C1(new_n319), .C2(new_n317), .ZN(new_n320));
  INV_X1    g119(.A(G120gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G113gat), .ZN(new_n322));
  INV_X1    g121(.A(G113gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G120gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n315), .A2(G127gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n317), .A2(new_n314), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT71), .B(G113gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n322), .B1(new_n330), .B2(new_n321), .ZN(new_n331));
  INV_X1    g130(.A(G127gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(G134gat), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n333), .A2(new_n327), .A3(KEYINPUT1), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n320), .A2(new_n329), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n285), .B1(new_n313), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n335), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n337), .A2(KEYINPUT77), .A3(new_n301), .A4(new_n312), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n288), .A2(new_n290), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n289), .A2(G148gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n293), .B1(new_n307), .B2(new_n342), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n341), .A2(new_n310), .B1(new_n343), .B2(new_n304), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n320), .A2(new_n329), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n331), .A2(new_n334), .ZN(new_n346));
  AND4_X1   g145(.A1(KEYINPUT4), .A2(new_n344), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT4), .B1(new_n335), .B2(new_n344), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(KEYINPUT5), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n339), .A2(new_n340), .A3(new_n349), .A4(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n349), .A2(new_n336), .A3(new_n338), .A4(new_n352), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT79), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n344), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n351), .B1(new_n337), .B2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n349), .A2(new_n336), .A3(new_n338), .A4(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n335), .B(new_n344), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(new_n351), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G1gat), .B(G29gat), .Z(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G57gat), .B(G85gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n364), .A2(KEYINPUT6), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n283), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n277), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n369), .A3(new_n363), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n353), .A2(new_n355), .B1(new_n359), .B2(new_n362), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(new_n369), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n371), .B(new_n373), .C1(new_n376), .C2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n202), .B1(new_n284), .B2(new_n379), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n377), .A2(new_n375), .A3(new_n369), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n370), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT6), .B1(new_n377), .B2(new_n369), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n273), .A2(new_n279), .A3(new_n203), .A4(new_n283), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n384), .A2(KEYINPUT86), .A3(new_n373), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n274), .A2(KEYINPUT37), .A3(new_n276), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT87), .A3(new_n283), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n279), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT87), .B1(new_n387), .B2(new_n283), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT38), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n380), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n274), .A2(new_n276), .A3(new_n283), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT30), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n373), .ZN(new_n395));
  INV_X1    g194(.A(new_n276), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n275), .B1(new_n253), .B2(new_n255), .ZN(new_n397));
  OAI211_X1 g196(.A(KEYINPUT30), .B(new_n372), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT75), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT75), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n277), .A2(new_n400), .A3(KEYINPUT30), .A4(new_n372), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n349), .A2(new_n336), .A3(new_n338), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n351), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n404), .A2(KEYINPUT39), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n404), .B(KEYINPUT39), .C1(new_n351), .C2(new_n361), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n369), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(KEYINPUT40), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n408), .A3(new_n382), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT85), .ZN(new_n410));
  XOR2_X1   g209(.A(G78gat), .B(G106gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT31), .ZN(new_n412));
  INV_X1    g211(.A(G50gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT29), .B1(new_n268), .B2(new_n269), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n357), .B1(new_n415), .B2(KEYINPUT3), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT29), .B1(new_n344), .B2(new_n302), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n416), .B1(new_n417), .B2(new_n270), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT82), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n417), .B2(new_n270), .ZN(new_n420));
  INV_X1    g219(.A(G228gat), .ZN(new_n421));
  INV_X1    g220(.A(G233gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n418), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  OAI221_X1 g224(.A(new_n416), .B1(new_n419), .B2(new_n423), .C1(new_n417), .C2(new_n270), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G22gat), .ZN(new_n428));
  INV_X1    g227(.A(G22gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n425), .A2(new_n429), .A3(new_n426), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n414), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n425), .B2(new_n426), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n432), .A2(KEYINPUT83), .ZN(new_n433));
  INV_X1    g232(.A(new_n414), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n432), .B2(KEYINPUT83), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n435), .A3(new_n430), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT84), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n433), .A2(new_n435), .A3(new_n438), .A4(new_n430), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n431), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n402), .A2(new_n408), .A3(new_n442), .A4(new_n382), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n392), .A2(new_n410), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT80), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n382), .B1(new_n383), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n374), .A2(new_n446), .A3(new_n375), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n445), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n376), .A2(KEYINPUT80), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(KEYINPUT81), .A3(new_n382), .A4(new_n448), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n371), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n402), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n440), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n233), .A2(new_n250), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n335), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n337), .B1(new_n233), .B2(new_n250), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G227gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n422), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT34), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n464));
  INV_X1    g263(.A(new_n462), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n458), .A2(new_n464), .A3(new_n465), .A4(new_n459), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G71gat), .B(G99gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT72), .ZN(new_n469));
  XNOR2_X1  g268(.A(G15gat), .B(G43gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n460), .A2(new_n462), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT33), .B1(new_n460), .B2(new_n462), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n463), .B(new_n466), .C1(new_n476), .C2(new_n471), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n479), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(new_n481), .A3(new_n477), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT73), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT36), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n475), .A2(new_n481), .A3(new_n477), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n481), .B1(new_n475), .B2(new_n477), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n484), .B(KEYINPUT36), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n444), .A2(new_n456), .A3(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n440), .A2(new_n486), .A3(new_n487), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n453), .A2(new_n492), .A3(new_n454), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT35), .ZN(new_n494));
  OR3_X1    g293(.A1(new_n402), .A2(new_n384), .A3(KEYINPUT88), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT88), .B1(new_n402), .B2(new_n384), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n492), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n491), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT16), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(G1gat), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(G1gat), .B2(new_n504), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(G8gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(G8gat), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT21), .ZN(new_n511));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G71gat), .B(G78gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n510), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G183gat), .ZN(new_n519));
  AND2_X1   g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G127gat), .B(G155gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(new_n262), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n521), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n517), .A2(new_n511), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n525), .B(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G29gat), .ZN(new_n530));
  INV_X1    g329(.A(G36gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT14), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(G29gat), .B2(G36gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT15), .ZN(new_n536));
  XOR2_X1   g335(.A(G43gat), .B(G50gat), .Z(new_n537));
  AOI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G29gat), .A2(G36gat), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n538), .B(new_n539), .C1(new_n536), .C2(new_n537), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n537), .A2(new_n536), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n535), .A2(KEYINPUT91), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n539), .B1(new_n535), .B2(KEYINPUT91), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT17), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  INV_X1    g346(.A(G85gat), .ZN(new_n548));
  AOI22_X1  g347(.A1(KEYINPUT8), .A2(new_n547), .B1(new_n548), .B2(new_n282), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT95), .ZN(new_n550));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT7), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G99gat), .B(G106gat), .Z(new_n554));
  OR2_X1    g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n546), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n556), .A3(new_n545), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT96), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n563), .B(new_n568), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n529), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n508), .A2(new_n509), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT92), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(KEYINPUT92), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n546), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT93), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n545), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT94), .Z(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT93), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n546), .A2(new_n574), .A3(new_n580), .A4(new_n573), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n576), .A2(new_n578), .A3(new_n579), .A4(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT18), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n572), .A2(new_n545), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n579), .B(KEYINPUT13), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n583), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(G169gat), .B(G197gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT12), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n584), .A2(new_n588), .A3(new_n589), .A4(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G230gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(new_n422), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n557), .A2(new_n517), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n555), .A2(new_n556), .A3(new_n516), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n605), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n606), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n603), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n208), .ZN(new_n615));
  INV_X1    g414(.A(G204gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n610), .A2(new_n612), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n601), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n571), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n501), .A2(new_n503), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n501), .A2(KEYINPUT97), .A3(new_n503), .A4(new_n624), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n453), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g431(.A(KEYINPUT16), .B(G8gat), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n491), .A2(new_n499), .A3(new_n502), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n502), .B1(new_n491), .B2(new_n499), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT97), .B1(new_n636), .B2(new_n624), .ZN(new_n637));
  INV_X1    g436(.A(new_n628), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n402), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n629), .A2(KEYINPUT98), .A3(new_n402), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n633), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT99), .B1(new_n643), .B2(KEYINPUT42), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n639), .A2(new_n645), .A3(new_n633), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT98), .B1(new_n629), .B2(new_n402), .ZN(new_n647));
  AOI211_X1 g446(.A(new_n640), .B(new_n454), .C1(new_n627), .C2(new_n628), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n646), .B1(new_n649), .B2(G8gat), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n651), .B(new_n645), .C1(new_n649), .C2(new_n633), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n644), .A2(new_n650), .A3(new_n652), .ZN(G1325gat));
  INV_X1    g452(.A(new_n483), .ZN(new_n654));
  AOI21_X1  g453(.A(G15gat), .B1(new_n629), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n483), .A2(new_n484), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT36), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n488), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT100), .B1(new_n485), .B2(new_n489), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n627), .B2(new_n628), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n655), .B1(new_n663), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g463(.A1(new_n629), .A2(new_n440), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT43), .B(G22gat), .Z(new_n666));
  AND2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n667), .B2(new_n668), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(G1327gat));
  NAND4_X1  g472(.A1(new_n636), .A2(new_n570), .A3(new_n529), .A4(new_n623), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n530), .A3(new_n630), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT45), .ZN(new_n677));
  INV_X1    g476(.A(new_n662), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n444), .A2(new_n456), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n499), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n680), .A2(new_n681), .A3(new_n570), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n501), .A2(new_n503), .A3(new_n570), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(KEYINPUT44), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n623), .A2(new_n529), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT103), .Z(new_n686));
  NOR3_X1   g485(.A1(new_n684), .A2(new_n453), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n677), .B1(new_n687), .B2(new_n530), .ZN(G1328gat));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n674), .A2(G36gat), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(new_n402), .ZN(new_n691));
  NOR4_X1   g490(.A1(new_n674), .A2(KEYINPUT104), .A3(G36gat), .A4(new_n454), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT46), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR3_X1    g494(.A1(new_n691), .A2(KEYINPUT46), .A3(new_n692), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n683), .A2(KEYINPUT44), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n681), .A3(new_n570), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n686), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n402), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G36gat), .ZN(new_n702));
  OAI211_X1 g501(.A(KEYINPUT105), .B(KEYINPUT46), .C1(new_n691), .C2(new_n692), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n695), .A2(new_n696), .A3(new_n702), .A4(new_n703), .ZN(G1329gat));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n684), .A2(new_n662), .A3(new_n686), .ZN(new_n706));
  INV_X1    g505(.A(G43gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n675), .A2(new_n707), .A3(new_n654), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n706), .B2(new_n707), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI221_X1 g511(.A(new_n709), .B1(new_n705), .B2(KEYINPUT47), .C1(new_n706), .C2(new_n707), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1330gat));
  OAI21_X1  g513(.A(new_n413), .B1(new_n674), .B2(new_n441), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n699), .A2(G50gat), .A3(new_n700), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(new_n441), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g517(.A1(new_n680), .A2(new_n622), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n571), .A2(new_n601), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n630), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n722), .A2(new_n402), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n726), .B(new_n727), .Z(G1333gat));
  NAND3_X1  g527(.A1(new_n722), .A2(G71gat), .A3(new_n678), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n722), .A2(new_n654), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(G71gat), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n722), .A2(new_n440), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g533(.A1(new_n529), .A2(new_n601), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n622), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT108), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n740), .A3(new_n622), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n697), .B2(new_n698), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n630), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(KEYINPUT109), .A3(new_n630), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(G85gat), .A3(new_n747), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n680), .A2(new_n570), .A3(new_n737), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n680), .A2(new_n570), .A3(new_n737), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT51), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(new_n622), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n548), .A3(new_n630), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n748), .A2(new_n756), .ZN(G1336gat));
  NAND2_X1  g556(.A1(new_n750), .A2(KEYINPUT110), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n749), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n454), .A2(G92gat), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n759), .A2(new_n622), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n282), .B1(new_n743), .B2(new_n402), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT52), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND4_X1   g562(.A1(new_n622), .A2(new_n751), .A3(new_n753), .A4(new_n760), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765));
  NOR4_X1   g564(.A1(new_n762), .A2(new_n764), .A3(new_n765), .A4(KEYINPUT52), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n739), .A2(new_n741), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n699), .A2(new_n402), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(new_n768), .B2(G92gat), .ZN(new_n769));
  INV_X1    g568(.A(new_n764), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT111), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n763), .B1(new_n766), .B2(new_n771), .ZN(G1337gat));
  INV_X1    g571(.A(G99gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n773), .A3(new_n654), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n684), .A2(new_n662), .A3(new_n742), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(G1338gat));
  NOR2_X1   g575(.A1(KEYINPUT112), .A2(G106gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n743), .B2(new_n440), .ZN(new_n778));
  NAND2_X1  g577(.A1(KEYINPUT112), .A2(G106gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n441), .A2(G106gat), .A3(new_n621), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT53), .B1(new_n754), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n778), .A2(new_n779), .B1(new_n759), .B2(new_n781), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(G1339gat));
  NAND3_X1  g585(.A1(new_n607), .A2(new_n608), .A3(new_n603), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n610), .A2(KEYINPUT54), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n609), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT113), .B1(new_n790), .B2(new_n617), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n792), .B(new_n619), .C1(new_n609), .C2(new_n789), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n788), .B(KEYINPUT55), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n620), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n788), .B1(new_n791), .B2(new_n793), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n797), .A2(KEYINPUT114), .A3(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n578), .A2(new_n585), .A3(new_n587), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n578), .A2(new_n805), .A3(new_n585), .A4(new_n587), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n576), .A2(new_n581), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n579), .B1(new_n808), .B2(new_n578), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n595), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n599), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n801), .A3(new_n802), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n811), .B1(new_n599), .B2(new_n810), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n813), .A2(new_n569), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n796), .A2(new_n801), .A3(new_n600), .A4(new_n802), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n622), .A2(new_n599), .A3(new_n810), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n570), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n529), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n571), .A2(new_n601), .A3(new_n621), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(new_n492), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n453), .A2(new_n402), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n600), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G113gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n330), .B2(new_n824), .ZN(G1340gat));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n823), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n621), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(new_n321), .ZN(G1341gat));
  NOR2_X1   g628(.A1(new_n827), .A2(new_n529), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT117), .B(G127gat), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n830), .B(new_n831), .ZN(G1342gat));
  NOR2_X1   g631(.A1(new_n827), .A2(new_n569), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI22_X1  g635(.A1(new_n836), .A2(G134gat), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n315), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n837), .B(new_n838), .C1(new_n315), .C2(new_n833), .ZN(G1343gat));
  NAND2_X1  g638(.A1(new_n662), .A2(new_n823), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n797), .A2(new_n798), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n795), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n799), .A2(KEYINPUT119), .A3(new_n620), .A4(new_n794), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n600), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n570), .B1(new_n847), .B2(new_n817), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n529), .B1(new_n848), .B2(new_n815), .ZN(new_n849));
  AOI211_X1 g648(.A(new_n842), .B(new_n441), .C1(new_n849), .C2(new_n820), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT57), .B1(new_n821), .B2(new_n440), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n841), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G141gat), .B1(new_n852), .B2(new_n601), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n441), .B1(new_n819), .B2(new_n820), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n841), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n289), .A3(new_n600), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n308), .A3(new_n622), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n622), .B(new_n841), .C1(new_n850), .C2(new_n851), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  INV_X1    g661(.A(new_n308), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n821), .A2(new_n440), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT57), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n820), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n571), .A2(KEYINPUT120), .A3(new_n601), .A4(new_n621), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n849), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n842), .A3(new_n440), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n866), .A2(new_n871), .A3(new_n622), .A4(new_n841), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n862), .B1(new_n872), .B2(G148gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n860), .B1(new_n864), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(KEYINPUT121), .B(new_n860), .C1(new_n864), .C2(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1345gat));
  INV_X1    g677(.A(G155gat), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n852), .A2(new_n879), .A3(new_n529), .ZN(new_n880));
  INV_X1    g679(.A(new_n529), .ZN(new_n881));
  AOI21_X1  g680(.A(G155gat), .B1(new_n856), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(G1346gat));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n852), .A2(new_n569), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G162gat), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n855), .A2(G162gat), .A3(new_n569), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n884), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT122), .B(new_n887), .C1(new_n885), .C2(G162gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n630), .A2(new_n454), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n821), .A2(new_n492), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n601), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(new_n207), .ZN(G1348gat));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n621), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(new_n208), .ZN(G1349gat));
  NAND2_X1  g696(.A1(new_n242), .A2(new_n244), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n822), .A2(new_n898), .A3(new_n881), .A4(new_n892), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  OAI21_X1  g699(.A(G183gat), .B1(new_n893), .B2(new_n529), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT124), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n902), .B(new_n904), .C1(new_n900), .C2(new_n899), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n903), .A2(KEYINPUT124), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n905), .B(new_n906), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n822), .A2(new_n570), .A3(new_n892), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(G190gat), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n909), .A2(KEYINPUT61), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(KEYINPUT61), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n910), .B(new_n911), .C1(new_n240), .C2(new_n908), .ZN(G1351gat));
  XNOR2_X1  g711(.A(KEYINPUT125), .B(G197gat), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n866), .A2(new_n871), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n662), .A2(new_n892), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n916), .B2(new_n601), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n854), .A2(new_n915), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n601), .A2(new_n913), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(G1352gat));
  NAND3_X1  g719(.A1(new_n914), .A2(new_n622), .A3(new_n915), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT127), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n914), .A2(new_n923), .A3(new_n622), .A4(new_n915), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n922), .A2(G204gat), .A3(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n918), .A2(G204gat), .A3(new_n621), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930));
  OR3_X1    g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n928), .B2(new_n929), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n925), .A2(new_n931), .A3(new_n932), .ZN(G1353gat));
  INV_X1    g732(.A(new_n918), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n262), .A3(new_n881), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n914), .A2(new_n881), .A3(new_n915), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  OAI21_X1  g738(.A(G218gat), .B1(new_n916), .B2(new_n569), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n263), .A3(new_n570), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1355gat));
endmodule


