//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n204));
  NAND2_X1  g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT83), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT83), .A2(G29gat), .A3(G36gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n204), .A2(new_n207), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G43gat), .ZN(new_n213));
  INV_X1    g012(.A(G43gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G50gat), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT15), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT15), .B1(new_n213), .B2(new_n215), .ZN(new_n217));
  NOR3_X1   g016(.A1(new_n211), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n204), .A2(new_n209), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n219), .B1(new_n221), .B2(new_n205), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT17), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n217), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n207), .A2(new_n210), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n224), .A2(new_n221), .A3(new_n219), .A4(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n227));
  INV_X1    g026(.A(new_n205), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n216), .B1(new_n220), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT85), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(G1gat), .ZN(new_n234));
  INV_X1    g033(.A(G8gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(G1gat), .B1(new_n233), .B2(KEYINPUT84), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT16), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G22gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G15gat), .ZN(new_n242));
  INV_X1    g041(.A(G15gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G22gat), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n242), .A2(new_n244), .A3(KEYINPUT84), .A4(G1gat), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n236), .A2(new_n238), .A3(new_n240), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n245), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n235), .B(new_n234), .C1(new_n247), .C2(new_n237), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G229gat), .A2(G233gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n226), .A2(new_n229), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n252), .A3(new_n248), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT18), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n250), .A2(KEYINPUT18), .A3(new_n251), .A4(new_n253), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n251), .B(KEYINPUT13), .Z(new_n258));
  INV_X1    g057(.A(new_n253), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n252), .B1(new_n246), .B2(new_n248), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n256), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G113gat), .B(G141gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G169gat), .B(G197gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT12), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n256), .A2(new_n257), .A3(new_n261), .A4(new_n268), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT28), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT27), .B(G183gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n278), .B2(G190gat), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n277), .B(new_n280), .C1(new_n275), .C2(KEYINPUT28), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n279), .A2(new_n281), .B1(G183gat), .B2(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT65), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT26), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  OAI22_X1  g087(.A1(new_n288), .A2(KEYINPUT69), .B1(KEYINPUT26), .B2(new_n286), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n282), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n285), .B(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n293), .A2(new_n284), .ZN(new_n294));
  NOR2_X1   g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT66), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n295), .A2(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT67), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n297), .A2(new_n301), .A3(new_n305), .A4(new_n302), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n294), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT25), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT25), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n302), .A2(new_n310), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n299), .A2(new_n300), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(new_n313), .A3(new_n296), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n294), .B(new_n309), .C1(new_n311), .C2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n291), .A2(new_n308), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G113gat), .B2(G120gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n318), .B1(G113gat), .B2(G120gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(G127gat), .B(G134gat), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI22_X1  g120(.A1(KEYINPUT71), .A2(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(KEYINPUT71), .B2(KEYINPUT1), .ZN(new_n323));
  INV_X1    g122(.A(G113gat), .ZN(new_n324));
  XOR2_X1   g123(.A(KEYINPUT70), .B(G120gat), .Z(new_n325));
  OAI211_X1 g124(.A(new_n323), .B(new_n320), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n274), .B1(new_n316), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n308), .A2(new_n315), .ZN(new_n329));
  INV_X1    g128(.A(new_n327), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n329), .A2(KEYINPUT72), .A3(new_n330), .A4(new_n291), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n327), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G227gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT32), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(G15gat), .B(G43gat), .Z(new_n340));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n337), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n328), .A2(new_n331), .A3(new_n334), .A4(new_n332), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT34), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT32), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n333), .B2(new_n335), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT33), .B1(new_n333), .B2(new_n335), .ZN(new_n349));
  INV_X1    g148(.A(new_n342), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n343), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n343), .A2(KEYINPUT74), .A3(new_n346), .A4(new_n351), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n357));
  AOI221_X4 g156(.A(new_n347), .B1(KEYINPUT33), .B2(new_n342), .C1(new_n333), .C2(new_n335), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT73), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n346), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n361), .A3(new_n351), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G141gat), .B(G148gat), .Z(new_n364));
  INV_X1    g163(.A(G155gat), .ZN(new_n365));
  INV_X1    g164(.A(G162gat), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT2), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G155gat), .B(G162gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n364), .A2(new_n369), .A3(new_n367), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n377));
  OR2_X1    g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(G197gat), .A2(G204gat), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n380), .A2(new_n381), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT3), .B1(new_n387), .B2(new_n375), .ZN(new_n388));
  INV_X1    g187(.A(new_n373), .ZN(new_n389));
  OAI22_X1  g188(.A1(new_n376), .A2(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G78gat), .B(G106gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(new_n241), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT31), .B(G50gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n392), .B(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n387), .ZN(new_n398));
  AND2_X1   g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n316), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n316), .B2(new_n375), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n329), .B2(new_n291), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n387), .B(new_n400), .C1(new_n404), .C2(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n403), .A2(new_n405), .A3(KEYINPUT30), .A4(new_n409), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT76), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n374), .A2(new_n327), .A3(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n321), .A2(new_n326), .A3(new_n371), .A4(new_n372), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT4), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n416), .A2(new_n419), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n327), .A2(new_n373), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n417), .ZN(new_n426));
  INV_X1    g225(.A(new_n420), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n327), .A2(KEYINPUT78), .A3(new_n373), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(KEYINPUT5), .A3(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n415), .A2(new_n327), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n431), .B2(new_n374), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n417), .A2(new_n421), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n418), .A2(KEYINPUT4), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G1gat), .B(G29gat), .Z(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G57gat), .B(G85gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n444));
  INV_X1    g243(.A(new_n442), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n436), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n437), .A2(KEYINPUT6), .A3(new_n442), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n403), .A2(new_n409), .A3(new_n405), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n447), .A2(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT76), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n411), .A2(new_n452), .A3(new_n412), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n414), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n356), .A2(new_n363), .A3(new_n397), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n447), .A2(new_n448), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT35), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n397), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n450), .A2(new_n449), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(new_n411), .A3(new_n412), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n360), .B1(new_n357), .B2(new_n358), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n356), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n356), .A2(new_n462), .A3(KEYINPUT81), .A4(new_n463), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n456), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n397), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n435), .A2(new_n434), .ZN(new_n470));
  INV_X1    g269(.A(new_n416), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n427), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n426), .A2(new_n428), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n420), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(KEYINPUT39), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT39), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n476), .B(new_n427), .C1(new_n470), .C2(new_n471), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n445), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT40), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n443), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n472), .A2(KEYINPUT39), .A3(new_n474), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n477), .A2(new_n445), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT80), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n478), .A2(KEYINPUT80), .A3(new_n479), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n480), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n469), .B1(new_n487), .B2(new_n461), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n409), .B1(new_n406), .B2(KEYINPUT37), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(KEYINPUT37), .B2(new_n406), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT38), .ZN(new_n491));
  INV_X1    g290(.A(new_n457), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n489), .B(new_n493), .C1(KEYINPUT37), .C2(new_n406), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n491), .A2(new_n492), .A3(new_n450), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n414), .A2(new_n451), .A3(new_n453), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n488), .A2(new_n495), .B1(new_n469), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n356), .A2(new_n498), .A3(new_n463), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n356), .A2(new_n363), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n497), .B(new_n499), .C1(new_n500), .C2(new_n498), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n273), .B1(new_n468), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT21), .ZN(new_n503));
  OR2_X1    g302(.A1(G57gat), .A2(G64gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(G57gat), .A2(G64gat), .ZN(new_n505));
  AND2_X1   g304(.A1(G71gat), .A2(G78gat), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(KEYINPUT9), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G71gat), .B(G78gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n249), .B1(new_n503), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(G231gat), .A3(G233gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(G231gat), .A2(G233gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n511), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G127gat), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n519), .A2(G127gat), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n513), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n522), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n512), .A3(new_n520), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT88), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G155gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(G183gat), .B(G211gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT89), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n528), .B(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n523), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n523), .B2(new_n525), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G190gat), .B(G218gat), .Z(new_n535));
  NAND2_X1  g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536));
  INV_X1    g335(.A(G85gat), .ZN(new_n537));
  INV_X1    g336(.A(G92gat), .ZN(new_n538));
  AOI22_X1  g337(.A1(KEYINPUT8), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT90), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n543));
  AND2_X1   g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT91), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n541), .A2(new_n543), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n542), .B2(KEYINPUT7), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n545), .B1(new_n550), .B2(new_n541), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n539), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G99gat), .B(G106gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n553), .B(new_n539), .C1(new_n549), .C2(new_n551), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(KEYINPUT92), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n552), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n559), .A3(new_n553), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n231), .A3(new_n560), .ZN(new_n561));
  AND3_X1   g360(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n557), .A2(new_n560), .B1(new_n229), .B2(new_n226), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n535), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n557), .A2(new_n560), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n252), .ZN(new_n568));
  INV_X1    g367(.A(new_n535), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n561), .A4(new_n563), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G134gat), .B(G162gat), .Z(new_n572));
  AOI21_X1  g371(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT93), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n574), .B(KEYINPUT93), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n566), .A2(new_n570), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n534), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n534), .A2(KEYINPUT94), .A3(new_n579), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G176gat), .B(G204gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT95), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n557), .A2(new_n511), .A3(new_n560), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g391(.A(new_n511), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n556), .A3(new_n555), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n567), .A2(KEYINPUT10), .A3(new_n593), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n589), .B1(new_n591), .B2(new_n594), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n588), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n601), .B(new_n588), .C1(new_n597), .C2(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n589), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n595), .B2(new_n596), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n605), .A2(new_n588), .A3(new_n598), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n584), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n502), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n492), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g412(.A(new_n235), .B1(new_n611), .B2(new_n461), .ZN(new_n614));
  INV_X1    g413(.A(new_n461), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT16), .B(G8gat), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n610), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT42), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(KEYINPUT42), .B2(new_n617), .ZN(G1325gat));
  OAI21_X1  g418(.A(new_n499), .B1(new_n500), .B2(new_n498), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(G15gat), .B1(new_n610), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n356), .A2(new_n463), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n243), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n622), .B1(new_n610), .B2(new_n625), .ZN(G1326gat));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n469), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT43), .B(G22gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n628), .B(new_n630), .ZN(G1327gat));
  NOR3_X1   g430(.A1(new_n608), .A2(new_n534), .A3(new_n579), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n502), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n202), .A3(new_n492), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT45), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n468), .A2(new_n501), .ZN(new_n637));
  INV_X1    g436(.A(new_n579), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(KEYINPUT99), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n637), .A2(KEYINPUT99), .A3(KEYINPUT44), .A4(new_n638), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n606), .B1(new_n600), .B2(new_n602), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT98), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n646), .A2(new_n273), .A3(new_n534), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n643), .A2(new_n492), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n636), .B1(new_n202), .B2(new_n648), .ZN(G1328gat));
  NAND4_X1  g448(.A1(new_n641), .A2(new_n461), .A3(new_n642), .A4(new_n647), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n203), .B1(new_n650), .B2(KEYINPUT100), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(KEYINPUT100), .B2(new_n650), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n633), .A2(G36gat), .A3(new_n615), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT46), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(G1329gat));
  NAND4_X1  g454(.A1(new_n641), .A2(new_n620), .A3(new_n642), .A4(new_n647), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(G43gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n634), .A2(new_n214), .A3(new_n624), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT101), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT47), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1330gat));
  INV_X1    g460(.A(KEYINPUT48), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n641), .A2(new_n469), .A3(new_n642), .A4(new_n647), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G50gat), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n664), .B2(KEYINPUT103), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n634), .A2(KEYINPUT102), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667));
  AOI211_X1 g466(.A(G50gat), .B(new_n397), .C1(new_n633), .C2(new_n667), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n666), .A2(new_n668), .B1(new_n663), .B2(G50gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n665), .B(new_n669), .ZN(G1331gat));
  NOR3_X1   g469(.A1(new_n584), .A2(new_n272), .A3(new_n645), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n637), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n457), .B(KEYINPUT104), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g474(.A(new_n615), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT105), .Z(new_n677));
  NAND2_X1  g476(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(G1333gat));
  INV_X1    g479(.A(G71gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n672), .A2(new_n681), .A3(new_n624), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n672), .A2(new_n620), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g484(.A1(new_n672), .A2(new_n469), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g486(.A1(new_n534), .A2(new_n644), .A3(new_n272), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n643), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G85gat), .B1(new_n689), .B2(new_n457), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n534), .A2(new_n272), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n637), .A2(new_n638), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT51), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n694), .A2(new_n537), .A3(new_n492), .A4(new_n608), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n690), .A2(new_n695), .ZN(G1336gat));
  INV_X1    g495(.A(KEYINPUT52), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n641), .A2(new_n461), .A3(new_n642), .A4(new_n688), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G92gat), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n645), .A2(G92gat), .A3(new_n615), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n694), .A2(KEYINPUT109), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT109), .B1(new_n694), .B2(new_n700), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n697), .B(new_n699), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n692), .A2(KEYINPUT107), .A3(new_n693), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n693), .A2(KEYINPUT107), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n637), .A2(new_n638), .A3(new_n691), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n700), .B(KEYINPUT106), .Z(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n699), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT108), .B1(new_n710), .B2(KEYINPUT52), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n712), .B(new_n697), .C1(new_n699), .C2(new_n709), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n703), .B1(new_n711), .B2(new_n713), .ZN(G1337gat));
  OAI21_X1  g513(.A(G99gat), .B1(new_n689), .B2(new_n621), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n623), .A2(G99gat), .A3(new_n644), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n694), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(G1338gat));
  NAND4_X1  g517(.A1(new_n641), .A2(new_n469), .A3(new_n642), .A4(new_n688), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G106gat), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n645), .A2(G106gat), .A3(new_n397), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n707), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT53), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT53), .B1(new_n694), .B2(new_n721), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n725), .A2(KEYINPUT110), .A3(new_n720), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT110), .B1(new_n725), .B2(new_n720), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(G1339gat));
  NAND4_X1  g527(.A1(new_n582), .A2(new_n273), .A3(new_n583), .A4(new_n644), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n595), .A2(new_n596), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n589), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n595), .A2(new_n596), .A3(new_n590), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(KEYINPUT54), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n587), .B1(new_n597), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(KEYINPUT55), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(new_n607), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n595), .A2(new_n596), .A3(new_n590), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT54), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n740), .A2(new_n605), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n590), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n730), .A2(new_n743), .A3(new_n734), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n588), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n739), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n251), .B1(new_n250), .B2(new_n253), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n259), .A2(new_n260), .A3(new_n258), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n267), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n271), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n576), .B2(new_n578), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n737), .A2(new_n738), .A3(new_n746), .A4(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n746), .A2(new_n751), .A3(new_n607), .A4(new_n736), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT112), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756));
  INV_X1    g555(.A(new_n750), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n608), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT113), .B1(new_n644), .B2(new_n750), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n746), .A2(new_n272), .A3(new_n607), .A4(new_n736), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n755), .B1(new_n579), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n729), .B1(new_n762), .B2(new_n534), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n763), .A2(new_n615), .A3(new_n673), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n500), .A2(new_n397), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n766), .A2(G113gat), .A3(new_n273), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n761), .A2(new_n579), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n752), .A2(new_n754), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n534), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n729), .ZN(new_n771));
  OAI211_X1 g570(.A(KEYINPUT114), .B(new_n397), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT114), .B1(new_n763), .B2(new_n397), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n615), .A2(new_n492), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n623), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n272), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n767), .B1(new_n779), .B2(G113gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT115), .ZN(G1340gat));
  INV_X1    g580(.A(new_n778), .ZN(new_n782));
  OAI21_X1  g581(.A(G120gat), .B1(new_n782), .B2(new_n645), .ZN(new_n783));
  INV_X1    g582(.A(new_n766), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n325), .A3(new_n608), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1341gat));
  INV_X1    g585(.A(new_n534), .ZN(new_n787));
  OAI21_X1  g586(.A(G127gat), .B1(new_n782), .B2(new_n787), .ZN(new_n788));
  OR3_X1    g587(.A1(new_n766), .A2(G127gat), .A3(new_n787), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1342gat));
  NOR3_X1   g589(.A1(new_n766), .A2(G134gat), .A3(new_n579), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT56), .ZN(new_n792));
  OAI21_X1  g591(.A(G134gat), .B1(new_n782), .B2(new_n579), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1343gat));
  NOR2_X1   g593(.A1(new_n620), .A2(new_n397), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n764), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(G141gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n798), .A3(new_n272), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n763), .A2(new_n800), .A3(new_n469), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n620), .A2(new_n776), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n608), .A2(new_n757), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n733), .A2(new_n735), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT55), .B1(new_n805), .B2(KEYINPUT116), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n733), .A2(new_n807), .A3(new_n735), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n737), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n272), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n736), .A2(new_n607), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n806), .B2(new_n808), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(KEYINPUT117), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n804), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n579), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n534), .B1(new_n817), .B2(new_n769), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n469), .B1(new_n818), .B2(new_n771), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n803), .B1(new_n819), .B2(KEYINPUT57), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n272), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n799), .B1(new_n821), .B2(new_n798), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g622(.A(G148gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n797), .A2(new_n824), .A3(new_n608), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n763), .A2(KEYINPUT57), .A3(new_n469), .ZN(new_n827));
  INV_X1    g626(.A(new_n753), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n816), .B2(new_n579), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n729), .B1(new_n829), .B2(new_n534), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT57), .B1(new_n830), .B2(new_n469), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n273), .B1(new_n814), .B2(KEYINPUT117), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n810), .A2(new_n811), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n834), .A2(new_n835), .B1(new_n608), .B2(new_n757), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n753), .B1(new_n836), .B2(new_n638), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n771), .B1(new_n837), .B2(new_n787), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n800), .B1(new_n838), .B2(new_n397), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n608), .B(new_n802), .C1(new_n833), .C2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n826), .B1(new_n841), .B2(G148gat), .ZN(new_n842));
  AOI211_X1 g641(.A(KEYINPUT59), .B(new_n824), .C1(new_n820), .C2(new_n608), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n825), .B1(new_n842), .B2(new_n843), .ZN(G1345gat));
  NAND3_X1  g643(.A1(new_n797), .A2(new_n365), .A3(new_n534), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n820), .A2(new_n534), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n365), .ZN(G1346gat));
  AOI21_X1  g646(.A(G162gat), .B1(new_n797), .B2(new_n638), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n579), .A2(new_n366), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n820), .B2(new_n849), .ZN(G1347gat));
  NOR2_X1   g649(.A1(new_n673), .A2(new_n615), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n624), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n773), .B2(new_n774), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n855), .A2(G169gat), .A3(new_n272), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n768), .A2(new_n769), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n771), .B1(new_n857), .B2(new_n787), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n492), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n765), .A2(new_n461), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G169gat), .B1(new_n862), .B2(new_n272), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n856), .A2(new_n863), .ZN(G1348gat));
  NOR3_X1   g663(.A1(new_n861), .A2(G176gat), .A3(new_n644), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n855), .A2(new_n646), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(G176gat), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT119), .ZN(G1349gat));
  NOR2_X1   g667(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n869));
  OAI21_X1  g668(.A(G183gat), .B1(new_n854), .B2(new_n787), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n862), .A2(new_n277), .A3(new_n534), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n872), .B(new_n873), .Z(G1350gat));
  NOR2_X1   g673(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n638), .B(new_n853), .C1(new_n773), .C2(new_n774), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n876), .A2(KEYINPUT121), .A3(G190gat), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT121), .B1(new_n876), .B2(G190gat), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n858), .B2(new_n469), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n579), .B(new_n852), .C1(new_n882), .C2(new_n772), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n880), .B1(new_n883), .B2(new_n280), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n876), .A2(KEYINPUT121), .A3(G190gat), .ZN(new_n885));
  XOR2_X1   g684(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n862), .A2(new_n280), .A3(new_n638), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n879), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n879), .A2(new_n887), .A3(KEYINPUT123), .A4(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1351gat));
  NAND2_X1  g692(.A1(new_n621), .A2(new_n851), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n894), .B(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n827), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n839), .B2(KEYINPUT118), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n831), .A2(new_n832), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G197gat), .B1(new_n901), .B2(new_n273), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n795), .A2(new_n461), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT124), .ZN(new_n904));
  INV_X1    g703(.A(new_n859), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n273), .A2(G197gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(KEYINPUT125), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n906), .A2(new_n910), .A3(new_n907), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n902), .B1(new_n909), .B2(new_n911), .ZN(G1352gat));
  OAI21_X1  g711(.A(G204gat), .B1(new_n901), .B2(new_n645), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n644), .A2(G204gat), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OR3_X1    g714(.A1(new_n906), .A2(KEYINPUT62), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT62), .B1(new_n906), .B2(new_n915), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n913), .A2(new_n916), .A3(new_n917), .ZN(G1353gat));
  NOR3_X1   g717(.A1(new_n620), .A2(new_n615), .A3(new_n673), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n534), .B(new_n919), .C1(new_n833), .C2(new_n840), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n920), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT63), .B1(new_n920), .B2(G211gat), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n787), .A2(G211gat), .ZN(new_n923));
  OAI22_X1  g722(.A1(new_n921), .A2(new_n922), .B1(new_n906), .B2(new_n923), .ZN(G1354gat));
  OAI21_X1  g723(.A(new_n638), .B1(new_n900), .B2(KEYINPUT127), .ZN(new_n925));
  INV_X1    g724(.A(new_n896), .ZN(new_n926));
  OAI211_X1 g725(.A(KEYINPUT127), .B(new_n926), .C1(new_n833), .C2(new_n840), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G218gat), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  OR3_X1    g728(.A1(new_n906), .A2(G218gat), .A3(new_n579), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1355gat));
endmodule


