//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(KEYINPUT92), .A3(new_n205), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n206), .B(G8gat), .C1(KEYINPUT92), .C2(new_n205), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(new_n208), .A3(new_n205), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n209), .A2(KEYINPUT93), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(KEYINPUT93), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(new_n212), .B(KEYINPUT94), .Z(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n214), .B(KEYINPUT14), .Z(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT89), .B(G29gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT90), .B(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  AND2_X1   g019(.A1(G43gat), .A2(G50gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G43gat), .A2(G50gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OR3_X1    g022(.A1(new_n219), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT91), .B(G43gat), .Z(new_n225));
  INV_X1    g024(.A(G50gat), .ZN(new_n226));
  AOI211_X1 g025(.A(KEYINPUT15), .B(new_n221), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n227), .A2(new_n219), .B1(new_n220), .B2(new_n223), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT17), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n213), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n229), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n212), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n212), .B(new_n229), .Z(new_n237));
  XOR2_X1   g036(.A(new_n235), .B(KEYINPUT13), .Z(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n231), .A2(new_n235), .A3(new_n233), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G197gat), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT11), .B(G169gat), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT12), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n248), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n236), .A2(new_n250), .A3(new_n239), .A4(new_n242), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n254));
  NAND2_X1  g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255));
  INV_X1    g054(.A(G169gat), .ZN(new_n256));
  INV_X1    g055(.A(G176gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT26), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT26), .B1(new_n256), .B2(new_n257), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT65), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(G183gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT27), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT27), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G183gat), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n265), .A2(new_n267), .A3(new_n269), .A4(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT65), .B(G190gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT27), .B(G183gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n278));
  AND3_X1   g077(.A1(new_n273), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT68), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n274), .A2(new_n275), .A3(new_n282), .A4(KEYINPUT28), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n263), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(G127gat), .A2(G134gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT69), .B(G134gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(G127gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(G113gat), .B2(G120gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G113gat), .ZN(new_n292));
  INV_X1    g091(.A(G120gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n286), .ZN(new_n295));
  NAND2_X1  g094(.A1(G127gat), .A2(G134gat), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n290), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT70), .B(G120gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G113gat), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n288), .A2(new_n294), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n255), .A2(KEYINPUT24), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n306));
  OR3_X1    g105(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n258), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT23), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n261), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n301), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n312), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n274), .A2(new_n268), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n305), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT25), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n285), .A2(new_n300), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n273), .A2(new_n277), .A3(new_n278), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n281), .A3(new_n283), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n323), .A2(new_n263), .B1(new_n313), .B2(new_n317), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(KEYINPUT71), .A3(new_n300), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n285), .A2(new_n318), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n288), .A2(new_n294), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n297), .A2(new_n299), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n321), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n254), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n300), .B1(new_n285), .B2(new_n318), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n320), .B2(new_n319), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT34), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n332), .A4(new_n325), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT32), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n331), .B2(new_n333), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT33), .B1(new_n331), .B2(new_n333), .ZN(new_n342));
  XNOR2_X1  g141(.A(G15gat), .B(G43gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(KEYINPUT72), .ZN(new_n344));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n341), .A2(new_n342), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(KEYINPUT33), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(KEYINPUT32), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n339), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT74), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n355), .B(new_n339), .C1(new_n348), .C2(new_n352), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n358));
  OR2_X1    g157(.A1(KEYINPUT81), .A2(G148gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(KEYINPUT81), .A2(G148gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(G141gat), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G148gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(G141gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  OR2_X1    g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n361), .A2(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT82), .B(G162gat), .ZN(new_n368));
  INV_X1    g167(.A(G155gat), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT2), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G141gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(G148gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT2), .ZN(new_n374));
  OAI22_X1  g173(.A1(new_n363), .A2(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n365), .A2(new_n373), .ZN(new_n376));
  NAND3_X1  g175(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n376), .A2(new_n366), .A3(new_n377), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n367), .A2(new_n370), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(new_n300), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT83), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n358), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n375), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n365), .ZN(new_n385));
  INV_X1    g184(.A(new_n360), .ZN(new_n386));
  NOR2_X1   g185(.A1(KEYINPUT81), .A2(G148gat), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n386), .A2(new_n387), .A3(new_n371), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n385), .B1(new_n388), .B2(new_n363), .ZN(new_n389));
  XOR2_X1   g188(.A(KEYINPUT82), .B(G162gat), .Z(new_n390));
  AOI21_X1  g189(.A(new_n374), .B1(new_n390), .B2(G155gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n384), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n395), .A3(new_n329), .ZN(new_n396));
  INV_X1    g195(.A(new_n382), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(new_n392), .B2(new_n329), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n300), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n396), .A2(new_n397), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n403), .A2(new_n358), .A3(new_n397), .A4(new_n396), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT0), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT84), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n409), .B1(new_n402), .B2(new_n404), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT6), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n414), .A2(KEYINPUT6), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n404), .A3(new_n409), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G226gat), .ZN(new_n422));
  INV_X1    g221(.A(G233gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n326), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n424), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n324), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G197gat), .B(G204gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT22), .ZN(new_n430));
  INV_X1    g229(.A(G211gat), .ZN(new_n431));
  INV_X1    g230(.A(G218gat), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G211gat), .B(G218gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n429), .A3(new_n433), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n426), .A2(new_n428), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(KEYINPUT77), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n427), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n326), .A2(new_n424), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT78), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G8gat), .B(G36gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(G64gat), .B(G92gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n441), .B1(new_n426), .B2(new_n428), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT78), .ZN(new_n452));
  INV_X1    g251(.A(new_n439), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n443), .A2(new_n453), .A3(new_n444), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n446), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n450), .B1(new_n451), .B2(new_n454), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(KEYINPUT30), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT79), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n457), .A2(new_n459), .A3(KEYINPUT30), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n457), .B2(KEYINPUT30), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n456), .B(new_n458), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n439), .A2(new_n425), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT3), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n465), .B2(new_n464), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n395), .A2(new_n425), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n467), .A2(new_n392), .B1(new_n453), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(G228gat), .A2(G233gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n464), .A2(new_n379), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n393), .A2(new_n470), .ZN(new_n473));
  AOI211_X1 g272(.A(new_n472), .B(new_n473), .C1(new_n442), .C2(new_n468), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G78gat), .B(G106gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT31), .B(G50gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G22gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(KEYINPUT86), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n480), .B1(new_n482), .B2(new_n478), .ZN(new_n483));
  XOR2_X1   g282(.A(new_n475), .B(new_n483), .Z(new_n484));
  NAND2_X1  g283(.A1(new_n349), .A2(KEYINPUT32), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n349), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n487), .A3(new_n346), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n351), .A2(new_n334), .A3(new_n338), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n484), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n357), .A2(new_n421), .A3(new_n463), .A4(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n461), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n457), .A2(new_n459), .A3(KEYINPUT30), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n458), .A2(new_n456), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n421), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n497), .A2(KEYINPUT35), .A3(new_n484), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT76), .B1(new_n348), .B2(new_n489), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT76), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n334), .A2(new_n338), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n488), .A2(new_n500), .A3(new_n501), .A4(new_n351), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n353), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n492), .A2(KEYINPUT35), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n490), .B2(new_n488), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n354), .A2(new_n356), .A3(new_n510), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n508), .A2(new_n511), .B1(new_n484), .B2(new_n497), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n446), .A2(KEYINPUT37), .A3(new_n455), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n451), .A2(new_n454), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n449), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT38), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n413), .A2(new_n416), .B1(new_n419), .B2(new_n418), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n426), .A2(new_n428), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n516), .B1(new_n521), .B2(new_n442), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n439), .B1(new_n426), .B2(new_n428), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT38), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n457), .B1(new_n524), .B2(new_n517), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n329), .B1(new_n379), .B2(new_n394), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n367), .A2(new_n370), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n528), .A2(new_n394), .A3(new_n384), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n399), .B(new_n400), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n382), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT87), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT87), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n533), .A3(new_n382), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT39), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n410), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n380), .A2(new_n382), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(new_n536), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n532), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT40), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n530), .A2(new_n533), .A3(new_n382), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n533), .B1(new_n530), .B2(new_n382), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n536), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n544), .A2(new_n540), .A3(KEYINPUT40), .A4(new_n409), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n411), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n462), .ZN(new_n548));
  INV_X1    g347(.A(new_n484), .ZN(new_n549));
  AND4_X1   g348(.A1(new_n513), .A2(new_n526), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n484), .B1(new_n547), .B2(new_n462), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n513), .B1(new_n551), .B2(new_n526), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n512), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n253), .B1(new_n506), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT96), .ZN(new_n556));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G71gat), .B(G78gat), .ZN(new_n560));
  INV_X1    g359(.A(G57gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(KEYINPUT95), .A3(G64gat), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n556), .A2(new_n559), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT97), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(new_n560), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(KEYINPUT21), .ZN(new_n569));
  AND2_X1   g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G127gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n212), .B1(new_n568), .B2(KEYINPUT21), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT98), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G155gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n576), .B(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n583), .A2(KEYINPUT99), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT7), .B1(new_n583), .B2(KEYINPUT99), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n586), .B(new_n590), .C1(new_n584), .C2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  NOR2_X1   g393(.A1(new_n230), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n232), .A2(new_n594), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT41), .ZN(new_n597));
  NAND2_X1  g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n597), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n602), .A2(KEYINPUT100), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n605), .B(KEYINPUT100), .Z(new_n608));
  NOR2_X1   g407(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n568), .A2(new_n594), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n568), .A2(new_n594), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT10), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(new_n616), .A3(new_n613), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n568), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n615), .B1(new_n619), .B2(new_n611), .ZN(new_n620));
  INV_X1    g419(.A(new_n611), .ZN(new_n621));
  AOI211_X1 g420(.A(KEYINPUT101), .B(new_n621), .C1(new_n617), .C2(new_n618), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OR4_X1    g425(.A1(new_n614), .A2(new_n620), .A3(new_n622), .A4(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n619), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n621), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n626), .B1(new_n629), .B2(new_n614), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n582), .A2(new_n610), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n554), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(new_n421), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(G1gat), .Z(G1324gat));
  INV_X1    g434(.A(KEYINPUT42), .ZN(new_n636));
  OAI21_X1  g435(.A(G8gat), .B1(new_n633), .B2(new_n463), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT16), .B(G8gat), .Z(new_n638));
  NAND4_X1  g437(.A1(new_n554), .A2(new_n462), .A3(new_n632), .A4(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n636), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n636), .B2(new_n639), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT102), .Z(G1325gat));
  NAND2_X1  g441(.A1(new_n508), .A2(new_n511), .ZN(new_n643));
  OAI21_X1  g442(.A(G15gat), .B1(new_n633), .B2(new_n643), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n503), .A2(G15gat), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n633), .B2(new_n645), .ZN(G1326gat));
  NOR2_X1   g445(.A1(new_n633), .A2(new_n549), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT43), .B(G22gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n553), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n512), .B(KEYINPUT104), .C1(new_n550), .C2(new_n552), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n505), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n610), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n506), .A2(new_n553), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(KEYINPUT44), .A3(new_n610), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n582), .B(KEYINPUT103), .ZN(new_n660));
  INV_X1    g459(.A(new_n631), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n252), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n216), .B1(new_n664), .B2(new_n421), .ZN(new_n665));
  INV_X1    g464(.A(new_n582), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n666), .A2(new_n655), .A3(new_n631), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n554), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(new_n421), .A3(new_n216), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT45), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n670), .ZN(G1328gat));
  OAI21_X1  g470(.A(new_n217), .B1(new_n664), .B2(new_n463), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n668), .A2(new_n463), .A3(new_n217), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT46), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(G1329gat));
  INV_X1    g474(.A(new_n643), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n663), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n225), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n668), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n504), .A3(new_n225), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT47), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685));
  AOI211_X1 g484(.A(KEYINPUT105), .B(new_n685), .C1(new_n679), .C2(new_n681), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n684), .A2(new_n686), .ZN(G1330gat));
  AND2_X1   g486(.A1(new_n680), .A2(KEYINPUT106), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n680), .A2(KEYINPUT106), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n484), .A2(new_n226), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n663), .A2(new_n484), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n692), .B2(G50gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g493(.A1(new_n666), .A2(new_n253), .A3(new_n655), .A4(new_n631), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n654), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n520), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g497(.A(new_n463), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT107), .ZN(new_n701));
  NOR2_X1   g500(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1333gat));
  INV_X1    g502(.A(G71gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n696), .A2(new_n704), .A3(new_n504), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n654), .A2(new_n643), .A3(new_n695), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(new_n704), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g507(.A1(new_n696), .A2(new_n484), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT108), .B(G78gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1335gat));
  AND2_X1   g510(.A1(new_n656), .A2(new_n658), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n666), .A2(new_n252), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n661), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G85gat), .B1(new_n716), .B2(new_n421), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n551), .A2(new_n526), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT88), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n551), .A2(new_n513), .A3(new_n526), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT104), .B1(new_n721), .B2(new_n512), .ZN(new_n722));
  INV_X1    g521(.A(new_n653), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n506), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n725), .A3(new_n610), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT109), .B1(new_n654), .B2(new_n655), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(new_n727), .A3(new_n713), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n652), .A2(new_n653), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n655), .B1(new_n731), .B2(new_n506), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n714), .B1(new_n732), .B2(new_n725), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n727), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n631), .A2(new_n588), .A3(new_n520), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n717), .B1(new_n736), .B2(new_n737), .ZN(G1336gat));
  NOR3_X1   g537(.A1(new_n661), .A2(G92gat), .A3(new_n463), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT51), .B1(new_n733), .B2(new_n727), .ZN(new_n740));
  AND4_X1   g539(.A1(KEYINPUT51), .A2(new_n726), .A3(new_n727), .A4(new_n713), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n656), .A2(new_n462), .A3(new_n658), .A4(new_n715), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(G92gat), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT52), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(new_n735), .B2(new_n739), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n712), .A2(KEYINPUT110), .A3(new_n462), .A4(new_n715), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n589), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n747), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  AND4_X1   g553(.A1(new_n747), .A2(new_n752), .A3(new_n742), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n746), .B1(new_n753), .B2(new_n755), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n716), .B2(new_n643), .ZN(new_n757));
  OR3_X1    g556(.A1(new_n661), .A2(G99gat), .A3(new_n503), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n736), .B2(new_n758), .ZN(G1338gat));
  NOR3_X1   g558(.A1(new_n661), .A2(G106gat), .A3(new_n549), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n735), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n656), .A2(new_n484), .A3(new_n658), .A4(new_n715), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G106gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n760), .B(KEYINPUT112), .Z(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n740), .B2(new_n741), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n764), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT113), .B1(new_n768), .B2(KEYINPUT53), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n770), .B(new_n762), .C1(new_n767), .C2(new_n764), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n765), .B1(new_n769), .B2(new_n771), .ZN(G1339gat));
  NAND2_X1  g571(.A1(new_n357), .A2(new_n491), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n421), .A2(new_n462), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT54), .B1(new_n619), .B2(new_n611), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n777), .A2(new_n620), .A3(new_n622), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n619), .A2(new_n611), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n626), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n776), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n781), .ZN(new_n783));
  INV_X1    g582(.A(new_n620), .ZN(new_n784));
  INV_X1    g583(.A(new_n622), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g585(.A(KEYINPUT55), .B(new_n783), .C1(new_n786), .C2(new_n777), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n782), .A2(new_n787), .A3(new_n627), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT115), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n782), .A2(new_n787), .A3(new_n627), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n252), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n234), .A2(new_n235), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n237), .A2(new_n238), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n247), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n251), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n631), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n610), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n796), .A2(new_n610), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n789), .A3(new_n791), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n660), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NOR4_X1   g601(.A1(new_n582), .A2(new_n252), .A3(new_n610), .A4(new_n631), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n773), .B(new_n775), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n292), .A3(new_n252), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n484), .B1(new_n802), .B2(new_n804), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n775), .A2(new_n503), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(KEYINPUT116), .A3(new_n808), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n252), .A3(new_n812), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n813), .A2(KEYINPUT117), .A3(G113gat), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT117), .B1(new_n813), .B2(G113gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n806), .B1(new_n814), .B2(new_n815), .ZN(G1340gat));
  NAND2_X1  g615(.A1(new_n811), .A2(new_n812), .ZN(new_n817));
  OAI21_X1  g616(.A(G120gat), .B1(new_n817), .B2(new_n661), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n661), .A2(new_n298), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n805), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1341gat));
  OAI21_X1  g620(.A(G127gat), .B1(new_n817), .B2(new_n660), .ZN(new_n822));
  INV_X1    g621(.A(G127gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n805), .A2(new_n823), .A3(new_n666), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1342gat));
  NOR2_X1   g624(.A1(new_n655), .A2(new_n287), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n805), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT56), .Z(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n817), .B2(new_n655), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1343gat));
  AOI21_X1  g629(.A(new_n549), .B1(new_n802), .B2(new_n804), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n643), .A2(new_n774), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n797), .B1(new_n253), .B2(new_n788), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n655), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n666), .B1(new_n836), .B2(new_n800), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n484), .B1(new_n837), .B2(new_n803), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n834), .B1(new_n838), .B2(KEYINPUT57), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n833), .A2(new_n839), .A3(new_n252), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(G141gat), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n775), .B1(new_n802), .B2(new_n804), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n676), .A2(new_n549), .ZN(new_n843));
  AND4_X1   g642(.A1(new_n371), .A2(new_n842), .A3(new_n252), .A4(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(KEYINPUT118), .B(KEYINPUT58), .C1(new_n841), .C2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n840), .B2(G141gat), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT58), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n851), .B1(new_n850), .B2(new_n844), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n845), .B(new_n849), .C1(new_n841), .C2(new_n852), .ZN(G1344gat));
  AND2_X1   g652(.A1(new_n842), .A2(new_n843), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n386), .A2(new_n387), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n855), .A3(new_n631), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT120), .Z(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(KEYINPUT59), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n833), .A2(new_n839), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n661), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT121), .B(new_n858), .C1(new_n859), .C2(new_n661), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n799), .A2(new_n627), .A3(new_n787), .A4(new_n782), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n666), .B1(new_n836), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n832), .B(new_n484), .C1(new_n865), .C2(new_n803), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n834), .A2(new_n661), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n866), .B(new_n867), .C1(new_n831), .C2(new_n832), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT59), .B1(new_n869), .B2(new_n362), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n862), .A2(new_n863), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n857), .A2(new_n871), .ZN(G1345gat));
  INV_X1    g671(.A(new_n859), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n660), .A2(new_n369), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT122), .B1(new_n854), .B2(new_n666), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n842), .A2(KEYINPUT122), .A3(new_n666), .A4(new_n843), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n369), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT123), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n875), .B(new_n881), .C1(new_n876), .C2(new_n878), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1346gat));
  AOI21_X1  g682(.A(new_n390), .B1(new_n854), .B2(new_n610), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n655), .A2(new_n368), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n873), .B2(new_n885), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n463), .A2(new_n520), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n807), .A2(new_n504), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(new_n256), .A3(new_n253), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n802), .A2(new_n804), .ZN(new_n890));
  INV_X1    g689(.A(new_n887), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n773), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(G169gat), .B1(new_n894), .B2(new_n252), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n889), .A2(new_n895), .ZN(G1348gat));
  OAI21_X1  g695(.A(G176gat), .B1(new_n888), .B2(new_n661), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n257), .A3(new_n631), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1349gat));
  OAI21_X1  g698(.A(G183gat), .B1(new_n888), .B2(new_n660), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n666), .A2(new_n275), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n893), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g702(.A1(new_n894), .A2(new_n274), .A3(new_n610), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT124), .Z(new_n905));
  NOR2_X1   g704(.A1(new_n888), .A2(new_n655), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n264), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(G1351gat));
  NOR2_X1   g709(.A1(new_n676), .A2(new_n891), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n831), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n912), .A2(new_n252), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n866), .B(new_n911), .C1(new_n831), .C2(new_n832), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n252), .A2(G197gat), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n913), .A2(G197gat), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(G1352gat));
  INV_X1    g716(.A(G204gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n912), .A2(new_n918), .A3(new_n631), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT62), .Z(new_n920));
  OAI21_X1  g719(.A(G204gat), .B1(new_n914), .B2(new_n661), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1353gat));
  OAI21_X1  g721(.A(G211gat), .B1(new_n914), .B2(new_n582), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g724(.A(KEYINPUT63), .B(G211gat), .C1(new_n914), .C2(new_n582), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(KEYINPUT125), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n431), .A3(new_n666), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n927), .B(new_n928), .C1(KEYINPUT125), .C2(new_n925), .ZN(G1354gat));
  NAND3_X1  g728(.A1(new_n831), .A2(new_n610), .A3(new_n911), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n432), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n610), .A2(G218gat), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT126), .Z(new_n933));
  OAI21_X1  g732(.A(new_n931), .B1(new_n914), .B2(new_n933), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT127), .Z(G1355gat));
endmodule


