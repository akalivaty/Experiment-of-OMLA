//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT86), .Z(new_n208));
  NOR2_X1   g007(.A1(new_n202), .A2(new_n203), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(KEYINPUT15), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(new_n211), .C1(KEYINPUT15), .C2(new_n210), .ZN(new_n212));
  OAI211_X1 g011(.A(KEYINPUT15), .B(new_n210), .C1(new_n207), .C2(new_n209), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G1gat), .ZN(new_n217));
  INV_X1    g016(.A(G8gat), .ZN(new_n218));
  OAI221_X1 g017(.A(new_n217), .B1(KEYINPUT87), .B2(new_n218), .C1(G1gat), .C2(new_n215), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(KEYINPUT87), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT88), .ZN(new_n223));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n214), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n221), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n223), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT18), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n221), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n224), .B(KEYINPUT13), .Z(new_n232));
  AOI22_X1  g031(.A1(new_n228), .A2(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(new_n229), .B2(new_n228), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G141gat), .ZN(new_n235));
  INV_X1    g034(.A(G197gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT11), .B(G169gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT89), .ZN(new_n242));
  OR3_X1    g041(.A1(new_n234), .A2(KEYINPUT90), .A3(new_n240), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT90), .B1(new_n234), .B2(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n248));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G120gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(KEYINPUT1), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n251), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n249), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n259), .A2(new_n260), .B1(KEYINPUT23), .B2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n262), .B(KEYINPUT68), .Z(new_n263));
  INV_X1    g062(.A(KEYINPUT24), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(G183gat), .A3(G190gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(G183gat), .B(G190gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(new_n264), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n261), .B2(KEYINPUT23), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n271), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(KEYINPUT25), .A3(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n263), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n273), .A2(KEYINPUT66), .A3(new_n262), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT66), .B1(new_n273), .B2(new_n262), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n277), .A2(new_n278), .A3(new_n267), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n279), .B2(KEYINPUT25), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(new_n262), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n273), .A2(new_n262), .A3(KEYINPUT66), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(new_n268), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT67), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n275), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT27), .B(G183gat), .ZN(new_n289));
  INV_X1    g088(.A(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n289), .B(new_n290), .C1(new_n291), .C2(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n259), .A2(new_n260), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT26), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n261), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G183gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(new_n290), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n301), .A2(KEYINPUT70), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(KEYINPUT70), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n294), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n256), .B1(new_n288), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n275), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n267), .B1(new_n281), .B2(new_n282), .ZN(new_n307));
  AOI211_X1 g106(.A(new_n276), .B(KEYINPUT25), .C1(new_n307), .C2(new_n284), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT67), .B1(new_n285), .B2(new_n286), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n252), .A2(new_n255), .ZN(new_n311));
  INV_X1    g110(.A(new_n304), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n305), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G227gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n248), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  AOI211_X1 g116(.A(KEYINPUT71), .B(new_n315), .C1(new_n305), .C2(new_n313), .ZN(new_n318));
  XOR2_X1   g117(.A(KEYINPUT72), .B(KEYINPUT33), .Z(new_n319));
  OAI22_X1  g118(.A1(new_n317), .A2(new_n318), .B1(KEYINPUT32), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G71gat), .B(G99gat), .Z(new_n321));
  XNOR2_X1  g120(.A(G15gat), .B(G43gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n288), .A2(new_n256), .A3(new_n304), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n311), .B1(new_n310), .B2(new_n312), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n316), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT71), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n314), .A2(new_n248), .A3(new_n316), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n319), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n333), .A2(KEYINPUT32), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n325), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n334), .ZN(new_n336));
  AOI211_X1 g135(.A(KEYINPUT73), .B(new_n336), .C1(new_n329), .C2(new_n330), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n324), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n305), .A2(new_n315), .A3(new_n313), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n339), .B(KEYINPUT34), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G78gat), .B(G106gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT31), .B(G50gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT83), .ZN(new_n346));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G155gat), .B(G162gat), .ZN(new_n351));
  INV_X1    g150(.A(G162gat), .ZN(new_n352));
  INV_X1    g151(.A(G155gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT79), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G155gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT2), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n350), .B(new_n351), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT2), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n360), .A2(KEYINPUT78), .A3(new_n351), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n362));
  INV_X1    g161(.A(new_n351), .ZN(new_n363));
  INV_X1    g162(.A(new_n349), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n358), .A3(new_n347), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n359), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G197gat), .B(G204gat), .ZN(new_n368));
  XOR2_X1   g167(.A(KEYINPUT74), .B(G218gat), .Z(new_n369));
  INV_X1    g168(.A(G211gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n368), .B1(new_n371), .B2(KEYINPUT22), .ZN(new_n372));
  XNOR2_X1  g171(.A(G211gat), .B(G218gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(KEYINPUT29), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n367), .B1(new_n375), .B2(KEYINPUT3), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n367), .A2(KEYINPUT3), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n374), .B1(new_n378), .B2(KEYINPUT29), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(G22gat), .ZN(new_n381));
  INV_X1    g180(.A(G228gat), .ZN(new_n382));
  INV_X1    g181(.A(G233gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G22gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n380), .B(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(new_n384), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n346), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n384), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n381), .A2(new_n385), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT83), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .A4(new_n345), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n334), .B1(new_n317), .B2(new_n318), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT73), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n331), .A2(new_n325), .A3(new_n334), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n340), .A3(new_n324), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n342), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n310), .A2(new_n312), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n405), .B(KEYINPUT75), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n374), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n402), .A2(new_n406), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G8gat), .B(G36gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(G64gat), .B(G92gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  NAND2_X1  g213(.A1(new_n280), .A2(new_n287), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n304), .B1(new_n415), .B2(new_n306), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT76), .B1(new_n416), .B2(new_n407), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT76), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n418), .A3(new_n406), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n417), .A2(new_n419), .B1(new_n404), .B2(new_n407), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n411), .B(new_n414), .C1(new_n420), .C2(new_n409), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT77), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT30), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(KEYINPUT77), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n411), .B1(new_n420), .B2(new_n409), .ZN(new_n426));
  INV_X1    g225(.A(new_n414), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n367), .A2(new_n256), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT78), .B1(new_n360), .B2(new_n351), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n363), .A2(new_n365), .A3(new_n362), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n434), .A2(new_n359), .B1(new_n255), .B2(new_n252), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n430), .B(KEYINPUT5), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n367), .A2(new_n256), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n311), .A2(new_n434), .A3(new_n359), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT5), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT81), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n437), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n311), .B1(new_n367), .B2(KEYINPUT3), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n449), .B1(new_n377), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT82), .B1(new_n431), .B2(new_n445), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n431), .A2(new_n447), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n455), .A3(KEYINPUT4), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  AOI211_X1 g256(.A(KEYINPUT5), .B(new_n449), .C1(new_n377), .C2(new_n450), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n444), .A2(new_n452), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT0), .ZN(new_n461));
  XNOR2_X1  g260(.A(G57gat), .B(G85gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n461), .B(new_n462), .Z(new_n463));
  OAI21_X1  g262(.A(KEYINPUT84), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT6), .B1(new_n459), .B2(new_n463), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n466));
  INV_X1    g265(.A(new_n463), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n438), .A2(new_n443), .B1(new_n448), .B2(new_n451), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n458), .A2(new_n457), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n464), .A2(new_n465), .A3(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT6), .B(new_n467), .C1(new_n468), .C2(new_n470), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n401), .A2(new_n429), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n465), .B1(new_n463), .B2(new_n459), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n473), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n423), .A2(new_n480), .A3(new_n425), .A4(new_n428), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n482), .A2(new_n395), .A3(new_n342), .A4(new_n400), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n478), .B1(new_n483), .B2(KEYINPUT35), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n478), .B(KEYINPUT35), .C1(new_n401), .C2(new_n481), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n477), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n488));
  INV_X1    g287(.A(new_n400), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n340), .B1(new_n399), .B2(new_n324), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n342), .A2(KEYINPUT36), .A3(new_n400), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n390), .A2(new_n394), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n472), .A2(new_n421), .A3(new_n473), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n427), .A2(KEYINPUT37), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n428), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n420), .A2(new_n374), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n416), .A2(new_n407), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n407), .B2(new_n404), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n500), .B2(new_n374), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT38), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n494), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n426), .A2(KEYINPUT37), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n427), .B1(new_n426), .B2(KEYINPUT37), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT38), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n493), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n464), .A2(new_n471), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n377), .A2(new_n450), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n437), .B1(new_n457), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT39), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n467), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n436), .A2(new_n437), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT39), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT40), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n429), .A2(new_n508), .A3(new_n516), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n491), .A2(new_n492), .B1(new_n507), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n481), .A2(new_n493), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n247), .B1(new_n487), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522));
  INV_X1    g321(.A(G85gat), .ZN(new_n523));
  INV_X1    g322(.A(G92gat), .ZN(new_n524));
  AOI22_X1  g323(.A1(KEYINPUT8), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT93), .ZN(new_n526));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G99gat), .B(G106gat), .Z(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n530), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n226), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n536), .B(new_n537), .C1(new_n214), .C2(new_n535), .ZN(new_n538));
  XNOR2_X1  g337(.A(G190gat), .B(G218gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT95), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n539), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G134gat), .B(G162gat), .Z(new_n544));
  AOI21_X1  g343(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT92), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n546), .B1(new_n542), .B2(KEYINPUT96), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n541), .B(new_n549), .C1(KEYINPUT96), .C2(new_n542), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  INV_X1    g351(.A(G71gat), .ZN(new_n553));
  INV_X1    g352(.A(G78gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G71gat), .B(G78gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G127gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n221), .B1(new_n562), .B2(new_n563), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(new_n353), .ZN(new_n571));
  XOR2_X1   g370(.A(G183gat), .B(G211gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(new_n574), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OR3_X1    g377(.A1(new_n551), .A2(KEYINPUT97), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT97), .B1(new_n551), .B2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n535), .A2(new_n562), .ZN(new_n582));
  INV_X1    g381(.A(new_n562), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(new_n534), .A3(new_n531), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(KEYINPUT10), .ZN(new_n586));
  OAI22_X1  g385(.A1(new_n585), .A2(KEYINPUT10), .B1(new_n535), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G230gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(new_n383), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n589), .B2(new_n585), .ZN(new_n592));
  XNOR2_X1  g391(.A(G120gat), .B(G148gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  OR2_X1    g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n581), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n521), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(new_n480), .ZN(new_n601));
  XOR2_X1   g400(.A(KEYINPUT98), .B(G1gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(G1324gat));
  NAND3_X1  g402(.A1(new_n521), .A2(new_n599), .A3(new_n429), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n604), .A2(G8gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT16), .B(G8gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT42), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(KEYINPUT42), .B2(new_n607), .ZN(G1325gat));
  INV_X1    g408(.A(new_n599), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n342), .A2(new_n400), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n610), .A2(G15gat), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n521), .ZN(new_n613));
  INV_X1    g412(.A(new_n491), .ZN(new_n614));
  INV_X1    g413(.A(new_n492), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(G15gat), .B1(new_n600), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n618), .ZN(G1326gat));
  NOR2_X1   g418(.A1(new_n600), .A2(new_n395), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT99), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT43), .B(G22gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(G1327gat));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n519), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n481), .A2(KEYINPUT101), .A3(new_n493), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n518), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n518), .B2(new_n628), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT35), .B1(new_n401), .B2(new_n481), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT85), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n485), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n635), .B2(new_n477), .ZN(new_n636));
  AOI211_X1 g435(.A(KEYINPUT103), .B(new_n476), .C1(new_n634), .C2(new_n485), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n631), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n551), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n487), .A2(new_n520), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(KEYINPUT44), .A3(new_n551), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n598), .B(KEYINPUT100), .Z(new_n645));
  NOR3_X1   g444(.A1(new_n645), .A2(new_n247), .A3(new_n577), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(G29gat), .B1(new_n647), .B2(new_n480), .ZN(new_n648));
  INV_X1    g447(.A(new_n551), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n649), .A2(new_n577), .A3(new_n598), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n521), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n651), .A2(G29gat), .A3(new_n480), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT45), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n653), .ZN(G1328gat));
  INV_X1    g453(.A(new_n429), .ZN(new_n655));
  OAI21_X1  g454(.A(G36gat), .B1(new_n647), .B2(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n651), .A2(G36gat), .A3(new_n655), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT46), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(G1329gat));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660));
  OAI21_X1  g459(.A(G43gat), .B1(new_n647), .B2(new_n617), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n651), .A2(G43gat), .A3(new_n611), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT105), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n660), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g464(.A(G50gat), .B1(new_n647), .B2(new_n395), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n651), .A2(G50gat), .A3(new_n395), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT107), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(KEYINPUT107), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n666), .A2(new_n669), .A3(KEYINPUT48), .A4(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n672), .A2(new_n673), .A3(new_n667), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n671), .B1(new_n674), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g474(.A(new_n638), .ZN(new_n676));
  INV_X1    g475(.A(new_n645), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n676), .A2(new_n246), .A3(new_n581), .A4(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n480), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT108), .B(G57gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1332gat));
  AOI21_X1  g481(.A(new_n655), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT109), .Z(new_n685));
  NOR2_X1   g484(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1333gat));
  AOI21_X1  g486(.A(new_n553), .B1(new_n678), .B2(new_n616), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n611), .A2(G71gat), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n678), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1334gat));
  NAND2_X1  g491(.A1(new_n678), .A2(new_n493), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g493(.A1(new_n246), .A2(new_n577), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n598), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n644), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n679), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n523), .B1(new_n700), .B2(KEYINPUT111), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(KEYINPUT111), .B2(new_n700), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT51), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n638), .A2(new_n704), .A3(new_n551), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n695), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n638), .B2(new_n551), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n639), .A2(KEYINPUT112), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n709), .A2(KEYINPUT51), .A3(new_n695), .A4(new_n705), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n598), .A2(new_n523), .A3(new_n679), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT113), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n702), .B1(new_n712), .B2(new_n714), .ZN(G1336gat));
  NOR3_X1   g514(.A1(new_n677), .A2(G92gat), .A3(new_n655), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n487), .A2(KEYINPUT103), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n635), .A2(new_n632), .A3(new_n477), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n649), .B1(new_n719), .B2(new_n631), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n696), .B1(new_n720), .B2(new_n704), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT51), .B1(new_n721), .B2(new_n709), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n706), .A2(new_n703), .A3(new_n707), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n716), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n641), .A2(new_n429), .A3(new_n643), .A4(new_n698), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G92gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT116), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT115), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT114), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n724), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n716), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n708), .B2(new_n710), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT114), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n733), .A2(new_n736), .A3(new_n727), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n731), .B1(new_n737), .B2(KEYINPUT52), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n727), .B1(new_n735), .B2(KEYINPUT114), .ZN(new_n739));
  AOI211_X1 g538(.A(new_n732), .B(new_n734), .C1(new_n708), .C2(new_n710), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n731), .B(KEYINPUT52), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n730), .B1(new_n738), .B2(new_n742), .ZN(G1337gat));
  NOR4_X1   g542(.A1(new_n712), .A2(G99gat), .A3(new_n611), .A4(new_n697), .ZN(new_n744));
  INV_X1    g543(.A(G99gat), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n699), .B2(new_n616), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n744), .A2(new_n746), .ZN(G1338gat));
  NAND2_X1  g546(.A1(new_n699), .A2(new_n493), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n677), .A2(G106gat), .A3(new_n395), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n748), .A2(G106gat), .B1(new_n711), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT53), .Z(G1339gat));
  NAND2_X1  g550(.A1(new_n599), .A2(new_n247), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n591), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n590), .B2(new_n587), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n595), .B1(new_n591), .B2(new_n753), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT55), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n597), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n757), .A2(KEYINPUT55), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n223), .A2(new_n227), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(G229gat), .A3(G233gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n231), .B2(new_n232), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n243), .A2(new_n244), .B1(new_n239), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n761), .A2(new_n551), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n598), .ZN(new_n767));
  INV_X1    g566(.A(new_n761), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(new_n247), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n766), .B1(new_n769), .B2(new_n649), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n752), .B1(new_n770), .B2(new_n577), .ZN(new_n771));
  INV_X1    g570(.A(new_n401), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n429), .A2(new_n480), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n246), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G113gat), .ZN(G1340gat));
  AOI21_X1  g575(.A(G120gat), .B1(new_n774), .B2(new_n598), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n645), .A2(G120gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n774), .B2(new_n778), .ZN(G1341gat));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n774), .B(new_n577), .C1(new_n780), .C2(G127gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(KEYINPUT118), .B2(G127gat), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n781), .B(new_n782), .Z(G1342gat));
  AOI21_X1  g582(.A(new_n649), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n774), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n785), .B(new_n786), .Z(G1343gat));
  INV_X1    g586(.A(G141gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n616), .A2(new_n395), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(KEYINPUT122), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n790), .A2(KEYINPUT122), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n788), .B1(new_n793), .B2(new_n247), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n616), .A2(new_n480), .A3(new_n429), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n493), .A2(KEYINPUT57), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT120), .B1(new_n759), .B2(new_n760), .ZN(new_n797));
  INV_X1    g596(.A(new_n760), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n798), .A2(new_n799), .A3(new_n597), .A4(new_n758), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n800), .A3(new_n246), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n767), .B(KEYINPUT119), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n551), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n578), .B1(new_n803), .B2(new_n766), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n804), .A2(new_n805), .B1(new_n247), .B2(new_n599), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n796), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT57), .B1(new_n771), .B2(new_n493), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n795), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n247), .A2(new_n788), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n794), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n794), .B(KEYINPUT58), .C1(new_n810), .C2(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1344gat));
  OR3_X1    g616(.A1(new_n810), .A2(KEYINPUT59), .A3(new_n697), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT59), .B1(new_n793), .B2(new_n697), .ZN(new_n819));
  INV_X1    g618(.A(G148gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n752), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT57), .B1(new_n822), .B2(new_n493), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n771), .A2(KEYINPUT57), .A3(new_n493), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n795), .A2(new_n598), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT59), .B(G148gat), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n818), .A2(new_n821), .A3(new_n827), .ZN(G1345gat));
  NAND2_X1  g627(.A1(new_n354), .A2(new_n356), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n810), .B2(new_n578), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n577), .A2(new_n354), .A3(new_n356), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n793), .B2(new_n831), .ZN(G1346gat));
  OAI21_X1  g631(.A(G162gat), .B1(new_n810), .B2(new_n649), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n791), .A2(new_n352), .A3(new_n551), .A4(new_n792), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(KEYINPUT123), .A3(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1347gat));
  NAND2_X1  g638(.A1(new_n771), .A2(new_n480), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n401), .A2(new_n655), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(KEYINPUT124), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(KEYINPUT124), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(G169gat), .B1(new_n844), .B2(new_n246), .ZN(new_n845));
  INV_X1    g644(.A(new_n841), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n246), .A2(G169gat), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(G1348gat));
  INV_X1    g648(.A(G176gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n844), .A2(new_n850), .A3(new_n598), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n840), .A2(new_n677), .A3(new_n846), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(G1349gat));
  AOI21_X1  g652(.A(new_n300), .B1(new_n847), .B2(new_n577), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n577), .A2(new_n289), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n844), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g656(.A(new_n290), .B1(new_n847), .B2(new_n551), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT61), .Z(new_n859));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n290), .A3(new_n551), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1351gat));
  INV_X1    g660(.A(new_n840), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n790), .A2(new_n429), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT125), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n863), .A2(KEYINPUT125), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(G197gat), .B1(new_n867), .B2(new_n246), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n616), .A2(new_n679), .A3(new_n655), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n825), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n247), .A2(new_n236), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(G1352gat));
  OR3_X1    g672(.A1(new_n866), .A2(G204gat), .A3(new_n697), .ZN(new_n874));
  AND2_X1   g673(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n875));
  NOR2_X1   g674(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n871), .A2(new_n645), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G204gat), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n877), .B(new_n879), .C1(new_n875), .C2(new_n874), .ZN(G1353gat));
  NAND3_X1  g679(.A1(new_n867), .A2(new_n370), .A3(new_n577), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n871), .A2(new_n577), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT63), .B1(new_n882), .B2(G211gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(G1354gat));
  NOR2_X1   g684(.A1(new_n649), .A2(new_n369), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n869), .B(new_n886), .C1(new_n823), .C2(new_n824), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n866), .A2(new_n649), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(G218gat), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


