//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954;
  INV_X1    g000(.A(G127gat), .ZN(new_n202));
  INV_X1    g001(.A(G134gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G127gat), .A2(G134gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(G113gat), .A2(G120gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G113gat), .A2(G120gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(KEYINPUT72), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210));
  AND2_X1   g009(.A1(G113gat), .A2(G120gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G113gat), .A2(G120gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n206), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G127gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n202), .A2(KEYINPUT69), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n203), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n202), .A2(KEYINPUT69), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(G127gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(G134gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT70), .A3(new_n208), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(new_n211), .B2(new_n212), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n222), .A2(new_n227), .A3(KEYINPUT71), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT71), .B1(new_n222), .B2(new_n227), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n214), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT73), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  INV_X1    g032(.A(G176gat), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT23), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n235), .B1(G169gat), .B2(G176gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT66), .B(G169gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(KEYINPUT23), .A3(new_n234), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT23), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n236), .A2(new_n243), .A3(KEYINPUT25), .A4(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT67), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT26), .ZN(new_n251));
  NAND2_X1  g050(.A1(G169gat), .A2(G176gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT67), .A4(KEYINPUT26), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n240), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n253), .A2(new_n257), .A3(new_n240), .A4(new_n254), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT27), .B(G183gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT28), .B1(new_n260), .B2(G190gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n262));
  INV_X1    g061(.A(G190gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n256), .A2(new_n258), .A3(new_n261), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(KEYINPUT73), .B(new_n214), .C1(new_n228), .C2(new_n229), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n232), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n261), .A2(new_n258), .A3(new_n264), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n269), .A2(new_n256), .B1(new_n246), .B2(new_n248), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(new_n231), .A3(new_n230), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n274), .B(KEYINPUT64), .Z(new_n275));
  XOR2_X1   g074(.A(new_n275), .B(KEYINPUT65), .Z(new_n276));
  NOR3_X1   g075(.A1(new_n273), .A2(KEYINPUT34), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT76), .B1(new_n268), .B2(new_n271), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(new_n275), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(new_n272), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n281), .B2(KEYINPUT34), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n271), .A3(new_n276), .ZN(new_n284));
  XOR2_X1   g083(.A(G15gat), .B(G43gat), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(KEYINPUT74), .ZN(new_n286));
  XNOR2_X1  g085(.A(G71gat), .B(G99gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT33), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(KEYINPUT32), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT75), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n284), .A2(KEYINPUT75), .A3(KEYINPUT32), .A4(new_n289), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n284), .A2(KEYINPUT32), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT33), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n298), .A3(new_n288), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n294), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n295), .B1(new_n294), .B2(new_n299), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n283), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n294), .A2(new_n299), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT77), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n294), .A2(new_n295), .A3(new_n299), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n282), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307));
  INV_X1    g106(.A(G211gat), .ZN(new_n308));
  INV_X1    g107(.A(G218gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(KEYINPUT22), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G211gat), .B(G218gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n312), .B(new_n307), .C1(KEYINPUT22), .C2(new_n310), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT3), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G141gat), .B(G148gat), .Z(new_n319));
  XNOR2_X1  g118(.A(G155gat), .B(G162gat), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  INV_X1    g120(.A(G162gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT2), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n320), .B1(new_n319), .B2(new_n323), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OR3_X1    g126(.A1(new_n318), .A2(KEYINPUT85), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n317), .ZN(new_n331));
  INV_X1    g130(.A(new_n316), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(G228gat), .A2(G233gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT85), .B1(new_n318), .B2(new_n327), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n328), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT86), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G22gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n314), .A2(KEYINPUT83), .A3(new_n315), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT83), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n311), .A2(new_n340), .A3(new_n313), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n317), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT84), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n339), .A2(KEYINPUT84), .A3(new_n317), .A4(new_n341), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n329), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n327), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n346), .A2(new_n347), .B1(new_n332), .B2(new_n331), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n336), .B(new_n338), .C1(new_n348), .C2(new_n334), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n337), .A2(G22gat), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT31), .B(G50gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n349), .B2(new_n350), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n336), .B1(new_n348), .B2(new_n334), .ZN(new_n356));
  AND2_X1   g155(.A1(KEYINPUT87), .A2(G22gat), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n354), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(new_n356), .B2(new_n357), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n351), .A2(new_n355), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n302), .A2(new_n306), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT35), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n249), .B2(new_n265), .ZN(new_n367));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n366), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(KEYINPUT79), .B(new_n368), .C1(new_n270), .C2(KEYINPUT29), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n368), .B(KEYINPUT78), .Z(new_n372));
  NAND2_X1  g171(.A1(new_n266), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n316), .A4(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n367), .A2(new_n372), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n270), .A2(new_n368), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n332), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n365), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n374), .A2(new_n377), .A3(KEYINPUT30), .A4(new_n381), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n378), .B2(new_n382), .ZN(new_n386));
  AOI211_X1 g185(.A(KEYINPUT80), .B(new_n381), .C1(new_n374), .C2(new_n377), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n383), .B(new_n384), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n230), .A2(new_n347), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n214), .B(new_n327), .C1(new_n228), .C2(new_n229), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(KEYINPUT82), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n230), .A2(new_n394), .A3(new_n347), .ZN(new_n395));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT5), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n393), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n214), .ZN(new_n401));
  INV_X1    g200(.A(new_n229), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n222), .A2(new_n227), .A3(KEYINPUT71), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n327), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n392), .A2(KEYINPUT4), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT3), .B1(new_n325), .B2(new_n326), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n330), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n230), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n396), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT81), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n406), .A2(new_n407), .B1(new_n230), .B2(new_n410), .ZN(new_n415));
  INV_X1    g214(.A(new_n413), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n396), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n400), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G1gat), .B(G29gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT0), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n390), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n412), .A2(new_n413), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n416), .B1(new_n415), .B2(new_n396), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n423), .B(new_n399), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n399), .B1(new_n425), .B2(new_n426), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n430), .A2(new_n390), .A3(new_n422), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n389), .B(KEYINPUT89), .C1(new_n429), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n363), .A2(new_n364), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n302), .A2(new_n306), .A3(new_n362), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT35), .B1(new_n435), .B2(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n408), .A2(new_n411), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT39), .ZN(new_n439));
  INV_X1    g238(.A(new_n396), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT39), .B1(new_n415), .B2(new_n396), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n440), .B1(new_n393), .B2(new_n395), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n441), .B(new_n422), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT40), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n427), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n442), .A2(new_n443), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n441), .A2(new_n422), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT40), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n361), .B1(new_n450), .B2(new_n388), .ZN(new_n451));
  INV_X1    g250(.A(new_n431), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n430), .A2(new_n422), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n390), .A3(new_n427), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT88), .B(KEYINPUT37), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n382), .B1(new_n378), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n374), .B2(new_n377), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT38), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n378), .A2(new_n382), .ZN(new_n461));
  INV_X1    g260(.A(new_n457), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n375), .A2(new_n376), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n458), .B1(new_n463), .B2(new_n316), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n370), .A2(new_n371), .A3(new_n332), .A4(new_n373), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT38), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n461), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n452), .A2(new_n454), .A3(new_n460), .A4(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n389), .B1(new_n429), .B2(new_n431), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n451), .A2(new_n468), .B1(new_n469), .B2(new_n361), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n302), .A2(new_n306), .A3(KEYINPUT36), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT36), .B1(new_n302), .B2(new_n306), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n437), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G71gat), .ZN(new_n476));
  INV_X1    g275(.A(G78gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G71gat), .A2(G78gat), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G57gat), .B(G64gat), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n481), .A2(KEYINPUT94), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT9), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n481), .B2(KEYINPUT94), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n480), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G57gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT95), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT95), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G57gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n490), .A3(G64gat), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n487), .A2(G64gat), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT96), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(KEYINPUT96), .A3(new_n492), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n479), .B1(new_n478), .B2(new_n483), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n486), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT98), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT98), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n486), .B(new_n499), .C1(new_n493), .C2(new_n496), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT21), .ZN(new_n502));
  XOR2_X1   g301(.A(G15gat), .B(G22gat), .Z(new_n503));
  OR2_X1    g302(.A1(new_n503), .A2(KEYINPUT16), .ZN(new_n504));
  INV_X1    g303(.A(G1gat), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n503), .B2(KEYINPUT91), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(G1gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n504), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G8gat), .ZN(new_n511));
  INV_X1    g310(.A(G8gat), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n504), .A2(new_n506), .A3(new_n512), .A4(new_n509), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n502), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n496), .A2(new_n493), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT21), .B1(new_n518), .B2(new_n486), .ZN(new_n519));
  AND2_X1   g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G127gat), .B(G155gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(KEYINPUT20), .Z(new_n523));
  XNOR2_X1  g322(.A(new_n521), .B(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(G183gat), .B(G211gat), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n523), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n521), .B(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n525), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n517), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n517), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n525), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n524), .A2(new_n526), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT102), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT101), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT7), .ZN(new_n539));
  INV_X1    g338(.A(G85gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(G92gat), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n544));
  AND2_X1   g343(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(KEYINPUT100), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT100), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(G99gat), .A3(G106gat), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n543), .A2(new_n546), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G99gat), .B(G106gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n538), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n551), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n539), .A2(new_n540), .A3(G92gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n544), .A2(new_n545), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n555), .B(new_n553), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n555), .B1(new_n557), .B2(new_n556), .ZN(new_n561));
  INV_X1    g360(.A(new_n553), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n561), .A2(new_n538), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n537), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(new_n538), .A3(new_n558), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n567), .A3(KEYINPUT102), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G29gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n570), .A2(KEYINPUT14), .ZN(new_n572));
  INV_X1    g371(.A(G36gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n570), .B2(KEYINPUT14), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n571), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n575), .A2(KEYINPUT15), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(KEYINPUT15), .ZN(new_n577));
  XNOR2_X1  g376(.A(G43gat), .B(G50gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(KEYINPUT17), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n564), .A2(new_n582), .A3(new_n568), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT103), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n588), .A2(KEYINPUT103), .A3(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n589), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT99), .Z(new_n598));
  AND2_X1   g397(.A1(new_n590), .A2(new_n597), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n594), .A2(new_n598), .B1(new_n593), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n536), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n602));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  AND4_X1   g403(.A1(new_n511), .A2(new_n513), .A3(new_n579), .A4(new_n580), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n511), .A2(new_n513), .B1(new_n579), .B2(new_n580), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT93), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n584), .A2(new_n514), .A3(new_n581), .ZN(new_n609));
  INV_X1    g408(.A(new_n606), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n603), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G169gat), .B(G197gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n608), .A2(new_n613), .A3(new_n614), .A4(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n565), .A2(new_n497), .A3(new_n567), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n518), .A2(new_n486), .A3(new_n558), .A4(new_n566), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n627), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT106), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n630), .A2(new_n627), .A3(new_n632), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI211_X1 g436(.A(KEYINPUT105), .B(new_n631), .C1(new_n628), .C2(new_n629), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT106), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n498), .A2(KEYINPUT10), .A3(new_n500), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n645), .B1(new_n569), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n631), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT104), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n650), .A3(new_n631), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n640), .A2(new_n643), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n643), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n636), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n501), .A2(KEYINPUT10), .A3(new_n568), .A4(new_n564), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n632), .B1(new_n655), .B2(new_n645), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n601), .A2(new_n626), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n475), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n429), .A2(new_n431), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n505), .ZN(G1324gat));
  INV_X1    g463(.A(new_n660), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n512), .B1(new_n665), .B2(new_n388), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT16), .B(G8gat), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n660), .A2(new_n389), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT42), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(KEYINPUT42), .B2(new_n668), .ZN(G1325gat));
  NOR3_X1   g469(.A1(new_n300), .A2(new_n283), .A3(new_n301), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n282), .B1(new_n304), .B2(new_n305), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n660), .A2(G15gat), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT36), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n671), .B2(new_n672), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n471), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n665), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n675), .B1(G15gat), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT107), .Z(G1326gat));
  NOR2_X1   g481(.A1(new_n660), .A2(new_n362), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n436), .A2(new_n434), .B1(new_n678), .B2(new_n470), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n687), .B2(new_n600), .ZN(new_n688));
  INV_X1    g487(.A(new_n600), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n475), .A2(KEYINPUT44), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n536), .A2(new_n626), .A3(new_n658), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n662), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n600), .B1(new_n437), .B2(new_n474), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n695), .A2(new_n570), .A3(new_n661), .A4(new_n692), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n697), .B2(new_n699), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n694), .B1(new_n700), .B2(new_n701), .ZN(G1328gat));
  NAND2_X1  g501(.A1(new_n695), .A2(new_n692), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(G36gat), .A3(new_n389), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n693), .B2(new_n389), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1329gat));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n679), .A3(new_n692), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G43gat), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n703), .A2(G43gat), .A3(new_n674), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT47), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n709), .B(new_n710), .C1(new_n712), .C2(KEYINPUT47), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1330gat));
  INV_X1    g515(.A(G50gat), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n688), .A2(new_n690), .A3(new_n361), .A4(new_n692), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(KEYINPUT112), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT112), .B2(new_n718), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n695), .A2(KEYINPUT110), .A3(new_n692), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n722), .A2(new_n717), .A3(new_n361), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n720), .A2(KEYINPUT48), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n718), .A2(G50gat), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT48), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(KEYINPUT111), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  AOI211_X1 g528(.A(new_n729), .B(KEYINPUT48), .C1(new_n724), .C2(new_n726), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n725), .B1(new_n728), .B2(new_n730), .ZN(G1331gat));
  INV_X1    g530(.A(new_n658), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n601), .A2(new_n625), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n475), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n662), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n488), .A2(new_n490), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1332gat));
  NOR2_X1   g536(.A1(new_n734), .A2(new_n389), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  AND2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n738), .B2(new_n739), .ZN(G1333gat));
  NOR3_X1   g541(.A1(new_n734), .A2(G71gat), .A3(new_n674), .ZN(new_n743));
  INV_X1    g542(.A(new_n734), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n679), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n743), .B1(G71gat), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n734), .A2(new_n362), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n477), .ZN(G1335gat));
  NOR2_X1   g548(.A1(new_n536), .A2(new_n625), .ZN(new_n750));
  AND4_X1   g549(.A1(KEYINPUT51), .A2(new_n475), .A3(new_n689), .A4(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT51), .B1(new_n695), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n754), .A2(new_n540), .A3(new_n661), .A4(new_n658), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n536), .A2(new_n625), .A3(new_n732), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n691), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(new_n661), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n758), .B2(new_n540), .ZN(G1336gat));
  NAND3_X1  g558(.A1(new_n691), .A2(new_n388), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n732), .A2(new_n389), .A3(G92gat), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT113), .Z(new_n763));
  NAND2_X1  g562(.A1(new_n754), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT52), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n761), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1337gat));
  AND2_X1   g568(.A1(new_n757), .A2(new_n679), .ZN(new_n770));
  INV_X1    g569(.A(G99gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n673), .A2(new_n771), .A3(new_n658), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n770), .A2(new_n771), .B1(new_n753), .B2(new_n772), .ZN(G1338gat));
  NAND4_X1  g572(.A1(new_n688), .A2(new_n690), .A3(new_n361), .A4(new_n756), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G106gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n362), .A2(new_n732), .A3(G106gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n751), .B2(new_n752), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n774), .A2(KEYINPUT114), .A3(G106gat), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT115), .B(new_n778), .C1(new_n751), .C2(new_n752), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n777), .A2(new_n781), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT53), .ZN(new_n785));
  INV_X1    g584(.A(G106gat), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n774), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n787), .B2(new_n774), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n790), .A3(new_n779), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n791), .ZN(G1339gat));
  INV_X1    g591(.A(new_n536), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n645), .B(new_n632), .C1(new_n569), .C2(new_n646), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(KEYINPUT54), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n649), .A2(new_n796), .A3(new_n651), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n643), .B1(new_n656), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(KEYINPUT55), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n652), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT55), .B1(new_n797), .B2(new_n799), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n794), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n797), .A2(new_n799), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n806), .A2(KEYINPUT118), .A3(new_n652), .A4(new_n800), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n803), .A2(new_n625), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n603), .B1(new_n609), .B2(new_n610), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n605), .A2(new_n606), .A3(new_n604), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n620), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n624), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n732), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n689), .B1(new_n808), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n812), .B(KEYINPUT119), .ZN(new_n816));
  AND4_X1   g615(.A1(new_n689), .A2(new_n803), .A3(new_n816), .A4(new_n807), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n793), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n536), .A2(new_n600), .A3(new_n626), .A4(new_n732), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n362), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n661), .A2(new_n389), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n674), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n625), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n822), .A2(KEYINPUT120), .A3(new_n362), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT120), .B1(new_n822), .B2(new_n362), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n829), .A2(new_n830), .A3(new_n826), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n625), .A2(G113gat), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(G1340gat));
  INV_X1    g632(.A(G120gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n827), .A2(new_n834), .A3(new_n658), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n658), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n836), .A2(KEYINPUT121), .A3(G120gat), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT121), .B1(new_n836), .B2(G120gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(G1341gat));
  NAND3_X1  g638(.A1(new_n827), .A2(new_n202), .A3(new_n536), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n831), .A2(new_n536), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n202), .ZN(G1342gat));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n600), .A2(G134gat), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n822), .A2(new_n362), .A3(new_n825), .A4(new_n844), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT56), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n831), .A2(new_n689), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n843), .B(new_n847), .C1(new_n848), .C2(new_n203), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n203), .B1(new_n831), .B2(new_n689), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT122), .B1(new_n850), .B2(new_n846), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(G1343gat));
  NOR2_X1   g651(.A1(new_n679), .A2(new_n824), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n802), .B(KEYINPUT123), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n626), .A2(new_n801), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n813), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n689), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n793), .B1(new_n858), .B2(new_n817), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n854), .B(new_n362), .C1(new_n859), .C2(new_n821), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(new_n822), .B2(new_n361), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n853), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G141gat), .B1(new_n862), .B2(new_n626), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n362), .B1(new_n818), .B2(new_n821), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n853), .ZN(new_n865));
  INV_X1    g664(.A(G141gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n866), .A3(new_n625), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT58), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n863), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1344gat));
  INV_X1    g671(.A(G148gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n865), .A2(new_n873), .A3(new_n658), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n862), .A2(new_n732), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(KEYINPUT59), .A3(new_n873), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n853), .B(KEYINPUT124), .ZN(new_n878));
  INV_X1    g677(.A(new_n819), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n806), .A2(new_n652), .A3(new_n800), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n689), .A2(new_n816), .ZN(new_n881));
  OAI22_X1  g680(.A1(new_n857), .A2(new_n689), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n879), .B1(new_n882), .B2(new_n793), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n854), .B1(new_n883), .B2(new_n362), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n854), .B(new_n362), .C1(new_n818), .C2(new_n821), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n864), .A2(new_n886), .A3(KEYINPUT57), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n658), .B(new_n878), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n877), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n874), .B1(new_n876), .B2(new_n890), .ZN(G1345gat));
  OAI21_X1  g690(.A(G155gat), .B1(new_n862), .B2(new_n793), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n865), .A2(new_n321), .A3(new_n536), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n862), .B2(new_n600), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n865), .A2(new_n322), .A3(new_n689), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n661), .A2(new_n389), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n674), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n829), .A2(new_n830), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n626), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n661), .B1(new_n818), .B2(new_n821), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n905), .A2(new_n388), .A3(new_n363), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n237), .A3(new_n625), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n829), .A2(new_n830), .A3(new_n901), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n233), .B1(new_n909), .B2(new_n625), .ZN(new_n910));
  INV_X1    g709(.A(new_n907), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT126), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n912), .ZN(G1348gat));
  OAI21_X1  g712(.A(G176gat), .B1(new_n902), .B2(new_n732), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n906), .A2(new_n234), .A3(new_n658), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1349gat));
  OAI21_X1  g715(.A(G183gat), .B1(new_n902), .B2(new_n793), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n906), .A2(new_n259), .A3(new_n536), .ZN(new_n918));
  XNOR2_X1  g717(.A(KEYINPUT127), .B(KEYINPUT60), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n919), .ZN(new_n921));
  INV_X1    g720(.A(G183gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n922), .B1(new_n909), .B2(new_n536), .ZN(new_n923));
  INV_X1    g722(.A(new_n918), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n920), .A2(new_n925), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n906), .A2(new_n263), .A3(new_n689), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n909), .A2(new_n689), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(G190gat), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT61), .B(new_n263), .C1(new_n909), .C2(new_n689), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(G1351gat));
  NOR3_X1   g731(.A1(new_n679), .A2(new_n362), .A3(new_n389), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n905), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n625), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n679), .A2(new_n899), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n887), .ZN(new_n938));
  INV_X1    g737(.A(new_n888), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n625), .A2(G197gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n935), .B1(new_n940), .B2(new_n941), .ZN(G1352gat));
  INV_X1    g741(.A(G204gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n934), .A2(new_n943), .A3(new_n658), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT62), .Z(new_n945));
  AOI211_X1 g744(.A(new_n732), .B(new_n937), .C1(new_n938), .C2(new_n939), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n943), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n934), .A2(new_n308), .A3(new_n536), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n536), .B(new_n936), .C1(new_n887), .C2(new_n888), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1354gat));
  NAND3_X1  g751(.A1(new_n934), .A2(new_n309), .A3(new_n689), .ZN(new_n953));
  AOI211_X1 g752(.A(new_n600), .B(new_n937), .C1(new_n938), .C2(new_n939), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n309), .ZN(G1355gat));
endmodule


