//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n218), .B1(new_n212), .B2(new_n211), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G226), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(new_n232), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  AOI21_X1  g0044(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT3), .B(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G1698), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  AND2_X1   g0049(.A1(new_n249), .A2(G223), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G222), .ZN(new_n253));
  INV_X1    g0053(.A(G77), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n246), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n245), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT66), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n260), .B(new_n206), .C1(G41), .C2(G45), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(G274), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n259), .A2(new_n263), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(G226), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n256), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G200), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT68), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n213), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G50), .B2(new_n273), .ZN(new_n279));
  INV_X1    g0079(.A(new_n276), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n207), .A2(G33), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n280), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT9), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT10), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n256), .A2(G190), .A3(new_n268), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n270), .A2(new_n289), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT71), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n270), .A2(new_n289), .A3(new_n291), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT72), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(KEYINPUT72), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n269), .A2(G169), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n269), .ZN(new_n301));
  INV_X1    g0101(.A(new_n287), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT75), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G58), .A2(G68), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n215), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n305), .B1(new_n307), .B2(G20), .ZN(new_n308));
  INV_X1    g0108(.A(new_n306), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n305), .B(G20), .C1(new_n309), .C2(new_n201), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n284), .A2(G159), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n257), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT74), .A2(G33), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(KEYINPUT3), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G33), .ZN(new_n319));
  AOI21_X1  g0119(.A(G20), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT7), .ZN(new_n321));
  OAI21_X1  g0121(.A(G68), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI211_X1 g0122(.A(KEYINPUT7), .B(G20), .C1(new_n317), .C2(new_n319), .ZN(new_n323));
  OAI211_X1 g0123(.A(KEYINPUT16), .B(new_n313), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT16), .ZN(new_n325));
  INV_X1    g0125(.A(G68), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n321), .A2(G20), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT3), .B1(new_n315), .B2(new_n316), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n327), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n321), .B1(new_n246), .B2(G20), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(G20), .B1(new_n309), .B2(new_n201), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT75), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(new_n310), .A3(new_n311), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n325), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n324), .A2(new_n337), .A3(new_n276), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n281), .B1(new_n206), .B2(G20), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(new_n277), .B1(new_n274), .B2(new_n281), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n259), .A2(G274), .A3(new_n261), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n264), .B1(new_n267), .B2(G232), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n251), .A2(G223), .ZN(new_n344));
  INV_X1    g0144(.A(G226), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(new_n251), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n317), .A2(new_n346), .A3(new_n319), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G87), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n342), .B(new_n343), .C1(new_n349), .C2(new_n259), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n259), .B1(new_n347), .B2(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n259), .A2(new_n263), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n262), .A2(new_n265), .B1(new_n353), .B2(new_n231), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n351), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n338), .A2(new_n340), .A3(new_n356), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n357), .A2(KEYINPUT17), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT76), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n338), .A2(new_n356), .A3(KEYINPUT76), .A4(new_n340), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT17), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n338), .A2(new_n340), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n352), .A2(new_n354), .A3(G179), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n342), .B1(new_n349), .B2(new_n259), .ZN(new_n367));
  INV_X1    g0167(.A(G169), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n249), .A2(G238), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n246), .A2(G232), .A3(new_n251), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n246), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n245), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n266), .B1(G244), .B2(new_n267), .ZN(new_n379));
  AOI21_X1  g0179(.A(G169), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT70), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n379), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(G179), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n378), .A2(KEYINPUT70), .A3(new_n300), .A4(new_n379), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n281), .A2(G20), .A3(G33), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT15), .B(G87), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n386), .A2(new_n282), .B1(new_n207), .B2(new_n254), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n276), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  XOR2_X1   g0188(.A(new_n388), .B(KEYINPUT69), .Z(new_n389));
  AOI21_X1  g0189(.A(new_n254), .B1(new_n206), .B2(G20), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n277), .A2(new_n390), .B1(new_n254), .B2(new_n274), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n392), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n382), .A2(G190), .ZN(new_n397));
  AOI21_X1  g0197(.A(G200), .B1(new_n378), .B2(new_n379), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT13), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n246), .A2(G232), .A3(G1698), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(new_n252), .C2(new_n345), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n245), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n341), .A2(new_n264), .B1(new_n267), .B2(G238), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n402), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT73), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n409), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n406), .A2(new_n402), .A3(new_n407), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n410), .A2(G179), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(G169), .C1(new_n412), .C2(new_n408), .ZN(new_n416));
  OAI21_X1  g0216(.A(G169), .B1(new_n412), .B2(new_n408), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT14), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G13), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n420), .A2(G1), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(G20), .A3(new_n326), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT12), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n277), .B(G68), .C1(G1), .C2(new_n207), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n284), .A2(G50), .B1(G20), .B2(new_n326), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n254), .B2(new_n282), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(KEYINPUT11), .A3(new_n276), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT11), .B1(new_n426), .B2(new_n276), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n419), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n412), .A2(new_n408), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n430), .B1(new_n432), .B2(G200), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n343), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n401), .A2(new_n436), .ZN(new_n437));
  OR3_X1    g0237(.A1(new_n304), .A2(new_n373), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G116), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n275), .A2(new_n213), .B1(G20), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G283), .ZN(new_n441));
  INV_X1    g0241(.A(G97), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(new_n207), .C1(G33), .C2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(KEYINPUT20), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT83), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT20), .B1(new_n440), .B2(new_n443), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT83), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n440), .A2(new_n448), .A3(new_n443), .A4(KEYINPUT20), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n207), .A2(G116), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(new_n421), .A3(KEYINPUT82), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT82), .B1(new_n451), .B2(new_n421), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n206), .A2(G33), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n273), .A2(new_n455), .A3(new_n213), .A4(new_n275), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n453), .A2(new_n454), .B1(new_n439), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n450), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n206), .A2(G45), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT5), .B(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n245), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n461), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n259), .A2(G274), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n463), .A2(G270), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G264), .A2(G1698), .ZN(new_n468));
  INV_X1    g0268(.A(G257), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(G1698), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n317), .A2(new_n319), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n319), .A2(new_n329), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G303), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n245), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n459), .A2(new_n476), .A3(KEYINPUT21), .A4(G169), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n462), .A2(new_n259), .A3(G274), .A4(new_n461), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n464), .A2(new_n259), .ZN(new_n479));
  INV_X1    g0279(.A(G270), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n259), .B1(new_n471), .B2(new_n473), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n459), .A2(new_n483), .A3(G179), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n446), .B1(KEYINPUT83), .B2(new_n444), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n457), .B1(new_n486), .B2(new_n449), .ZN(new_n487));
  AOI21_X1  g0287(.A(G200), .B1(new_n467), .B2(new_n475), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n481), .A2(new_n482), .A3(G190), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT21), .ZN(new_n491));
  OAI21_X1  g0291(.A(G169), .B1(new_n481), .B2(new_n482), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n485), .A2(KEYINPUT84), .A3(new_n490), .A4(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n490), .A2(new_n493), .A3(new_n477), .A4(new_n484), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT84), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G250), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(KEYINPUT79), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n461), .B1(new_n500), .B2(G274), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n460), .A2(KEYINPUT79), .A3(G250), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n245), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G244), .A2(G1698), .ZN(new_n505));
  INV_X1    g0305(.A(G238), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(G1698), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n317), .A2(new_n319), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n315), .A2(new_n316), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G116), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n504), .B1(new_n511), .B2(new_n259), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G200), .ZN(new_n513));
  NOR2_X1   g0313(.A1(G87), .A2(G97), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(new_n376), .B1(new_n404), .B2(new_n207), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT19), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n207), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n515), .A2(new_n516), .B1(new_n404), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n317), .A2(new_n207), .A3(G68), .A4(new_n319), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n280), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n386), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n521), .A2(new_n273), .ZN(new_n522));
  INV_X1    g0322(.A(G87), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n456), .A2(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n259), .B1(new_n508), .B2(new_n510), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n503), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G190), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n513), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT80), .ZN(new_n530));
  NOR4_X1   g0330(.A1(new_n526), .A2(new_n503), .A3(new_n530), .A4(G179), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n512), .B2(new_n368), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n512), .A2(G179), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT81), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n518), .A2(new_n519), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n522), .B1(new_n537), .B2(new_n276), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n456), .A2(new_n386), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NOR4_X1   g0341(.A1(new_n520), .A2(KEYINPUT81), .A3(new_n522), .A4(new_n539), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n529), .B1(new_n535), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n274), .A2(new_n442), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n545), .A2(KEYINPUT78), .ZN(new_n546));
  INV_X1    g0346(.A(new_n456), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(KEYINPUT78), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g0350(.A(G97), .B(G107), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT77), .ZN(new_n554));
  NAND2_X1  g0354(.A1(KEYINPUT6), .A2(G97), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n554), .B1(new_n555), .B2(G107), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n376), .A2(KEYINPUT77), .A3(KEYINPUT6), .A4(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n331), .A2(new_n332), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(new_n561), .B2(new_n376), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n550), .B1(new_n562), .B2(new_n276), .ZN(new_n563));
  INV_X1    g0363(.A(new_n319), .ZN(new_n564));
  AND2_X1   g0364(.A1(KEYINPUT74), .A2(G33), .ZN(new_n565));
  NOR2_X1   g0365(.A1(KEYINPUT74), .A2(G33), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n567), .B2(KEYINPUT3), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n251), .A2(G244), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT4), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n319), .A2(new_n329), .A3(G250), .A4(G1698), .ZN(new_n572));
  AND2_X1   g0372(.A1(KEYINPUT4), .A2(G244), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n319), .A2(new_n329), .A3(new_n573), .A4(new_n251), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n574), .A3(new_n441), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n245), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n478), .B1(new_n479), .B2(new_n469), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(G200), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n317), .A2(new_n319), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n569), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n572), .A2(new_n574), .A3(new_n441), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n259), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n584), .A2(G190), .A3(new_n577), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n563), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n559), .A2(G20), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n284), .A2(G77), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n376), .B1(new_n331), .B2(new_n332), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n276), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n550), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n368), .B1(new_n576), .B2(new_n578), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n584), .A2(new_n300), .A3(new_n577), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n586), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n544), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G257), .A2(G1698), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n499), .B2(G1698), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n317), .A2(new_n319), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n509), .A2(G294), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT86), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT86), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n605), .A3(new_n602), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n245), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n463), .A2(G264), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n607), .A2(G179), .A3(new_n478), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n245), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n605), .B1(new_n601), .B2(new_n602), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n478), .B(new_n608), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n609), .A2(KEYINPUT87), .B1(new_n612), .B2(G169), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n612), .A2(KEYINPUT87), .A3(G169), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT22), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n523), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n317), .A2(new_n207), .A3(new_n319), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n207), .A2(G87), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n615), .B1(new_n472), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n376), .A2(G20), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT23), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n509), .A2(new_n207), .A3(G116), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n617), .A2(new_n619), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n624), .A2(KEYINPUT24), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT24), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(KEYINPUT85), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n626), .A2(KEYINPUT85), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n280), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n421), .A2(G20), .A3(new_n376), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n630), .A2(KEYINPUT25), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(KEYINPUT25), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n631), .B(new_n632), .C1(new_n376), .C2(new_n456), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n613), .A2(new_n614), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(KEYINPUT85), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(KEYINPUT24), .B2(new_n624), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n626), .A2(KEYINPUT85), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n276), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n612), .A2(new_n351), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(G190), .B2(new_n612), .ZN(new_n640));
  INV_X1    g0440(.A(new_n633), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n498), .A2(new_n598), .A3(new_n634), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n438), .A2(new_n643), .ZN(G372));
  NAND2_X1  g0444(.A1(new_n395), .A2(new_n435), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n431), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n364), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n372), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n298), .B1(new_n302), .B2(new_n301), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n485), .A2(new_n493), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n634), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT88), .ZN(new_n652));
  OAI21_X1  g0452(.A(G169), .B1(new_n584), .B2(new_n577), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n576), .A2(G179), .A3(new_n578), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n653), .A2(new_n654), .B1(new_n591), .B2(new_n592), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n584), .A2(new_n577), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n343), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n576), .A2(new_n578), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n351), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n655), .B1(new_n563), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n642), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n527), .A2(new_n300), .ZN(new_n663));
  OAI221_X1 g0463(.A(new_n663), .B1(G169), .B2(new_n527), .C1(new_n541), .C2(new_n542), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n662), .A2(new_n529), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n651), .A2(KEYINPUT88), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n652), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(new_n655), .A3(new_n529), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT26), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n513), .A2(new_n525), .A3(new_n528), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n541), .A2(new_n542), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT80), .B1(new_n527), .B2(G169), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n531), .B1(new_n672), .B2(new_n663), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n670), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n655), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n669), .A2(new_n676), .A3(new_n664), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n667), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n649), .B1(new_n438), .B2(new_n679), .ZN(G369));
  NAND2_X1  g0480(.A1(new_n206), .A2(G13), .ZN(new_n681));
  OR3_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .A3(G20), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT27), .B1(new_n681), .B2(G20), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n487), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n650), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n498), .B2(new_n688), .ZN(new_n690));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n634), .A2(new_n687), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n686), .B1(new_n629), .B2(new_n633), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n634), .A2(new_n642), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n650), .A2(new_n686), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(new_n696), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n634), .B2(new_n686), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n698), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n210), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n514), .A2(new_n376), .A3(new_n439), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n704), .A2(new_n705), .A3(new_n206), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n217), .B2(new_n704), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  NAND2_X1  g0508(.A1(new_n662), .A2(new_n529), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n651), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n668), .A2(KEYINPUT26), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n711), .B(new_n664), .C1(new_n675), .C2(KEYINPUT26), .ZN(new_n712));
  OAI211_X1 g0512(.A(KEYINPUT29), .B(new_n687), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n686), .B1(new_n667), .B2(new_n677), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(KEYINPUT29), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n656), .A2(G179), .A3(new_n483), .A4(new_n527), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n607), .A2(new_n608), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n476), .A2(new_n512), .A3(new_n300), .ZN(new_n720));
  INV_X1    g0520(.A(new_n718), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(KEYINPUT30), .A4(new_n656), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n483), .A2(new_n527), .A3(G179), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n612), .A3(new_n658), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n719), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n726), .B(KEYINPUT89), .Z(new_n727));
  NAND4_X1  g0527(.A1(new_n634), .A2(new_n642), .A3(new_n661), .A4(new_n674), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n495), .B(KEYINPUT84), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT31), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n719), .A2(new_n722), .A3(new_n731), .A4(new_n724), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n686), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G330), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n715), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n708), .B1(new_n737), .B2(G1), .ZN(G364));
  INV_X1    g0538(.A(new_n704), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n420), .A2(G20), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G45), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n739), .A2(G1), .A3(new_n741), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n690), .A2(new_n691), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n743), .B2(new_n692), .ZN(new_n744));
  INV_X1    g0544(.A(new_n742), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n690), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n703), .A2(new_n472), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n750), .A2(G355), .B1(new_n439), .B2(new_n703), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n217), .A2(G45), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n240), .B2(G45), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n703), .A2(new_n568), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n751), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n213), .B1(G20), .B2(new_n368), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n300), .A2(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n207), .A2(G190), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n351), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G77), .A2(new_n763), .B1(new_n766), .B2(G107), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n207), .A2(new_n343), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n764), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n523), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n761), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G159), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT91), .B(KEYINPUT32), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n768), .A2(new_n760), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n472), .B1(new_n778), .B2(G58), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n207), .B1(new_n771), .B2(G190), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n776), .B(new_n779), .C1(new_n442), .C2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n207), .A2(new_n300), .A3(new_n351), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT90), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(KEYINPUT90), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n783), .A2(G190), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n770), .B(new_n781), .C1(G50), .C2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n783), .A2(new_n343), .A3(new_n784), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT92), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G68), .ZN(new_n793));
  INV_X1    g0593(.A(new_n780), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n786), .A2(G326), .B1(G294), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT93), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n472), .B1(new_n762), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n772), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G283), .A2(new_n766), .B1(new_n800), .B2(G329), .ZN(new_n801));
  INV_X1    g0601(.A(G303), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(new_n802), .B2(new_n769), .C1(new_n803), .C2(new_n777), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n797), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT94), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n792), .A2(new_n807), .B1(new_n795), .B2(new_n796), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n787), .A2(new_n793), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n757), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n759), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n745), .B1(new_n749), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n744), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT95), .Z(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NOR2_X1   g0615(.A1(new_n394), .A2(new_n686), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n392), .A2(new_n686), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n399), .A2(new_n817), .B1(new_n383), .B2(new_n393), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n714), .B(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n736), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n745), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n822), .B2(new_n821), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n786), .A2(G137), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G143), .A2(new_n778), .B1(new_n763), .B2(G159), .ZN(new_n826));
  INV_X1    g0626(.A(new_n792), .ZN(new_n827));
  INV_X1    g0627(.A(G150), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n825), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT34), .Z(new_n830));
  INV_X1    g0630(.A(new_n769), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G50), .A2(new_n831), .B1(new_n766), .B2(G68), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n772), .ZN(new_n834));
  INV_X1    g0634(.A(G58), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n568), .B1(new_n835), .B2(new_n780), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n830), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n785), .A2(new_n802), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n769), .A2(new_n376), .B1(new_n762), .B2(new_n439), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n246), .B(new_n839), .C1(G294), .C2(new_n778), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n765), .A2(new_n523), .B1(new_n772), .B2(new_n798), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT96), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n840), .B(new_n842), .C1(new_n442), .C2(new_n780), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n838), .B(new_n843), .C1(G283), .C2(new_n792), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n757), .B1(new_n837), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n757), .A2(new_n746), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n742), .B1(new_n254), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n845), .B(new_n847), .C1(new_n819), .C2(new_n747), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n824), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n431), .A2(new_n686), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n324), .A2(new_n276), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT7), .B1(new_n568), .B2(G20), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n320), .A2(new_n321), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n853), .A2(G68), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT16), .B1(new_n855), .B2(new_n313), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n340), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT98), .ZN(new_n858));
  INV_X1    g0658(.A(new_n684), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT98), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n860), .B(new_n340), .C1(new_n852), .C2(new_n856), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n858), .A2(new_n369), .A3(new_n861), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n862), .A2(new_n863), .A3(new_n360), .A4(new_n361), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n365), .A2(new_n859), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n370), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(new_n362), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT99), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n862), .B1(new_n364), .B2(new_n372), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n869), .B1(new_n864), .B2(KEYINPUT37), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT99), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n872), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n370), .A2(new_n866), .A3(new_n357), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n869), .B1(KEYINPUT37), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n866), .B1(new_n364), .B2(new_n372), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n877), .A2(new_n878), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n872), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n872), .B2(new_n876), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT39), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n884), .B1(new_n887), .B2(KEYINPUT100), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n877), .A2(new_n878), .A3(new_n883), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT100), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n851), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n372), .A2(new_n859), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n430), .A2(new_n686), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n431), .A2(new_n435), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n419), .A2(new_n430), .A3(new_n686), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT97), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n419), .A2(KEYINPUT97), .A3(new_n430), .A4(new_n686), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n895), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n714), .A2(new_n819), .ZN(new_n902));
  INV_X1    g0702(.A(new_n816), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n865), .A2(new_n875), .A3(new_n870), .ZN(new_n905));
  INV_X1    g0705(.A(new_n873), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n874), .A2(new_n875), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n879), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n877), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n893), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n892), .A2(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n715), .A2(new_n438), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n649), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n912), .B(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n733), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n643), .B2(KEYINPUT31), .ZN(new_n917));
  INV_X1    g0717(.A(new_n726), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n819), .B(new_n900), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT101), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n734), .A2(new_n726), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(KEYINPUT40), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n922), .A2(new_n819), .A3(new_n900), .A4(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n885), .A2(new_n886), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n919), .B1(new_n877), .B2(new_n883), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n925), .A2(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n438), .B1(new_n734), .B2(new_n726), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n929), .B(new_n930), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(G330), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n915), .A2(new_n932), .B1(new_n206), .B2(new_n740), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT102), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n915), .A2(new_n932), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(G116), .B(new_n214), .C1(new_n559), .C2(KEYINPUT35), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(KEYINPUT35), .B2(new_n559), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT36), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT36), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n306), .A2(G77), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n216), .A2(new_n943), .B1(G50), .B2(new_n326), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(G1), .A3(new_n420), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n938), .A2(new_n941), .A3(new_n942), .A4(new_n945), .ZN(G367));
  NAND2_X1  g0746(.A1(new_n664), .A2(new_n529), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n525), .A2(new_n687), .ZN(new_n948));
  MUX2_X1   g0748(.A(new_n947), .B(new_n664), .S(new_n948), .Z(new_n949));
  INV_X1    g0749(.A(KEYINPUT43), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n661), .B1(new_n563), .B2(new_n687), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n596), .B1(new_n952), .B2(new_n634), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n687), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n700), .A2(new_n952), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT42), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n958), .A2(KEYINPUT103), .B1(KEYINPUT42), .B2(new_n955), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n958), .A2(KEYINPUT103), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n951), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n949), .A2(new_n950), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n961), .B(new_n962), .Z(new_n963));
  NAND2_X1  g0763(.A1(new_n655), .A2(new_n686), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n952), .A2(new_n964), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n693), .A2(new_n697), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n963), .B(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n704), .B(KEYINPUT41), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n697), .A2(new_n699), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n700), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n692), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n737), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT104), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(KEYINPUT104), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n701), .A2(new_n965), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT44), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n701), .A2(new_n965), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n698), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n968), .B1(new_n982), .B2(new_n737), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n741), .A2(G1), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n967), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(KEYINPUT105), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT105), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n967), .B(new_n987), .C1(new_n983), .C2(new_n984), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n236), .A2(new_n755), .ZN(new_n990));
  INV_X1    g0790(.A(new_n758), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n703), .B2(new_n521), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n831), .A2(G116), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT46), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n568), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n995), .B2(new_n994), .C1(new_n376), .C2(new_n780), .ZN(new_n997));
  INV_X1    g0797(.A(G283), .ZN(new_n998));
  INV_X1    g0798(.A(G317), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n762), .A2(new_n998), .B1(new_n772), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n766), .A2(G97), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n802), .B2(new_n777), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n997), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(G294), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n827), .C1(new_n798), .C2(new_n785), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n246), .B1(new_n780), .B2(new_n326), .C1(new_n835), .C2(new_n769), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(KEYINPUT106), .B(G137), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n777), .A2(new_n828), .B1(new_n772), .B2(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n202), .A2(new_n762), .B1(new_n765), .B2(new_n254), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(G143), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n1011), .B2(new_n785), .C1(new_n827), .C2(new_n773), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1005), .A2(KEYINPUT47), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n757), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT47), .B1(new_n1005), .B2(new_n1012), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n745), .B1(new_n990), .B2(new_n993), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n949), .A2(new_n748), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n989), .A2(new_n1019), .ZN(G387));
  NAND2_X1  g0820(.A1(new_n750), .A2(new_n705), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(G107), .B2(new_n210), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n232), .A2(G45), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n281), .A2(G50), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT50), .ZN(new_n1025));
  AOI211_X1 g0825(.A(G45), .B(new_n705), .C1(G68), .C2(G77), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n755), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1022), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n745), .B1(new_n1028), .B2(new_n991), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n831), .A2(G77), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n800), .A2(G150), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1030), .A2(new_n1001), .A3(new_n1031), .A4(new_n568), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT107), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G50), .A2(new_n778), .B1(new_n763), .B2(G68), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n386), .B2(new_n780), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G159), .B2(new_n786), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1033), .B(new_n1036), .C1(new_n827), .C2(new_n281), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G116), .A2(new_n766), .B1(new_n800), .B2(G326), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n769), .A2(new_n1004), .B1(new_n780), .B2(new_n998), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G317), .A2(new_n778), .B1(new_n763), .B2(G303), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n785), .B2(new_n803), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n792), .B2(G311), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1039), .B1(new_n1042), .B2(KEYINPUT48), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(KEYINPUT48), .B2(new_n1042), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n581), .B(new_n1038), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1037), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1029), .B1(new_n1048), .B2(new_n757), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n697), .A2(new_n748), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT108), .Z(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n971), .B2(new_n984), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n739), .B1(new_n973), .B2(new_n974), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(KEYINPUT109), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n737), .A2(new_n971), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT110), .Z(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1054), .A2(KEYINPUT109), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1053), .B1(new_n1058), .B2(new_n1059), .ZN(G393));
  NAND2_X1  g0860(.A1(new_n982), .A2(new_n704), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n975), .A2(new_n981), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n984), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n981), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n965), .A2(new_n748), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n785), .A2(new_n999), .B1(new_n798), .B2(new_n777), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT52), .Z(new_n1068));
  OAI22_X1  g0868(.A1(new_n762), .A2(new_n1004), .B1(new_n772), .B2(new_n803), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n472), .B1(new_n780), .B2(new_n439), .C1(new_n376), .C2(new_n765), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G283), .C2(new_n831), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n827), .B2(new_n802), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n568), .B1(new_n254), .B2(new_n780), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n765), .A2(new_n523), .B1(new_n772), .B2(new_n1011), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n769), .A2(new_n326), .B1(new_n762), .B2(new_n281), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n827), .B2(new_n202), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n785), .A2(new_n828), .B1(new_n773), .B2(new_n777), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT51), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n1068), .A2(new_n1072), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n757), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n758), .B1(new_n442), .B2(new_n210), .C1(new_n755), .C2(new_n243), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1066), .A2(new_n745), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1065), .A2(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1063), .A2(new_n1084), .ZN(G390));
  AOI21_X1  g0885(.A(new_n878), .B1(new_n909), .B2(new_n877), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n889), .B1(new_n1086), .B2(new_n890), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n891), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n851), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n816), .B1(new_n714), .B2(new_n819), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n901), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1087), .A2(new_n1088), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n851), .B1(new_n877), .B2(new_n883), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n687), .B1(new_n710), .B2(new_n712), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n903), .B1(new_n1094), .B2(new_n818), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT111), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n900), .B(KEYINPUT112), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1093), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n922), .A2(G330), .A3(new_n819), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(new_n901), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT113), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT113), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1101), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n1092), .C2(new_n1098), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n736), .A2(new_n820), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n900), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1092), .A2(new_n1098), .A3(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(KEYINPUT114), .A3(new_n984), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT114), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n1064), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1090), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1107), .A2(new_n900), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n1101), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1096), .A2(new_n1108), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n930), .A2(G330), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n649), .A3(new_n913), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1112), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1124), .B(new_n1109), .C1(new_n1102), .C2(new_n1105), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n704), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1087), .A2(new_n1088), .A3(new_n746), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n742), .B1(new_n281), .B2(new_n846), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT115), .Z(new_n1131));
  OAI221_X1 g0931(.A(new_n472), .B1(new_n780), .B2(new_n254), .C1(new_n523), .C2(new_n769), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G68), .A2(new_n766), .B1(new_n800), .B2(G294), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n442), .B2(new_n762), .C1(new_n439), .C2(new_n777), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(G283), .C2(new_n786), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n376), .B2(new_n827), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT116), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n831), .A2(G150), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G50), .A2(new_n766), .B1(new_n800), .B2(G125), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n762), .B2(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n246), .B1(new_n780), .B2(new_n773), .C1(new_n833), .C2(new_n777), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1140), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(G128), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n785), .C1(new_n827), .C2(new_n1007), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1138), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1137), .B2(new_n1136), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1129), .B(new_n1131), .C1(new_n810), .C2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1114), .A2(new_n1128), .A3(new_n1150), .ZN(G378));
  XOR2_X1   g0951(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1152));
  NOR2_X1   g0952(.A1(new_n287), .A2(new_n684), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n298), .A2(new_n303), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1154), .B1(new_n298), .B2(new_n303), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1152), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1157), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1152), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n927), .A2(new_n928), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n921), .A2(new_n924), .B1(new_n909), .B2(new_n877), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1162), .B(G330), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1162), .B1(new_n929), .B2(G330), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1089), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n911), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1166), .A2(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT119), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(KEYINPUT120), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(G330), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1162), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1178), .A2(new_n892), .A3(new_n911), .A4(new_n1165), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT120), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1172), .A2(new_n1175), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1172), .B1(new_n1181), .B2(new_n1175), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1123), .B(KEYINPUT121), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1127), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1170), .A2(new_n1179), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(KEYINPUT57), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n704), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1178), .A2(new_n1165), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT119), .B1(new_n1193), .B2(new_n912), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT120), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1172), .A2(new_n1175), .A3(new_n1181), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n984), .A3(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G128), .A2(new_n778), .B1(new_n763), .B2(G137), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n769), .B2(new_n1142), .C1(new_n827), .C2(new_n833), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n786), .A2(G125), .B1(G150), .B2(new_n794), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT117), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n800), .A2(G124), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n766), .C2(G159), .ZN(new_n1208));
  AND4_X1   g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1030), .B1(new_n835), .B2(new_n765), .C1(new_n326), .C2(new_n780), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G107), .A2(new_n778), .B1(new_n800), .B2(G283), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n386), .B2(new_n762), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n581), .A2(new_n258), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n439), .B2(new_n785), .C1(new_n827), .C2(new_n442), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1213), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n757), .B1(new_n1209), .B2(new_n1220), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT118), .Z(new_n1222));
  AOI21_X1  g1022(.A(new_n742), .B1(new_n202), .B2(new_n846), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n1162), .C2(new_n747), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1199), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1192), .A2(new_n1225), .ZN(G375));
  AND3_X1   g1026(.A1(new_n1123), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n968), .B(KEYINPUT122), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1125), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT123), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1097), .A2(new_n746), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n757), .A2(G68), .A3(new_n746), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n777), .A2(new_n998), .B1(new_n780), .B2(new_n386), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT124), .Z(new_n1237));
  OAI21_X1  g1037(.A(new_n472), .B1(new_n765), .B2(new_n254), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n769), .A2(new_n442), .B1(new_n762), .B2(new_n376), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(G303), .C2(new_n800), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1237), .B(new_n1240), .C1(new_n1004), .C2(new_n785), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n827), .A2(new_n439), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n827), .A2(new_n1142), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n786), .A2(G132), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n777), .A2(new_n1007), .B1(new_n772), .B2(new_n1146), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G159), .B2(new_n831), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n794), .A2(G50), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n835), .A2(new_n765), .B1(new_n762), .B2(new_n828), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(new_n581), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1244), .A2(new_n1246), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n1241), .A2(new_n1242), .B1(new_n1243), .B2(new_n1250), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n742), .B(new_n1235), .C1(new_n1251), .C2(new_n757), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1120), .A2(new_n984), .B1(new_n1234), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1232), .A2(new_n1233), .A3(new_n1253), .ZN(G381));
  INV_X1    g1054(.A(new_n1225), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1191), .A2(G378), .A3(new_n1255), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1018), .B(G390), .C1(new_n986), .C2(new_n988), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G381), .A2(G384), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(G407));
  INV_X1    g1060(.A(new_n1256), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G407), .B(G213), .C1(G343), .C2(new_n1261), .ZN(G409));
  OAI211_X1 g1062(.A(G378), .B(new_n1225), .C1(new_n1187), .C2(new_n1190), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1114), .A2(new_n1128), .A3(new_n1150), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1186), .A2(new_n1197), .A3(new_n1198), .A4(new_n1229), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1188), .A2(new_n984), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1224), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1263), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n685), .A2(G213), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1228), .A2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1124), .A2(new_n739), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1228), .A2(KEYINPUT125), .A3(new_n1272), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT125), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1227), .B2(KEYINPUT60), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1273), .B(new_n1274), .C1(new_n1275), .C2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1253), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n849), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(G384), .A3(new_n1253), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .A4(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT61), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1263), .A2(new_n1268), .B1(G213), .B2(new_n685), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1286));
  INV_X1    g1086(.A(G2897), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1271), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1288), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1280), .A2(new_n1281), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1283), .B(new_n1284), .C1(new_n1285), .C2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1270), .B1(new_n1285), .B2(new_n1282), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT126), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(G390), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n989), .B2(new_n1019), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n989), .A2(new_n1019), .A3(new_n1296), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(G393), .B(new_n814), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1257), .B2(new_n1297), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1291), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1290), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1285), .A2(new_n1282), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT62), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1309), .A2(new_n1311), .A3(new_n1312), .A4(new_n1283), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1295), .A2(new_n1304), .A3(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(KEYINPUT63), .B1(new_n1292), .B2(new_n1285), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1310), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1304), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1282), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1316), .A2(new_n1317), .A3(new_n1284), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1314), .A2(new_n1319), .ZN(G405));
  NAND2_X1  g1120(.A1(G375), .A2(G378), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(new_n1261), .A3(new_n1286), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1264), .B1(new_n1192), .B2(new_n1225), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1282), .B1(new_n1323), .B2(new_n1256), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT127), .B1(new_n1325), .B2(new_n1304), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1317), .A2(new_n1322), .A3(new_n1327), .A4(new_n1324), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1325), .A2(new_n1304), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1326), .A2(new_n1328), .A3(new_n1329), .ZN(G402));
endmodule


