

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U552 ( .A1(n527), .A2(n526), .ZN(G160) );
  NOR2_X1 U553 ( .A1(n698), .A2(n972), .ZN(n691) );
  NOR2_X1 U554 ( .A1(n748), .A2(n968), .ZN(n751) );
  XNOR2_X1 U555 ( .A(n773), .B(KEYINPUT97), .ZN(n808) );
  NOR2_X1 U556 ( .A1(G651), .A2(n656), .ZN(n650) );
  XOR2_X1 U557 ( .A(n688), .B(KEYINPUT26), .Z(n517) );
  NOR2_X1 U558 ( .A1(n977), .A2(n517), .ZN(n690) );
  NOR2_X1 U559 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U560 ( .A1(G1966), .A2(n767), .ZN(n727) );
  NAND2_X1 U561 ( .A1(n775), .A2(n692), .ZN(n735) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n644) );
  XOR2_X1 U564 ( .A(KEYINPUT1), .B(n537), .Z(n654) );
  XOR2_X2 U565 ( .A(KEYINPUT17), .B(n518), .Z(n855) );
  NAND2_X1 U566 ( .A1(G137), .A2(n855), .ZN(n519) );
  XNOR2_X1 U567 ( .A(n519), .B(KEYINPUT64), .ZN(n527) );
  INV_X1 U568 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n522), .ZN(n859) );
  NAND2_X1 U570 ( .A1(G125), .A2(n859), .ZN(n521) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n860) );
  NAND2_X1 U572 ( .A1(G113), .A2(n860), .ZN(n520) );
  AND2_X1 U573 ( .A1(n521), .A2(n520), .ZN(n525) );
  AND2_X1 U574 ( .A1(n522), .A2(G2104), .ZN(n856) );
  NAND2_X1 U575 ( .A1(G101), .A2(n856), .ZN(n523) );
  XOR2_X1 U576 ( .A(KEYINPUT23), .B(n523), .Z(n524) );
  AND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U578 ( .A1(G138), .A2(n855), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G102), .A2(n856), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n533) );
  NAND2_X1 U581 ( .A1(G126), .A2(n859), .ZN(n531) );
  NAND2_X1 U582 ( .A1(G114), .A2(n860), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U584 ( .A1(n533), .A2(n532), .ZN(G164) );
  NAND2_X1 U585 ( .A1(G85), .A2(n644), .ZN(n535) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n656) );
  INV_X1 U587 ( .A(G651), .ZN(n536) );
  NOR2_X1 U588 ( .A1(n656), .A2(n536), .ZN(n645) );
  NAND2_X1 U589 ( .A1(G72), .A2(n645), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n541) );
  NOR2_X1 U591 ( .A1(G543), .A2(n536), .ZN(n537) );
  NAND2_X1 U592 ( .A1(G60), .A2(n654), .ZN(n539) );
  NAND2_X1 U593 ( .A1(G47), .A2(n650), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U595 ( .A1(n541), .A2(n540), .ZN(G290) );
  XNOR2_X1 U596 ( .A(G2451), .B(G2443), .ZN(n551) );
  XOR2_X1 U597 ( .A(G2446), .B(G2454), .Z(n543) );
  XNOR2_X1 U598 ( .A(KEYINPUT100), .B(G2435), .ZN(n542) );
  XNOR2_X1 U599 ( .A(n543), .B(n542), .ZN(n547) );
  XOR2_X1 U600 ( .A(KEYINPUT99), .B(G2438), .Z(n545) );
  XNOR2_X1 U601 ( .A(G1341), .B(G1348), .ZN(n544) );
  XNOR2_X1 U602 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U603 ( .A(n547), .B(n546), .Z(n549) );
  XNOR2_X1 U604 ( .A(G2430), .B(G2427), .ZN(n548) );
  XNOR2_X1 U605 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n551), .B(n550), .ZN(n552) );
  AND2_X1 U607 ( .A1(n552), .A2(G14), .ZN(G401) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  NAND2_X1 U610 ( .A1(G65), .A2(n654), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G53), .A2(n650), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G91), .A2(n644), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G78), .A2(n645), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U616 ( .A1(n558), .A2(n557), .ZN(n707) );
  INV_X1 U617 ( .A(n707), .ZN(G299) );
  NAND2_X1 U618 ( .A1(n650), .A2(G52), .ZN(n559) );
  XNOR2_X1 U619 ( .A(KEYINPUT65), .B(n559), .ZN(n568) );
  XOR2_X1 U620 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n560) );
  XNOR2_X1 U621 ( .A(KEYINPUT9), .B(n560), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G90), .A2(n644), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G77), .A2(n645), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U625 ( .A(n564), .B(n563), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G64), .A2(n654), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U628 ( .A1(n568), .A2(n567), .ZN(G171) );
  NAND2_X1 U629 ( .A1(G63), .A2(n654), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G51), .A2(n650), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U632 ( .A(KEYINPUT6), .B(n571), .ZN(n577) );
  NAND2_X1 U633 ( .A1(n644), .A2(G89), .ZN(n572) );
  XNOR2_X1 U634 ( .A(n572), .B(KEYINPUT4), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G76), .A2(n645), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U637 ( .A(n575), .B(KEYINPUT5), .Z(n576) );
  NOR2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT71), .B(n578), .Z(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT7), .B(n579), .Z(G168) );
  XOR2_X1 U641 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U642 ( .A1(G94), .A2(G452), .ZN(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT68), .B(n580), .Z(G173) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U646 ( .A(G223), .ZN(n826) );
  NAND2_X1 U647 ( .A1(n826), .A2(G567), .ZN(n582) );
  XOR2_X1 U648 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  NAND2_X1 U649 ( .A1(G56), .A2(n654), .ZN(n583) );
  XNOR2_X1 U650 ( .A(KEYINPUT14), .B(n583), .ZN(n584) );
  INV_X1 U651 ( .A(n584), .ZN(n590) );
  NAND2_X1 U652 ( .A1(n644), .A2(G81), .ZN(n585) );
  XNOR2_X1 U653 ( .A(n585), .B(KEYINPUT12), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G68), .A2(n645), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U656 ( .A(KEYINPUT13), .B(n588), .Z(n589) );
  NOR2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n650), .A2(G43), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n592), .A2(n591), .ZN(n977) );
  INV_X1 U660 ( .A(n977), .ZN(n593) );
  NAND2_X1 U661 ( .A1(n593), .A2(G860), .ZN(n594) );
  XNOR2_X1 U662 ( .A(KEYINPUT70), .B(n594), .ZN(G153) );
  INV_X1 U663 ( .A(G171), .ZN(G301) );
  NAND2_X1 U664 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U665 ( .A1(G79), .A2(n645), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G54), .A2(n650), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U668 ( .A1(G66), .A2(n654), .ZN(n598) );
  NAND2_X1 U669 ( .A1(G92), .A2(n644), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n601), .B(KEYINPUT15), .ZN(n972) );
  INV_X1 U673 ( .A(G868), .ZN(n669) );
  NAND2_X1 U674 ( .A1(n972), .A2(n669), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(G284) );
  NOR2_X1 U676 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U677 ( .A1(G286), .A2(n669), .ZN(n604) );
  NOR2_X1 U678 ( .A1(n605), .A2(n604), .ZN(G297) );
  INV_X1 U679 ( .A(G559), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G860), .A2(n606), .ZN(n607) );
  XNOR2_X1 U681 ( .A(n607), .B(KEYINPUT72), .ZN(n608) );
  NOR2_X1 U682 ( .A1(n972), .A2(n608), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT16), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT73), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n977), .ZN(n613) );
  INV_X1 U686 ( .A(n972), .ZN(n623) );
  NAND2_X1 U687 ( .A1(G868), .A2(n623), .ZN(n611) );
  NOR2_X1 U688 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U690 ( .A1(G123), .A2(n859), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n614), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n856), .A2(G99), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G135), .A2(n855), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G111), .A2(n860), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n914) );
  XNOR2_X1 U698 ( .A(G2096), .B(n914), .ZN(n622) );
  INV_X1 U699 ( .A(G2100), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U701 ( .A1(n623), .A2(G559), .ZN(n667) );
  XNOR2_X1 U702 ( .A(n977), .B(n667), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n624), .A2(G860), .ZN(n631) );
  NAND2_X1 U704 ( .A1(G67), .A2(n654), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G93), .A2(n644), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G80), .A2(n645), .ZN(n628) );
  NAND2_X1 U708 ( .A1(G55), .A2(n650), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  OR2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n670) );
  XOR2_X1 U711 ( .A(n631), .B(n670), .Z(G145) );
  NAND2_X1 U712 ( .A1(G73), .A2(n645), .ZN(n632) );
  XNOR2_X1 U713 ( .A(n632), .B(KEYINPUT2), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G61), .A2(n654), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G86), .A2(n644), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G48), .A2(n650), .ZN(n635) );
  XNOR2_X1 U718 ( .A(KEYINPUT75), .B(n635), .ZN(n636) );
  NOR2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U721 ( .A(KEYINPUT76), .B(n640), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G62), .A2(n654), .ZN(n642) );
  NAND2_X1 U723 ( .A1(G50), .A2(n650), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U725 ( .A(KEYINPUT77), .B(n643), .ZN(n649) );
  NAND2_X1 U726 ( .A1(G88), .A2(n644), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G75), .A2(n645), .ZN(n646) );
  AND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(G303) );
  INV_X1 U730 ( .A(G303), .ZN(G166) );
  NAND2_X1 U731 ( .A1(G49), .A2(n650), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U734 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n655), .B(KEYINPUT74), .ZN(n658) );
  NAND2_X1 U736 ( .A1(G87), .A2(n656), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(G288) );
  XOR2_X1 U738 ( .A(KEYINPUT19), .B(KEYINPUT78), .Z(n660) );
  XNOR2_X1 U739 ( .A(n707), .B(KEYINPUT79), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n660), .B(n659), .ZN(n663) );
  XNOR2_X1 U741 ( .A(G166), .B(G288), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n661), .B(n977), .ZN(n662) );
  XNOR2_X1 U743 ( .A(n663), .B(n662), .ZN(n665) );
  XOR2_X1 U744 ( .A(G290), .B(n670), .Z(n664) );
  XNOR2_X1 U745 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U746 ( .A(G305), .B(n666), .ZN(n895) );
  XNOR2_X1 U747 ( .A(n667), .B(n895), .ZN(n668) );
  NAND2_X1 U748 ( .A1(n668), .A2(G868), .ZN(n672) );
  NAND2_X1 U749 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U755 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U757 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NOR2_X1 U758 ( .A1(G219), .A2(G220), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U760 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U761 ( .A1(G96), .A2(n679), .ZN(n831) );
  AND2_X1 U762 ( .A1(G2106), .A2(n831), .ZN(n684) );
  NAND2_X1 U763 ( .A1(G108), .A2(G120), .ZN(n680) );
  NOR2_X1 U764 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U765 ( .A1(G69), .A2(n681), .ZN(n830) );
  NAND2_X1 U766 ( .A1(G567), .A2(n830), .ZN(n682) );
  XOR2_X1 U767 ( .A(KEYINPUT80), .B(n682), .Z(n683) );
  NOR2_X1 U768 ( .A1(n684), .A2(n683), .ZN(G319) );
  INV_X1 U769 ( .A(G319), .ZN(n902) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n685) );
  NOR2_X1 U771 ( .A1(n902), .A2(n685), .ZN(n829) );
  NAND2_X1 U772 ( .A1(n829), .A2(G36), .ZN(G176) );
  NOR2_X2 U773 ( .A1(G164), .A2(G1384), .ZN(n775) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n774) );
  INV_X1 U775 ( .A(n774), .ZN(n692) );
  NAND2_X1 U776 ( .A1(G8), .A2(n735), .ZN(n767) );
  AND2_X1 U777 ( .A1(G160), .A2(G40), .ZN(n687) );
  AND2_X1 U778 ( .A1(G1996), .A2(n775), .ZN(n686) );
  NAND2_X1 U779 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U780 ( .A1(G1341), .A2(n735), .ZN(n689) );
  NAND2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n698) );
  XNOR2_X1 U782 ( .A(n691), .B(KEYINPUT87), .ZN(n697) );
  AND2_X1 U783 ( .A1(n775), .A2(n692), .ZN(n712) );
  AND2_X1 U784 ( .A1(n712), .A2(G2067), .ZN(n693) );
  XOR2_X1 U785 ( .A(n693), .B(KEYINPUT88), .Z(n695) );
  NAND2_X1 U786 ( .A1(n735), .A2(G1348), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n698), .A2(n972), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n705) );
  NAND2_X1 U791 ( .A1(n712), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U792 ( .A(n701), .B(KEYINPUT27), .ZN(n703) );
  INV_X1 U793 ( .A(G1956), .ZN(n991) );
  NOR2_X1 U794 ( .A1(n991), .A2(n712), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U799 ( .A(n708), .B(KEYINPUT28), .Z(n709) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U801 ( .A(KEYINPUT29), .B(n711), .Z(n716) );
  INV_X1 U802 ( .A(G1961), .ZN(n1002) );
  NAND2_X1 U803 ( .A1(n735), .A2(n1002), .ZN(n714) );
  XNOR2_X1 U804 ( .A(KEYINPUT25), .B(G2078), .ZN(n945) );
  NAND2_X1 U805 ( .A1(n712), .A2(n945), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U807 ( .A1(G171), .A2(n717), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n725) );
  NOR2_X1 U809 ( .A1(G171), .A2(n717), .ZN(n722) );
  NOR2_X1 U810 ( .A1(G2084), .A2(n735), .ZN(n728) );
  NOR2_X1 U811 ( .A1(n727), .A2(n728), .ZN(n718) );
  NAND2_X1 U812 ( .A1(G8), .A2(n718), .ZN(n719) );
  XNOR2_X1 U813 ( .A(KEYINPUT30), .B(n719), .ZN(n720) );
  NOR2_X1 U814 ( .A1(G168), .A2(n720), .ZN(n721) );
  XOR2_X1 U815 ( .A(KEYINPUT31), .B(n723), .Z(n724) );
  NAND2_X1 U816 ( .A1(n725), .A2(n724), .ZN(n732) );
  XNOR2_X1 U817 ( .A(n732), .B(KEYINPUT89), .ZN(n726) );
  NOR2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U819 ( .A1(G8), .A2(n728), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n747) );
  AND2_X1 U821 ( .A1(G286), .A2(G8), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n742) );
  INV_X1 U823 ( .A(G8), .ZN(n740) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n767), .ZN(n733) );
  XNOR2_X1 U825 ( .A(n733), .B(KEYINPUT90), .ZN(n734) );
  NOR2_X1 U826 ( .A1(G166), .A2(n734), .ZN(n738) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n735), .ZN(n736) );
  XNOR2_X1 U828 ( .A(n736), .B(KEYINPUT91), .ZN(n737) );
  NAND2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n739) );
  OR2_X1 U830 ( .A1(n740), .A2(n739), .ZN(n741) );
  AND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n745) );
  XOR2_X1 U832 ( .A(KEYINPUT92), .B(KEYINPUT32), .Z(n743) );
  XNOR2_X1 U833 ( .A(KEYINPUT93), .B(n743), .ZN(n744) );
  XNOR2_X1 U834 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n765) );
  INV_X1 U836 ( .A(n765), .ZN(n748) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n968) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n749) );
  XOR2_X1 U839 ( .A(n749), .B(KEYINPUT94), .Z(n750) );
  NAND2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U841 ( .A1(G288), .A2(G1976), .ZN(n752) );
  XOR2_X1 U842 ( .A(KEYINPUT95), .B(n752), .Z(n970) );
  NAND2_X1 U843 ( .A1(n753), .A2(n970), .ZN(n754) );
  NOR2_X1 U844 ( .A1(n767), .A2(n754), .ZN(n755) );
  OR2_X2 U845 ( .A1(KEYINPUT33), .A2(n755), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n968), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U847 ( .A1(n756), .A2(n767), .ZN(n758) );
  XOR2_X1 U848 ( .A(G305), .B(G1981), .Z(n959) );
  INV_X1 U849 ( .A(n959), .ZN(n757) );
  NOR2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n772) );
  NOR2_X1 U852 ( .A1(G305), .A2(G1981), .ZN(n761) );
  XOR2_X1 U853 ( .A(n761), .B(KEYINPUT24), .Z(n762) );
  OR2_X1 U854 ( .A1(n767), .A2(n762), .ZN(n770) );
  NOR2_X1 U855 ( .A1(G2090), .A2(G303), .ZN(n763) );
  NAND2_X1 U856 ( .A1(G8), .A2(n763), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U859 ( .A(n768), .B(KEYINPUT96), .ZN(n769) );
  AND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n821) );
  XNOR2_X1 U863 ( .A(G2067), .B(KEYINPUT37), .ZN(n818) );
  NAND2_X1 U864 ( .A1(G140), .A2(n855), .ZN(n777) );
  NAND2_X1 U865 ( .A1(G104), .A2(n856), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U867 ( .A(KEYINPUT34), .B(n778), .ZN(n785) );
  XNOR2_X1 U868 ( .A(KEYINPUT35), .B(KEYINPUT82), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n860), .A2(G116), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n859), .A2(G128), .ZN(n779) );
  XOR2_X1 U871 ( .A(KEYINPUT81), .B(n779), .Z(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U873 ( .A(n783), .B(n782), .Z(n784) );
  NOR2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U875 ( .A(KEYINPUT36), .B(n786), .ZN(n872) );
  NOR2_X1 U876 ( .A1(n818), .A2(n872), .ZN(n919) );
  NAND2_X1 U877 ( .A1(n821), .A2(n919), .ZN(n816) );
  XOR2_X1 U878 ( .A(KEYINPUT84), .B(G1991), .Z(n936) );
  NAND2_X1 U879 ( .A1(G95), .A2(n856), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G107), .A2(n860), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U882 ( .A1(G131), .A2(n855), .ZN(n790) );
  NAND2_X1 U883 ( .A1(G119), .A2(n859), .ZN(n789) );
  NAND2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U886 ( .A(n793), .B(KEYINPUT83), .Z(n849) );
  NOR2_X1 U887 ( .A1(n936), .A2(n849), .ZN(n804) );
  NAND2_X1 U888 ( .A1(n855), .A2(G141), .ZN(n794) );
  XNOR2_X1 U889 ( .A(KEYINPUT86), .B(n794), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G129), .A2(n859), .ZN(n796) );
  NAND2_X1 U891 ( .A1(G117), .A2(n860), .ZN(n795) );
  NAND2_X1 U892 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n856), .A2(G105), .ZN(n797) );
  XOR2_X1 U894 ( .A(KEYINPUT38), .B(n797), .Z(n798) );
  NOR2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U896 ( .A(KEYINPUT85), .B(n800), .Z(n801) );
  NAND2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n867) );
  AND2_X1 U898 ( .A1(n867), .A2(G1996), .ZN(n803) );
  NOR2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n921) );
  INV_X1 U900 ( .A(n821), .ZN(n805) );
  NOR2_X1 U901 ( .A1(n921), .A2(n805), .ZN(n813) );
  INV_X1 U902 ( .A(n813), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n816), .A2(n806), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n810) );
  XNOR2_X1 U905 ( .A(G1986), .B(G290), .ZN(n964) );
  NAND2_X1 U906 ( .A1(n964), .A2(n821), .ZN(n809) );
  NAND2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n824) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n867), .ZN(n924) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n811) );
  AND2_X1 U910 ( .A1(n936), .A2(n849), .ZN(n915) );
  NOR2_X1 U911 ( .A1(n811), .A2(n915), .ZN(n812) );
  NOR2_X1 U912 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U913 ( .A1(n924), .A2(n814), .ZN(n815) );
  XNOR2_X1 U914 ( .A(n815), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n818), .A2(n872), .ZN(n912) );
  NAND2_X1 U917 ( .A1(n819), .A2(n912), .ZN(n820) );
  XNOR2_X1 U918 ( .A(KEYINPUT98), .B(n820), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U924 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n829), .A2(n828), .ZN(G188) );
  XNOR2_X1 U927 ( .A(G120), .B(KEYINPUT101), .ZN(G236) );
  NOR2_X1 U928 ( .A1(n831), .A2(n830), .ZN(G325) );
  XOR2_X1 U929 ( .A(KEYINPUT102), .B(G325), .Z(G261) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NAND2_X1 U933 ( .A1(G100), .A2(n856), .ZN(n833) );
  NAND2_X1 U934 ( .A1(G112), .A2(n860), .ZN(n832) );
  NAND2_X1 U935 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n834), .B(KEYINPUT105), .ZN(n836) );
  NAND2_X1 U937 ( .A1(G136), .A2(n855), .ZN(n835) );
  NAND2_X1 U938 ( .A1(n836), .A2(n835), .ZN(n839) );
  NAND2_X1 U939 ( .A1(n859), .A2(G124), .ZN(n837) );
  XOR2_X1 U940 ( .A(KEYINPUT44), .B(n837), .Z(n838) );
  NOR2_X1 U941 ( .A1(n839), .A2(n838), .ZN(G162) );
  NAND2_X1 U942 ( .A1(G142), .A2(n855), .ZN(n841) );
  NAND2_X1 U943 ( .A1(G106), .A2(n856), .ZN(n840) );
  NAND2_X1 U944 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n842), .B(KEYINPUT45), .ZN(n847) );
  NAND2_X1 U946 ( .A1(G130), .A2(n859), .ZN(n844) );
  NAND2_X1 U947 ( .A1(G118), .A2(n860), .ZN(n843) );
  NAND2_X1 U948 ( .A1(n844), .A2(n843), .ZN(n845) );
  XOR2_X1 U949 ( .A(KEYINPUT106), .B(n845), .Z(n846) );
  NAND2_X1 U950 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n848), .B(G162), .ZN(n871) );
  XOR2_X1 U952 ( .A(KEYINPUT107), .B(KEYINPUT46), .Z(n851) );
  XNOR2_X1 U953 ( .A(n849), .B(KEYINPUT108), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U955 ( .A(n852), .B(KEYINPUT109), .Z(n854) );
  XNOR2_X1 U956 ( .A(G164), .B(KEYINPUT48), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n866) );
  NAND2_X1 U958 ( .A1(G139), .A2(n855), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G103), .A2(n856), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G127), .A2(n859), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G115), .A2(n860), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(KEYINPUT47), .B(n863), .Z(n864) );
  NOR2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n907) );
  XOR2_X1 U966 ( .A(n866), .B(n907), .Z(n869) );
  XOR2_X1 U967 ( .A(G160), .B(n867), .Z(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n874) );
  XNOR2_X1 U970 ( .A(n872), .B(n914), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(n875) );
  NOR2_X1 U972 ( .A1(G37), .A2(n875), .ZN(G395) );
  XNOR2_X1 U973 ( .A(G1991), .B(KEYINPUT41), .ZN(n885) );
  XOR2_X1 U974 ( .A(G1966), .B(G1961), .Z(n877) );
  XNOR2_X1 U975 ( .A(G1996), .B(G1981), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(n881) );
  XOR2_X1 U977 ( .A(G1956), .B(G1971), .Z(n879) );
  XNOR2_X1 U978 ( .A(G1986), .B(G1976), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U980 ( .A(n881), .B(n880), .Z(n883) );
  XNOR2_X1 U981 ( .A(KEYINPUT104), .B(G2474), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(G229) );
  XOR2_X1 U984 ( .A(KEYINPUT103), .B(G2084), .Z(n887) );
  XNOR2_X1 U985 ( .A(G2090), .B(G2072), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U987 ( .A(n888), .B(G2096), .Z(n890) );
  XNOR2_X1 U988 ( .A(G2067), .B(G2078), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n894) );
  XOR2_X1 U990 ( .A(KEYINPUT43), .B(G2678), .Z(n892) );
  XNOR2_X1 U991 ( .A(G2100), .B(KEYINPUT42), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U993 ( .A(n894), .B(n893), .Z(G227) );
  XNOR2_X1 U994 ( .A(G171), .B(n972), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n897), .B(G286), .ZN(n898) );
  NOR2_X1 U997 ( .A1(G37), .A2(n898), .ZN(n899) );
  XNOR2_X1 U998 ( .A(KEYINPUT110), .B(n899), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G229), .A2(G227), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(KEYINPUT49), .B(n900), .ZN(n901) );
  NOR2_X1 U1001 ( .A1(G395), .A2(n901), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(G401), .A2(n902), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(KEYINPUT111), .B(n903), .ZN(n904) );
  NOR2_X1 U1004 ( .A1(G397), .A2(n904), .ZN(n905) );
  NAND2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1008 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n1020) );
  INV_X1 U1009 ( .A(KEYINPUT55), .ZN(n955) );
  XOR2_X1 U1010 ( .A(G2072), .B(n907), .Z(n909) );
  XOR2_X1 U1011 ( .A(G164), .B(G2078), .Z(n908) );
  NOR2_X1 U1012 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(KEYINPUT114), .B(n910), .ZN(n911) );
  XNOR2_X1 U1014 ( .A(n911), .B(KEYINPUT50), .ZN(n913) );
  NAND2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n930) );
  XNOR2_X1 U1016 ( .A(G160), .B(G2084), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT112), .B(n922), .ZN(n927) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n925), .B(KEYINPUT51), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n928), .B(KEYINPUT113), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n931), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n955), .A2(n932), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(G29), .ZN(n1017) );
  XNOR2_X1 U1031 ( .A(KEYINPUT115), .B(G2090), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(n934), .B(G35), .ZN(n953) );
  XNOR2_X1 U1033 ( .A(G2084), .B(G34), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(n935), .B(KEYINPUT54), .ZN(n951) );
  XNOR2_X1 U1035 ( .A(n936), .B(G25), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(G2067), .B(G26), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(G1996), .B(G32), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(G28), .A2(n939), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(KEYINPUT116), .B(G2072), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(G33), .B(n940), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G27), .B(n945), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(KEYINPUT117), .B(n946), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(n949), .B(KEYINPUT53), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(n955), .B(n954), .ZN(n957) );
  INV_X1 U1051 ( .A(G29), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(G11), .A2(n958), .ZN(n1015) );
  XNOR2_X1 U1054 ( .A(KEYINPUT56), .B(G16), .ZN(n983) );
  XNOR2_X1 U1055 ( .A(G168), .B(G1966), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(n961), .B(KEYINPUT57), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(KEYINPUT118), .B(n962), .ZN(n981) );
  XNOR2_X1 U1059 ( .A(G166), .B(G1971), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G1956), .B(G299), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(n971), .B(KEYINPUT119), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(G301), .B(G1961), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n972), .B(G1348), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G1341), .B(n977), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n1013) );
  XOR2_X1 U1074 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n990) );
  XNOR2_X1 U1075 ( .A(G1986), .B(G24), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(G1971), .B(G22), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1078 ( .A(G1976), .B(KEYINPUT122), .Z(n986) );
  XNOR2_X1 U1079 ( .A(G23), .B(n986), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(n990), .B(n989), .ZN(n1008) );
  XOR2_X1 U1082 ( .A(G1966), .B(G21), .Z(n1001) );
  XNOR2_X1 U1083 ( .A(G20), .B(n991), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G1981), .B(G6), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(G1341), .B(G19), .ZN(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n998) );
  XOR2_X1 U1088 ( .A(KEYINPUT59), .B(G1348), .Z(n996) );
  XNOR2_X1 U1089 ( .A(G4), .B(n996), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n999), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(KEYINPUT120), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1094 ( .A(G5), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1006), .B(KEYINPUT121), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(KEYINPUT61), .B(n1009), .Z(n1010) );
  NOR2_X1 U1099 ( .A1(G16), .A2(n1010), .ZN(n1011) );
  XOR2_X1 U1100 ( .A(KEYINPUT124), .B(n1011), .Z(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(n1018), .B(KEYINPUT62), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(n1020), .B(n1019), .ZN(G311) );
  XNOR2_X1 U1106 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

