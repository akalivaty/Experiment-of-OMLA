

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n669), .A2(n951), .ZN(n608) );
  AND2_X1 U553 ( .A1(n620), .A2(n619), .ZN(n521) );
  INV_X1 U554 ( .A(n992), .ZN(n619) );
  AND2_X1 U555 ( .A1(n621), .A2(n521), .ZN(n622) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n647) );
  XNOR2_X1 U557 ( .A(n648), .B(n647), .ZN(n653) );
  NAND2_X1 U558 ( .A1(n602), .A2(n711), .ZN(n669) );
  NOR2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n711) );
  NOR2_X1 U561 ( .A1(G651), .A2(n579), .ZN(n799) );
  OR2_X1 U562 ( .A1(n748), .A2(n747), .ZN(n762) );
  INV_X1 U563 ( .A(KEYINPUT87), .ZN(n539) );
  XOR2_X1 U564 ( .A(KEYINPUT65), .B(n533), .Z(G160) );
  INV_X1 U565 ( .A(G2105), .ZN(n536) );
  AND2_X1 U566 ( .A1(G2104), .A2(G101), .ZN(n522) );
  NAND2_X1 U567 ( .A1(n536), .A2(n522), .ZN(n523) );
  XNOR2_X1 U568 ( .A(n523), .B(KEYINPUT66), .ZN(n525) );
  INV_X1 U569 ( .A(KEYINPUT23), .ZN(n524) );
  XNOR2_X1 U570 ( .A(n525), .B(n524), .ZN(n527) );
  NOR2_X1 U571 ( .A1(G2104), .A2(n536), .ZN(n872) );
  NAND2_X1 U572 ( .A1(G125), .A2(n872), .ZN(n526) );
  NAND2_X1 U573 ( .A1(n527), .A2(n526), .ZN(n532) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n873) );
  NAND2_X1 U575 ( .A1(G113), .A2(n873), .ZN(n530) );
  XOR2_X2 U576 ( .A(KEYINPUT17), .B(n528), .Z(n878) );
  NAND2_X1 U577 ( .A1(G137), .A2(n878), .ZN(n529) );
  NAND2_X1 U578 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U579 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U580 ( .A1(G126), .A2(n872), .ZN(n535) );
  NAND2_X1 U581 ( .A1(G114), .A2(n873), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n542) );
  NAND2_X1 U583 ( .A1(G138), .A2(n878), .ZN(n538) );
  AND2_X1 U584 ( .A1(n536), .A2(G2104), .ZN(n876) );
  NAND2_X1 U585 ( .A1(G102), .A2(n876), .ZN(n537) );
  NAND2_X1 U586 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U587 ( .A(n540), .B(n539), .ZN(n541) );
  NOR2_X1 U588 ( .A1(n542), .A2(n541), .ZN(G164) );
  INV_X1 U589 ( .A(G651), .ZN(n549) );
  NOR2_X1 U590 ( .A1(G543), .A2(n549), .ZN(n544) );
  XNOR2_X1 U591 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n543) );
  XNOR2_X1 U592 ( .A(n544), .B(n543), .ZN(n798) );
  NAND2_X1 U593 ( .A1(n798), .A2(G65), .ZN(n545) );
  XOR2_X1 U594 ( .A(KEYINPUT71), .B(n545), .Z(n547) );
  XOR2_X1 U595 ( .A(G543), .B(KEYINPUT0), .Z(n579) );
  NAND2_X1 U596 ( .A1(n799), .A2(G53), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U598 ( .A(KEYINPUT72), .B(n548), .Z(n553) );
  NOR2_X1 U599 ( .A1(n579), .A2(n549), .ZN(n794) );
  NAND2_X1 U600 ( .A1(n794), .A2(G78), .ZN(n551) );
  NOR2_X1 U601 ( .A1(G651), .A2(G543), .ZN(n795) );
  NAND2_X1 U602 ( .A1(G91), .A2(n795), .ZN(n550) );
  AND2_X1 U603 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U604 ( .A1(n553), .A2(n552), .ZN(G299) );
  NAND2_X1 U605 ( .A1(G64), .A2(n798), .ZN(n555) );
  NAND2_X1 U606 ( .A1(G52), .A2(n799), .ZN(n554) );
  NAND2_X1 U607 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U608 ( .A1(G77), .A2(n794), .ZN(n557) );
  NAND2_X1 U609 ( .A1(G90), .A2(n795), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U612 ( .A1(n560), .A2(n559), .ZN(G171) );
  NAND2_X1 U613 ( .A1(G89), .A2(n795), .ZN(n561) );
  XNOR2_X1 U614 ( .A(n561), .B(KEYINPUT76), .ZN(n562) );
  XNOR2_X1 U615 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U616 ( .A1(G76), .A2(n794), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U618 ( .A(n565), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U619 ( .A1(G63), .A2(n798), .ZN(n567) );
  NAND2_X1 U620 ( .A1(G51), .A2(n799), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U622 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U623 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U624 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U625 ( .A1(n794), .A2(G75), .ZN(n572) );
  XNOR2_X1 U626 ( .A(n572), .B(KEYINPUT84), .ZN(n574) );
  NAND2_X1 U627 ( .A1(G88), .A2(n795), .ZN(n573) );
  NAND2_X1 U628 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U629 ( .A1(G62), .A2(n798), .ZN(n576) );
  NAND2_X1 U630 ( .A1(G50), .A2(n799), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U632 ( .A1(n578), .A2(n577), .ZN(G166) );
  XOR2_X1 U633 ( .A(KEYINPUT88), .B(G166), .Z(G303) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G49), .A2(n799), .ZN(n581) );
  NAND2_X1 U636 ( .A1(G87), .A2(n579), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U638 ( .A1(n798), .A2(n582), .ZN(n584) );
  NAND2_X1 U639 ( .A1(G651), .A2(G74), .ZN(n583) );
  NAND2_X1 U640 ( .A1(n584), .A2(n583), .ZN(G288) );
  NAND2_X1 U641 ( .A1(n799), .A2(G48), .ZN(n591) );
  NAND2_X1 U642 ( .A1(G86), .A2(n795), .ZN(n586) );
  NAND2_X1 U643 ( .A1(G61), .A2(n798), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U645 ( .A1(n794), .A2(G73), .ZN(n587) );
  XOR2_X1 U646 ( .A(KEYINPUT2), .B(n587), .Z(n588) );
  NOR2_X1 U647 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U648 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U649 ( .A(KEYINPUT83), .B(n592), .Z(G305) );
  NAND2_X1 U650 ( .A1(n794), .A2(G72), .ZN(n593) );
  XNOR2_X1 U651 ( .A(n593), .B(KEYINPUT68), .ZN(n600) );
  NAND2_X1 U652 ( .A1(n799), .A2(G47), .ZN(n595) );
  NAND2_X1 U653 ( .A1(n798), .A2(G60), .ZN(n594) );
  NAND2_X1 U654 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U655 ( .A1(G85), .A2(n795), .ZN(n596) );
  XNOR2_X1 U656 ( .A(KEYINPUT67), .B(n596), .ZN(n597) );
  NOR2_X1 U657 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U658 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U659 ( .A(KEYINPUT70), .B(n601), .ZN(G290) );
  AND2_X1 U660 ( .A1(G160), .A2(G40), .ZN(n602) );
  NAND2_X1 U661 ( .A1(G8), .A2(n669), .ZN(n704) );
  NOR2_X1 U662 ( .A1(G1966), .A2(n704), .ZN(n663) );
  INV_X1 U663 ( .A(G299), .ZN(n984) );
  INV_X1 U664 ( .A(n669), .ZN(n649) );
  NAND2_X1 U665 ( .A1(n649), .A2(G2072), .ZN(n603) );
  XNOR2_X1 U666 ( .A(n603), .B(KEYINPUT27), .ZN(n605) );
  AND2_X1 U667 ( .A1(G1956), .A2(n669), .ZN(n604) );
  NOR2_X1 U668 ( .A1(n605), .A2(n604), .ZN(n635) );
  NOR2_X1 U669 ( .A1(n984), .A2(n635), .ZN(n606) );
  XOR2_X1 U670 ( .A(n606), .B(KEYINPUT28), .Z(n646) );
  INV_X1 U671 ( .A(G1996), .ZN(n951) );
  INV_X1 U672 ( .A(KEYINPUT26), .ZN(n607) );
  XNOR2_X1 U673 ( .A(n608), .B(n607), .ZN(n621) );
  NAND2_X1 U674 ( .A1(n669), .A2(G1341), .ZN(n620) );
  NAND2_X1 U675 ( .A1(n795), .A2(G81), .ZN(n609) );
  XNOR2_X1 U676 ( .A(n609), .B(KEYINPUT12), .ZN(n611) );
  NAND2_X1 U677 ( .A1(G68), .A2(n794), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n613) );
  XOR2_X1 U679 ( .A(KEYINPUT13), .B(KEYINPUT74), .Z(n612) );
  XNOR2_X1 U680 ( .A(n613), .B(n612), .ZN(n616) );
  NAND2_X1 U681 ( .A1(n798), .A2(G56), .ZN(n614) );
  XOR2_X1 U682 ( .A(KEYINPUT14), .B(n614), .Z(n615) );
  NOR2_X1 U683 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U684 ( .A1(n799), .A2(G43), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n992) );
  XOR2_X1 U686 ( .A(KEYINPUT64), .B(n622), .Z(n640) );
  NAND2_X1 U687 ( .A1(G79), .A2(n794), .ZN(n624) );
  NAND2_X1 U688 ( .A1(G92), .A2(n795), .ZN(n623) );
  NAND2_X1 U689 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U690 ( .A1(G66), .A2(n798), .ZN(n626) );
  NAND2_X1 U691 ( .A1(G54), .A2(n799), .ZN(n625) );
  NAND2_X1 U692 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U693 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U694 ( .A(KEYINPUT15), .B(n629), .Z(n630) );
  XNOR2_X1 U695 ( .A(KEYINPUT75), .B(n630), .ZN(n977) );
  NOR2_X1 U696 ( .A1(n640), .A2(n977), .ZN(n631) );
  XOR2_X1 U697 ( .A(n631), .B(KEYINPUT98), .Z(n638) );
  AND2_X1 U698 ( .A1(n649), .A2(G2067), .ZN(n632) );
  XNOR2_X1 U699 ( .A(n632), .B(KEYINPUT99), .ZN(n634) );
  NAND2_X1 U700 ( .A1(n669), .A2(G1348), .ZN(n633) );
  NAND2_X1 U701 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U702 ( .A1(n984), .A2(n635), .ZN(n639) );
  AND2_X1 U703 ( .A1(n636), .A2(n639), .ZN(n637) );
  NAND2_X1 U704 ( .A1(n638), .A2(n637), .ZN(n644) );
  INV_X1 U705 ( .A(n639), .ZN(n642) );
  NAND2_X1 U706 ( .A1(n640), .A2(n977), .ZN(n641) );
  OR2_X1 U707 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U708 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U709 ( .A1(n646), .A2(n645), .ZN(n648) );
  OR2_X1 U710 ( .A1(n649), .A2(G1961), .ZN(n651) );
  XNOR2_X1 U711 ( .A(KEYINPUT25), .B(G2078), .ZN(n956) );
  NAND2_X1 U712 ( .A1(n649), .A2(n956), .ZN(n650) );
  NAND2_X1 U713 ( .A1(n651), .A2(n650), .ZN(n658) );
  NAND2_X1 U714 ( .A1(n658), .A2(G171), .ZN(n652) );
  NAND2_X1 U715 ( .A1(n653), .A2(n652), .ZN(n677) );
  NOR2_X1 U716 ( .A1(n669), .A2(G2084), .ZN(n654) );
  XNOR2_X1 U717 ( .A(n654), .B(KEYINPUT97), .ZN(n664) );
  NAND2_X1 U718 ( .A1(G8), .A2(n664), .ZN(n655) );
  NOR2_X1 U719 ( .A1(n663), .A2(n655), .ZN(n656) );
  XOR2_X1 U720 ( .A(KEYINPUT30), .B(n656), .Z(n657) );
  NOR2_X1 U721 ( .A1(G168), .A2(n657), .ZN(n660) );
  NOR2_X1 U722 ( .A1(G171), .A2(n658), .ZN(n659) );
  NOR2_X1 U723 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U724 ( .A(KEYINPUT31), .B(n661), .Z(n675) );
  AND2_X1 U725 ( .A1(n677), .A2(n675), .ZN(n662) );
  NOR2_X1 U726 ( .A1(n663), .A2(n662), .ZN(n667) );
  INV_X1 U727 ( .A(n664), .ZN(n665) );
  NAND2_X1 U728 ( .A1(G8), .A2(n665), .ZN(n666) );
  NAND2_X1 U729 ( .A1(n667), .A2(n666), .ZN(n685) );
  INV_X1 U730 ( .A(G8), .ZN(n674) );
  NOR2_X1 U731 ( .A1(G1971), .A2(n704), .ZN(n668) );
  XNOR2_X1 U732 ( .A(n668), .B(KEYINPUT100), .ZN(n671) );
  NOR2_X1 U733 ( .A1(n669), .A2(G2090), .ZN(n670) );
  NOR2_X1 U734 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U735 ( .A1(n672), .A2(G303), .ZN(n673) );
  OR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n678) );
  AND2_X1 U737 ( .A1(n675), .A2(n678), .ZN(n676) );
  NAND2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n681) );
  INV_X1 U739 ( .A(n678), .ZN(n679) );
  OR2_X1 U740 ( .A1(n679), .A2(G286), .ZN(n680) );
  NAND2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n683) );
  XOR2_X1 U742 ( .A(KEYINPUT101), .B(KEYINPUT32), .Z(n682) );
  XNOR2_X1 U743 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U744 ( .A1(n685), .A2(n684), .ZN(n703) );
  NOR2_X1 U745 ( .A1(G288), .A2(G1976), .ZN(n686) );
  XNOR2_X1 U746 ( .A(n686), .B(KEYINPUT102), .ZN(n981) );
  NOR2_X1 U747 ( .A1(G303), .A2(G1971), .ZN(n687) );
  XOR2_X1 U748 ( .A(n687), .B(KEYINPUT103), .Z(n688) );
  NOR2_X1 U749 ( .A1(n981), .A2(n688), .ZN(n689) );
  NAND2_X1 U750 ( .A1(n703), .A2(n689), .ZN(n690) );
  NAND2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n982) );
  NAND2_X1 U752 ( .A1(n690), .A2(n982), .ZN(n691) );
  NOR2_X1 U753 ( .A1(n691), .A2(n704), .ZN(n692) );
  OR2_X1 U754 ( .A1(n692), .A2(KEYINPUT33), .ZN(n698) );
  XOR2_X1 U755 ( .A(G1981), .B(KEYINPUT104), .Z(n693) );
  XNOR2_X1 U756 ( .A(G305), .B(n693), .ZN(n974) );
  INV_X1 U757 ( .A(n974), .ZN(n696) );
  NAND2_X1 U758 ( .A1(KEYINPUT33), .A2(n981), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n704), .A2(n694), .ZN(n695) );
  NOR2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n709) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n699) );
  XOR2_X1 U763 ( .A(n699), .B(KEYINPUT24), .Z(n700) );
  OR2_X1 U764 ( .A1(n704), .A2(n700), .ZN(n707) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n701) );
  NAND2_X1 U766 ( .A1(G8), .A2(n701), .ZN(n702) );
  NAND2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  AND2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n708) );
  AND2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n748) );
  XNOR2_X1 U771 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n710) );
  NOR2_X1 U773 ( .A1(n711), .A2(n710), .ZN(n759) );
  AND2_X1 U774 ( .A1(n978), .A2(n759), .ZN(n746) );
  XOR2_X1 U775 ( .A(KEYINPUT94), .B(G1991), .Z(n955) );
  NAND2_X1 U776 ( .A1(G107), .A2(n873), .ZN(n712) );
  XNOR2_X1 U777 ( .A(n712), .B(KEYINPUT92), .ZN(n715) );
  NAND2_X1 U778 ( .A1(G95), .A2(n876), .ZN(n713) );
  XOR2_X1 U779 ( .A(KEYINPUT93), .B(n713), .Z(n714) );
  NAND2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U781 ( .A1(G119), .A2(n872), .ZN(n717) );
  NAND2_X1 U782 ( .A1(G131), .A2(n878), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n889) );
  NOR2_X1 U785 ( .A1(n955), .A2(n889), .ZN(n730) );
  XOR2_X1 U786 ( .A(KEYINPUT38), .B(KEYINPUT96), .Z(n721) );
  NAND2_X1 U787 ( .A1(G105), .A2(n876), .ZN(n720) );
  XNOR2_X1 U788 ( .A(n721), .B(n720), .ZN(n726) );
  NAND2_X1 U789 ( .A1(G129), .A2(n872), .ZN(n723) );
  NAND2_X1 U790 ( .A1(G117), .A2(n873), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U792 ( .A(KEYINPUT95), .B(n724), .Z(n725) );
  NOR2_X1 U793 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U794 ( .A1(n878), .A2(G141), .ZN(n727) );
  NAND2_X1 U795 ( .A1(n728), .A2(n727), .ZN(n890) );
  AND2_X1 U796 ( .A1(n890), .A2(G1996), .ZN(n729) );
  NOR2_X1 U797 ( .A1(n730), .A2(n729), .ZN(n933) );
  INV_X1 U798 ( .A(n759), .ZN(n731) );
  NOR2_X1 U799 ( .A1(n933), .A2(n731), .ZN(n751) );
  INV_X1 U800 ( .A(n751), .ZN(n744) );
  NAND2_X1 U801 ( .A1(n873), .A2(G116), .ZN(n732) );
  XOR2_X1 U802 ( .A(KEYINPUT91), .B(n732), .Z(n734) );
  NAND2_X1 U803 ( .A1(n872), .A2(G128), .ZN(n733) );
  NAND2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U805 ( .A(KEYINPUT35), .B(n735), .Z(n742) );
  XNOR2_X1 U806 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n736) );
  XNOR2_X1 U807 ( .A(n736), .B(KEYINPUT34), .ZN(n740) );
  NAND2_X1 U808 ( .A1(G104), .A2(n876), .ZN(n738) );
  NAND2_X1 U809 ( .A1(G140), .A2(n878), .ZN(n737) );
  NAND2_X1 U810 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U811 ( .A(n740), .B(n739), .Z(n741) );
  NOR2_X1 U812 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U813 ( .A(KEYINPUT36), .B(n743), .ZN(n897) );
  XNOR2_X1 U814 ( .A(G2067), .B(KEYINPUT37), .ZN(n756) );
  NOR2_X1 U815 ( .A1(n897), .A2(n756), .ZN(n942) );
  NAND2_X1 U816 ( .A1(n759), .A2(n942), .ZN(n754) );
  NAND2_X1 U817 ( .A1(n744), .A2(n754), .ZN(n745) );
  OR2_X1 U818 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U819 ( .A1(G1996), .A2(n890), .ZN(n935) );
  NOR2_X1 U820 ( .A1(G1986), .A2(G290), .ZN(n749) );
  AND2_X1 U821 ( .A1(n955), .A2(n889), .ZN(n931) );
  NOR2_X1 U822 ( .A1(n749), .A2(n931), .ZN(n750) );
  NOR2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U824 ( .A1(n935), .A2(n752), .ZN(n753) );
  XNOR2_X1 U825 ( .A(n753), .B(KEYINPUT39), .ZN(n755) );
  NAND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n758) );
  AND2_X1 U827 ( .A1(n756), .A2(n897), .ZN(n757) );
  XNOR2_X1 U828 ( .A(n757), .B(KEYINPUT105), .ZN(n939) );
  NAND2_X1 U829 ( .A1(n758), .A2(n939), .ZN(n760) );
  NAND2_X1 U830 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U831 ( .A1(n762), .A2(n761), .ZN(n764) );
  XNOR2_X1 U832 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n763) );
  XNOR2_X1 U833 ( .A(n764), .B(n763), .ZN(G329) );
  AND2_X1 U834 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U835 ( .A(KEYINPUT79), .B(KEYINPUT18), .Z(n766) );
  NAND2_X1 U836 ( .A1(G123), .A2(n872), .ZN(n765) );
  XNOR2_X1 U837 ( .A(n766), .B(n765), .ZN(n773) );
  NAND2_X1 U838 ( .A1(G111), .A2(n873), .ZN(n768) );
  NAND2_X1 U839 ( .A1(G135), .A2(n878), .ZN(n767) );
  NAND2_X1 U840 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U841 ( .A1(n876), .A2(G99), .ZN(n769) );
  XOR2_X1 U842 ( .A(KEYINPUT80), .B(n769), .Z(n770) );
  NOR2_X1 U843 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U844 ( .A1(n773), .A2(n772), .ZN(n928) );
  XNOR2_X1 U845 ( .A(G2096), .B(n928), .ZN(n774) );
  OR2_X1 U846 ( .A1(G2100), .A2(n774), .ZN(G156) );
  INV_X1 U847 ( .A(G132), .ZN(G219) );
  INV_X1 U848 ( .A(G82), .ZN(G220) );
  NAND2_X1 U849 ( .A1(G7), .A2(G661), .ZN(n775) );
  XNOR2_X1 U850 ( .A(n775), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U851 ( .A(G223), .ZN(n824) );
  NAND2_X1 U852 ( .A1(n824), .A2(G567), .ZN(n776) );
  XOR2_X1 U853 ( .A(KEYINPUT11), .B(n776), .Z(G234) );
  INV_X1 U854 ( .A(G860), .ZN(n829) );
  OR2_X1 U855 ( .A1(n992), .A2(n829), .ZN(G153) );
  INV_X1 U856 ( .A(G171), .ZN(G301) );
  NAND2_X1 U857 ( .A1(G868), .A2(G301), .ZN(n778) );
  INV_X1 U858 ( .A(G868), .ZN(n809) );
  NAND2_X1 U859 ( .A1(n977), .A2(n809), .ZN(n777) );
  NAND2_X1 U860 ( .A1(n778), .A2(n777), .ZN(G284) );
  NOR2_X1 U861 ( .A1(G286), .A2(n809), .ZN(n780) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n779) );
  NOR2_X1 U863 ( .A1(n780), .A2(n779), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n829), .A2(G559), .ZN(n781) );
  INV_X1 U865 ( .A(n977), .ZN(n900) );
  NAND2_X1 U866 ( .A1(n781), .A2(n900), .ZN(n782) );
  XNOR2_X1 U867 ( .A(n782), .B(KEYINPUT77), .ZN(n783) );
  XOR2_X1 U868 ( .A(KEYINPUT16), .B(n783), .Z(G148) );
  NOR2_X1 U869 ( .A1(n977), .A2(n809), .ZN(n784) );
  XOR2_X1 U870 ( .A(KEYINPUT78), .B(n784), .Z(n785) );
  NOR2_X1 U871 ( .A1(G559), .A2(n785), .ZN(n787) );
  NOR2_X1 U872 ( .A1(G868), .A2(n992), .ZN(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(G282) );
  XNOR2_X1 U874 ( .A(KEYINPUT19), .B(KEYINPUT85), .ZN(n789) );
  XNOR2_X1 U875 ( .A(G288), .B(KEYINPUT86), .ZN(n788) );
  XNOR2_X1 U876 ( .A(n789), .B(n788), .ZN(n790) );
  XNOR2_X1 U877 ( .A(G305), .B(n790), .ZN(n792) );
  XNOR2_X1 U878 ( .A(G290), .B(G166), .ZN(n791) );
  XNOR2_X1 U879 ( .A(n792), .B(n791), .ZN(n793) );
  XNOR2_X1 U880 ( .A(n984), .B(n793), .ZN(n806) );
  NAND2_X1 U881 ( .A1(G80), .A2(n794), .ZN(n797) );
  NAND2_X1 U882 ( .A1(G93), .A2(n795), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n804) );
  NAND2_X1 U884 ( .A1(G67), .A2(n798), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G55), .A2(n799), .ZN(n800) );
  NAND2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U887 ( .A(KEYINPUT81), .B(n802), .Z(n803) );
  NOR2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U889 ( .A(KEYINPUT82), .B(n805), .Z(n830) );
  XOR2_X1 U890 ( .A(n806), .B(n830), .Z(n903) );
  NAND2_X1 U891 ( .A1(G559), .A2(n900), .ZN(n807) );
  XOR2_X1 U892 ( .A(n992), .B(n807), .Z(n828) );
  XNOR2_X1 U893 ( .A(n903), .B(n828), .ZN(n808) );
  NAND2_X1 U894 ( .A1(n808), .A2(G868), .ZN(n811) );
  NAND2_X1 U895 ( .A1(n809), .A2(n830), .ZN(n810) );
  NAND2_X1 U896 ( .A1(n811), .A2(n810), .ZN(G295) );
  NAND2_X1 U897 ( .A1(G2078), .A2(G2084), .ZN(n812) );
  XOR2_X1 U898 ( .A(KEYINPUT20), .B(n812), .Z(n813) );
  NAND2_X1 U899 ( .A1(G2090), .A2(n813), .ZN(n814) );
  XNOR2_X1 U900 ( .A(KEYINPUT21), .B(n814), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n815), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U902 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  XNOR2_X1 U903 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U904 ( .A1(G108), .A2(G120), .ZN(n816) );
  NOR2_X1 U905 ( .A1(G237), .A2(n816), .ZN(n817) );
  NAND2_X1 U906 ( .A1(G69), .A2(n817), .ZN(n832) );
  NAND2_X1 U907 ( .A1(n832), .A2(G567), .ZN(n822) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n818) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n818), .Z(n819) );
  NOR2_X1 U910 ( .A1(G218), .A2(n819), .ZN(n820) );
  NAND2_X1 U911 ( .A1(G96), .A2(n820), .ZN(n833) );
  NAND2_X1 U912 ( .A1(n833), .A2(G2106), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n834) );
  NAND2_X1 U914 ( .A1(G483), .A2(G661), .ZN(n823) );
  NOR2_X1 U915 ( .A1(n834), .A2(n823), .ZN(n827) );
  NAND2_X1 U916 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U919 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(G188) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n831) );
  XNOR2_X1 U924 ( .A(n831), .B(n830), .ZN(G145) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G108), .ZN(G238) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  INV_X1 U928 ( .A(G69), .ZN(G235) );
  NOR2_X1 U929 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  INV_X1 U931 ( .A(n834), .ZN(G319) );
  XOR2_X1 U932 ( .A(G2096), .B(KEYINPUT43), .Z(n836) );
  XNOR2_X1 U933 ( .A(G2090), .B(KEYINPUT110), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n837), .B(G2678), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2100), .Z(n841) );
  XNOR2_X1 U939 ( .A(G2078), .B(G2084), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U942 ( .A(G1956), .B(G1961), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1966), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U945 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U949 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n853) );
  XOR2_X1 U951 ( .A(G1981), .B(G2474), .Z(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U953 ( .A1(n872), .A2(G124), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U955 ( .A1(G136), .A2(n878), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U957 ( .A(KEYINPUT112), .B(n857), .ZN(n860) );
  NAND2_X1 U958 ( .A1(G100), .A2(n876), .ZN(n858) );
  XNOR2_X1 U959 ( .A(KEYINPUT113), .B(n858), .ZN(n859) );
  NOR2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n873), .A2(G112), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U963 ( .A(KEYINPUT114), .B(n863), .Z(G162) );
  NAND2_X1 U964 ( .A1(G103), .A2(n876), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G139), .A2(n878), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U967 ( .A1(n872), .A2(G127), .ZN(n866) );
  XOR2_X1 U968 ( .A(KEYINPUT117), .B(n866), .Z(n868) );
  NAND2_X1 U969 ( .A1(n873), .A2(G115), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n924) );
  NAND2_X1 U973 ( .A1(G130), .A2(n872), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G118), .A2(n873), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n883) );
  NAND2_X1 U976 ( .A1(n876), .A2(G106), .ZN(n877) );
  XOR2_X1 U977 ( .A(KEYINPUT115), .B(n877), .Z(n880) );
  NAND2_X1 U978 ( .A1(n878), .A2(G142), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U980 ( .A(KEYINPUT45), .B(n881), .Z(n882) );
  NOR2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U982 ( .A(n924), .B(n884), .Z(n885) );
  XNOR2_X1 U983 ( .A(G162), .B(n885), .ZN(n894) );
  XOR2_X1 U984 ( .A(KEYINPUT116), .B(KEYINPUT118), .Z(n887) );
  XNOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n928), .B(n888), .ZN(n892) );
  XOR2_X1 U988 ( .A(n890), .B(n889), .Z(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U990 ( .A(n894), .B(n893), .Z(n896) );
  XNOR2_X1 U991 ( .A(G164), .B(G160), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U994 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U995 ( .A(n992), .B(G286), .ZN(n902) );
  XNOR2_X1 U996 ( .A(G171), .B(n900), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U999 ( .A1(G37), .A2(n905), .ZN(G397) );
  XOR2_X1 U1000 ( .A(KEYINPUT109), .B(G2446), .Z(n907) );
  XNOR2_X1 U1001 ( .A(KEYINPUT107), .B(G2451), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1003 ( .A(n908), .B(G2430), .Z(n910) );
  XNOR2_X1 U1004 ( .A(G1348), .B(G1341), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1006 ( .A(G2438), .B(G2435), .Z(n912) );
  XNOR2_X1 U1007 ( .A(KEYINPUT108), .B(G2454), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1009 ( .A(n914), .B(n913), .Z(n916) );
  XNOR2_X1 U1010 ( .A(G2443), .B(G2427), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n917), .A2(G14), .ZN(n923) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n923), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(n923), .ZN(G401) );
  XOR2_X1 U1021 ( .A(G2072), .B(n924), .Z(n926) );
  XOR2_X1 U1022 ( .A(G164), .B(G2078), .Z(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1024 ( .A(KEYINPUT50), .B(n927), .Z(n945) );
  XNOR2_X1 U1025 ( .A(G160), .B(G2084), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n938) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(n936), .B(KEYINPUT51), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(KEYINPUT119), .B(n943), .ZN(n944) );
  NOR2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1037 ( .A(n946), .B(KEYINPUT52), .Z(n947) );
  XNOR2_X1 U1038 ( .A(KEYINPUT120), .B(n947), .ZN(n948) );
  NOR2_X1 U1039 ( .A1(KEYINPUT55), .A2(n948), .ZN(n949) );
  XNOR2_X1 U1040 ( .A(KEYINPUT121), .B(n949), .ZN(n950) );
  NAND2_X1 U1041 ( .A1(n950), .A2(G29), .ZN(n1028) );
  XOR2_X1 U1042 ( .A(G2090), .B(G35), .Z(n966) );
  XNOR2_X1 U1043 ( .A(G32), .B(n951), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(n952), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n960) );
  XOR2_X1 U1048 ( .A(n955), .B(G25), .Z(n958) );
  XOR2_X1 U1049 ( .A(n956), .B(G27), .Z(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1053 ( .A(KEYINPUT122), .B(n963), .Z(n964) );
  XNOR2_X1 U1054 ( .A(n964), .B(KEYINPUT53), .ZN(n965) );
  NAND2_X1 U1055 ( .A1(n966), .A2(n965), .ZN(n969) );
  XNOR2_X1 U1056 ( .A(G34), .B(G2084), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n967), .ZN(n968) );
  NOR2_X1 U1058 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1059 ( .A(n970), .B(KEYINPUT55), .ZN(n972) );
  XNOR2_X1 U1060 ( .A(G29), .B(KEYINPUT123), .ZN(n971) );
  NAND2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n973), .ZN(n1026) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n998) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G168), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(n976), .B(KEYINPUT57), .ZN(n996) );
  XNOR2_X1 U1067 ( .A(G1348), .B(n977), .ZN(n979) );
  NOR2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n990) );
  XNOR2_X1 U1069 ( .A(G1961), .B(G301), .ZN(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n983) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n988) );
  XOR2_X1 U1072 ( .A(G303), .B(G1971), .Z(n986) );
  XNOR2_X1 U1073 ( .A(n984), .B(G1956), .ZN(n985) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1076 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1077 ( .A(KEYINPUT124), .B(n991), .ZN(n994) );
  XNOR2_X1 U1078 ( .A(G1341), .B(n992), .ZN(n993) );
  NOR2_X1 U1079 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1080 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1081 ( .A1(n998), .A2(n997), .ZN(n1024) );
  INV_X1 U1082 ( .A(G16), .ZN(n1022) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G21), .ZN(n1000) );
  XNOR2_X1 U1084 ( .A(G5), .B(G1961), .ZN(n999) );
  NOR2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1012) );
  XOR2_X1 U1086 ( .A(KEYINPUT126), .B(G4), .Z(n1002) );
  XNOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT59), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n1002), .B(n1001), .ZN(n1005) );
  XOR2_X1 U1089 ( .A(KEYINPUT125), .B(G1341), .Z(n1003) );
  XNOR2_X1 U1090 ( .A(G19), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(G1956), .B(G20), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G6), .B(G1981), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1096 ( .A(KEYINPUT60), .B(n1010), .Z(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(G1986), .B(G24), .Z(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1109 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1029), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

