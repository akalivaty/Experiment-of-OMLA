//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT24), .B(G110), .Z(new_n191));
  XNOR2_X1  g005(.A(G119), .B(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G128), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n196), .B(new_n198), .C1(G119), .C2(new_n197), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G110), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT70), .ZN(new_n205));
  OR3_X1    g019(.A1(new_n201), .A2(KEYINPUT70), .A3(G125), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n202), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n208), .B1(new_n207), .B2(new_n210), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n193), .B(new_n200), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(new_n210), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n202), .A2(new_n204), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  OAI22_X1  g032(.A1(new_n199), .A2(G110), .B1(new_n192), .B2(new_n191), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G137), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n222), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n214), .A2(new_n220), .A3(new_n225), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(new_n188), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n190), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n227), .A2(new_n228), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n189), .A2(G902), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n208), .A2(G143), .ZN(new_n239));
  INV_X1    g053(.A(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G146), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G143), .B(G146), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G128), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G137), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT64), .A2(G134), .ZN(new_n250));
  NOR2_X1   g064(.A1(KEYINPUT64), .A2(G134), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .A3(G134), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(G137), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n252), .A2(G131), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n254), .A2(new_n255), .ZN(new_n259));
  INV_X1    g073(.A(new_n251), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(KEYINPUT11), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT64), .A2(G134), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n258), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n247), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT1), .B1(new_n240), .B2(G146), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n240), .A2(G146), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n208), .A2(G143), .ZN(new_n268));
  OAI211_X1 g082(.A(G128), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n239), .B(new_n241), .C1(KEYINPUT1), .C2(new_n197), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n258), .B1(G134), .B2(G137), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n250), .A2(new_n251), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n272), .B1(new_n274), .B2(G137), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n259), .A2(new_n263), .A3(new_n258), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT2), .B(G113), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT67), .A2(G116), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT67), .A2(G116), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n280), .A2(new_n281), .A3(new_n195), .ZN(new_n282));
  INV_X1    g096(.A(G116), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT66), .B1(new_n283), .B2(G119), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT66), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n195), .A3(G116), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n278), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(KEYINPUT2), .B(G113), .Z(new_n289));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n283), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(G119), .A3(new_n279), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n289), .A2(new_n292), .A3(new_n284), .A4(new_n286), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n265), .A2(new_n277), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n265), .A2(new_n277), .A3(KEYINPUT30), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n300));
  OAI21_X1  g114(.A(G131), .B1(new_n252), .B2(new_n256), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n276), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n300), .B1(new_n302), .B2(new_n247), .ZN(new_n303));
  AOI211_X1 g117(.A(KEYINPUT65), .B(new_n246), .C1(new_n301), .C2(new_n276), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n277), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT30), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n299), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n297), .B1(new_n307), .B2(new_n294), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT26), .B(G101), .ZN(new_n309));
  NOR2_X1   g123(.A1(G237), .A2(G953), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G210), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n309), .B(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT31), .B1(new_n308), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n277), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n265), .A2(KEYINPUT65), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n302), .A2(new_n300), .A3(new_n247), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n294), .B(new_n298), .C1(new_n319), .C2(KEYINPUT30), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n320), .A2(KEYINPUT31), .A3(new_n314), .A4(new_n296), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n296), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n277), .A2(new_n265), .A3(new_n295), .A4(KEYINPUT28), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n324), .B(new_n325), .C1(new_n319), .C2(new_n295), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI22_X1  g141(.A1(new_n315), .A2(new_n322), .B1(new_n314), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT32), .ZN(new_n329));
  NOR2_X1   g143(.A1(G472), .A2(G902), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n327), .A2(new_n314), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n320), .A2(new_n314), .A3(new_n296), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT31), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n332), .B1(new_n335), .B2(new_n321), .ZN(new_n336));
  INV_X1    g150(.A(new_n330), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT32), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n340));
  INV_X1    g154(.A(new_n314), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n326), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n314), .B1(new_n320), .B2(new_n296), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT69), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT69), .B1(new_n342), .B2(new_n344), .ZN(new_n348));
  INV_X1    g162(.A(new_n265), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n294), .B1(new_n349), .B2(new_n316), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n323), .B1(new_n350), .B2(new_n296), .ZN(new_n351));
  INV_X1    g165(.A(new_n324), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n341), .A2(new_n340), .ZN(new_n354));
  AOI21_X1  g168(.A(G902), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n347), .A2(new_n348), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G472), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n238), .B1(new_n339), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(G210), .B1(G237), .B2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n269), .A2(new_n203), .A3(new_n270), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n243), .B(G125), .C1(new_n244), .C2(new_n245), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n223), .A2(G224), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(new_n367), .B2(G107), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n369));
  INV_X1    g183(.A(G107), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(G104), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(G107), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G101), .ZN(new_n374));
  INV_X1    g188(.A(G101), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n368), .A2(new_n371), .A3(new_n375), .A4(new_n372), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(KEYINPUT4), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n373), .A2(new_n378), .A3(G101), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n294), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n292), .A2(KEYINPUT5), .A3(new_n284), .A4(new_n286), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n283), .A2(KEYINPUT5), .A3(G119), .ZN(new_n382));
  INV_X1    g196(.A(G113), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n367), .A2(G107), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n370), .A2(G104), .ZN(new_n387));
  OAI21_X1  g201(.A(G101), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n376), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n389), .A3(new_n293), .ZN(new_n390));
  XNOR2_X1  g204(.A(G110), .B(G122), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n380), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT73), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n380), .B2(new_n390), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n394), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n366), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n391), .B(KEYINPUT8), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT74), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n390), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n385), .A2(new_n293), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n376), .A2(new_n388), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n403), .A3(new_n406), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n402), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT75), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n364), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n361), .A2(new_n362), .A3(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n364), .A2(KEYINPUT7), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n361), .A2(new_n362), .A3(new_n412), .A4(new_n414), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n392), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n188), .B1(new_n410), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n360), .B1(new_n400), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n396), .B1(new_n394), .B2(new_n392), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n396), .A2(new_n394), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n365), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n389), .B1(new_n385), .B2(new_n293), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n425), .B1(new_n403), .B2(new_n390), .ZN(new_n426));
  INV_X1    g240(.A(new_n409), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n401), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n392), .A2(new_n418), .ZN(new_n429));
  AOI21_X1  g243(.A(G902), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n424), .A2(new_n430), .A3(new_n359), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n421), .A2(KEYINPUT76), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT76), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n424), .A2(new_n430), .A3(new_n433), .A4(new_n359), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n223), .A2(G952), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(G234), .B2(G237), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(G898), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT84), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n188), .B(new_n223), .C1(G234), .C2(G237), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n432), .A2(new_n434), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT9), .B(G234), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n446), .A2(new_n187), .A3(G953), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n291), .A2(G122), .A3(new_n279), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n283), .A2(G122), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n370), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT81), .B1(new_n197), .B2(G143), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n240), .A3(G128), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n240), .A2(G128), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n455), .A2(new_n273), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n273), .B1(new_n455), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n451), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT14), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n449), .A2(new_n461), .A3(new_n450), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n291), .A2(KEYINPUT14), .A3(G122), .A4(new_n279), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n462), .A2(G107), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT83), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n455), .A2(new_n457), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n274), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n455), .A2(new_n273), .A3(new_n457), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n462), .A2(G107), .A3(new_n463), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .A4(new_n451), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n449), .A2(new_n450), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G107), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n451), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n468), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n452), .A2(new_n454), .A3(KEYINPUT13), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT13), .B1(new_n452), .B2(new_n454), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n478), .A2(new_n479), .A3(new_n456), .ZN(new_n480));
  INV_X1    g294(.A(G134), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT82), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT13), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n455), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n452), .A2(new_n454), .A3(KEYINPUT13), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n457), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT82), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(G134), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n477), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n448), .B1(new_n473), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n458), .B1(new_n475), .B2(new_n451), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n456), .B1(new_n455), .B2(new_n483), .ZN(new_n492));
  AOI211_X1 g306(.A(KEYINPUT82), .B(new_n481), .C1(new_n492), .C2(new_n485), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n487), .B1(new_n486), .B2(G134), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(new_n465), .A3(new_n472), .A4(new_n447), .ZN(new_n496));
  AOI21_X1  g310(.A(G902), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G478), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(KEYINPUT15), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n497), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G237), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n223), .A3(G214), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n240), .A2(KEYINPUT77), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT77), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G143), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n310), .A2(G214), .B1(new_n504), .B2(G143), .ZN(new_n507));
  OAI21_X1  g321(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n502), .A2(new_n505), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT77), .B(G143), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n510), .B(new_n258), .C1(new_n502), .C2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n510), .B1(new_n511), .B2(new_n502), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(KEYINPUT17), .A3(G131), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n513), .A2(new_n216), .A3(new_n211), .A4(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G113), .B(G122), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(new_n367), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n205), .A2(new_n206), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n218), .B1(new_n519), .B2(new_n208), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(new_n258), .ZN(new_n522));
  OAI221_X1 g336(.A(new_n520), .B1(new_n514), .B2(new_n522), .C1(new_n508), .C2(new_n521), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n516), .A2(new_n518), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n518), .B1(new_n516), .B2(new_n523), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT79), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n516), .A2(new_n523), .ZN(new_n527));
  INV_X1    g341(.A(new_n518), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(KEYINPUT79), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n188), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT80), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT80), .ZN(new_n532));
  AOI21_X1  g346(.A(G902), .B1(new_n525), .B2(KEYINPUT79), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n528), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT79), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n532), .B(new_n533), .C1(new_n536), .C2(new_n524), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(G475), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(G475), .A2(G902), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n213), .B1(new_n508), .B2(new_n512), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT78), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n519), .A2(KEYINPUT19), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n217), .A2(KEYINPUT19), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n544), .B2(new_n208), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT19), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n205), .B2(new_n206), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n217), .A2(KEYINPUT19), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n541), .B(new_n208), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n540), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n518), .B1(new_n551), .B2(new_n523), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n539), .B1(new_n552), .B2(new_n524), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT20), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(new_n539), .C1(new_n552), .C2(new_n524), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n500), .A2(new_n538), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G221), .B1(new_n446), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n269), .A2(new_n376), .A3(new_n388), .A4(new_n270), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n270), .A2(new_n269), .B1(new_n376), .B2(new_n388), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n302), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT12), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n377), .A2(new_n247), .A3(new_n379), .ZN(new_n567));
  INV_X1    g381(.A(new_n302), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n271), .A2(new_n389), .A3(KEYINPUT10), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT10), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n223), .A2(G227), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT71), .ZN(new_n574));
  XNOR2_X1  g388(.A(G110), .B(G140), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n578), .B(new_n302), .C1(new_n563), .C2(new_n564), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n566), .A2(new_n572), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n302), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n577), .B1(new_n582), .B2(new_n572), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n583), .B2(KEYINPUT72), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n580), .A2(KEYINPUT72), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G469), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n188), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n188), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n566), .A2(new_n572), .A3(new_n579), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n576), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n582), .A2(new_n577), .A3(new_n572), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n589), .B1(new_n594), .B2(G469), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n561), .B1(new_n588), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n445), .A2(new_n559), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n358), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NAND2_X1  g414(.A1(new_n328), .A2(new_n330), .ZN(new_n601));
  OAI21_X1  g415(.A(G472), .B1(new_n336), .B2(G902), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n237), .A4(new_n596), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT85), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT87), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n496), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n490), .A2(new_n496), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n490), .B(new_n496), .C1(new_n606), .C2(new_n605), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(G478), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n498), .A2(new_n188), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n497), .B2(new_n498), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n538), .A2(new_n557), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n424), .A2(new_n430), .A3(KEYINPUT86), .A4(new_n359), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n617), .A2(new_n442), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT86), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n421), .A2(new_n619), .A3(new_n431), .ZN(new_n620));
  INV_X1    g434(.A(new_n441), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n604), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT34), .B(G104), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  XOR2_X1   g439(.A(new_n497), .B(new_n499), .Z(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n538), .A3(new_n557), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n604), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT88), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n226), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n221), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n235), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n233), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n601), .A2(new_n602), .A3(new_n636), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n597), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  AOI21_X1  g454(.A(new_n329), .B1(new_n328), .B2(new_n330), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n336), .A2(KEYINPUT32), .A3(new_n337), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n357), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AND4_X1   g457(.A1(new_n596), .A2(new_n620), .A3(new_n618), .A4(new_n636), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n440), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n436), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n627), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n643), .A2(new_n644), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  INV_X1    g466(.A(KEYINPUT91), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n648), .B(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n596), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT90), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n308), .A2(new_n341), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n350), .A2(new_n341), .A3(new_n296), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n188), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(new_n641), .B2(new_n642), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT89), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n432), .A2(new_n434), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT38), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n615), .A2(new_n626), .ZN(new_n668));
  NOR4_X1   g482(.A1(new_n667), .A2(new_n443), .A3(new_n636), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n653), .B1(new_n659), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n657), .A2(new_n658), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n672), .A2(KEYINPUT91), .A3(new_n665), .A4(new_n669), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  INV_X1    g489(.A(KEYINPUT92), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n614), .A2(new_n615), .A3(new_n676), .A4(new_n648), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n614), .A2(new_n615), .A3(new_n648), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT92), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n643), .A2(new_n644), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  NOR2_X1   g495(.A1(new_n616), .A2(new_n622), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n580), .A2(KEYINPUT72), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n562), .B(KEYINPUT10), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n568), .B1(new_n684), .B2(new_n567), .ZN(new_n685));
  INV_X1    g499(.A(new_n572), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n576), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT72), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n683), .B1(new_n689), .B2(new_n580), .ZN(new_n690));
  OAI21_X1  g504(.A(G469), .B1(new_n690), .B2(G902), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n560), .A3(new_n588), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n643), .A2(new_n237), .A3(new_n682), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NOR2_X1   g510(.A1(new_n627), .A2(new_n622), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n643), .A2(new_n237), .A3(new_n697), .A4(new_n693), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  AND3_X1   g513(.A1(new_n559), .A2(new_n621), .A3(new_n636), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n618), .A2(new_n620), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n643), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  INV_X1    g518(.A(KEYINPUT94), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n341), .B1(new_n351), .B2(new_n352), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(new_n315), .B2(new_n322), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n330), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n602), .A2(new_n708), .A3(new_n237), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT93), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n602), .A2(new_n708), .A3(KEYINPUT93), .A4(new_n237), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n615), .A2(new_n626), .A3(new_n618), .A4(new_n620), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n714), .A2(new_n441), .A3(new_n692), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n705), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n713), .A2(new_n715), .A3(new_n705), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  AND3_X1   g534(.A1(new_n679), .A2(new_n677), .A3(new_n702), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n602), .A2(new_n708), .A3(new_n636), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT95), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n602), .A2(new_n708), .A3(KEYINPUT95), .A4(new_n636), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  NAND2_X1  g542(.A1(new_n593), .A2(KEYINPUT96), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT96), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n591), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n587), .B1(new_n732), .B2(new_n188), .ZN(new_n733));
  INV_X1    g547(.A(new_n588), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n560), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n666), .A2(new_n442), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n677), .A3(new_n679), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n643), .A2(new_n237), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n738), .A2(new_n739), .A3(KEYINPUT42), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT97), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n331), .A2(new_n338), .B1(G472), .B2(new_n356), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(new_n238), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n679), .A2(new_n677), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n643), .A2(KEYINPUT97), .A3(new_n237), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n743), .A2(new_n745), .A3(new_n746), .A4(new_n737), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n740), .B1(KEYINPUT42), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  INV_X1    g563(.A(new_n736), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n735), .A2(new_n627), .A3(new_n649), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n358), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  OAI21_X1  g567(.A(G469), .B1(new_n594), .B2(KEYINPUT45), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n729), .A2(new_n731), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n754), .B1(new_n755), .B2(KEYINPUT45), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n589), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n588), .B1(new_n757), .B2(KEYINPUT46), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n560), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n654), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n614), .A2(new_n538), .A3(new_n557), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n601), .A2(new_n602), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n636), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n762), .A2(new_n769), .A3(new_n750), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT98), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n767), .B2(new_n768), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n767), .A2(new_n771), .A3(new_n768), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n253), .ZN(G39));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n760), .B(new_n776), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n744), .A2(new_n643), .A3(new_n237), .A4(new_n736), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  INV_X1    g594(.A(new_n691), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n734), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(KEYINPUT49), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n237), .A2(new_n442), .A3(new_n560), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n784), .A2(new_n763), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(KEYINPUT49), .B2(new_n783), .ZN(new_n787));
  INV_X1    g601(.A(new_n667), .ZN(new_n788));
  OR3_X1    g602(.A1(new_n787), .A2(new_n665), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n233), .A2(new_n635), .A3(new_n649), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n792), .B(new_n560), .C1(new_n733), .C2(new_n734), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n714), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n664), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n680), .A2(new_n651), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n679), .A2(new_n677), .A3(new_n702), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n724), .B2(new_n725), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT100), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n596), .A2(new_n620), .A3(new_n618), .A4(new_n636), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n339), .B2(new_n357), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n801), .A2(new_n650), .B1(new_n664), .B2(new_n794), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT100), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n727), .A3(new_n803), .A4(new_n680), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT52), .B1(new_n796), .B2(new_n798), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n615), .A2(new_n500), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n445), .A2(new_n810), .ZN(new_n811));
  OAI22_X1  g625(.A1(new_n597), .A2(new_n637), .B1(new_n603), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT99), .ZN(new_n814));
  OAI221_X1 g628(.A(new_n814), .B1(new_n603), .B2(new_n811), .C1(new_n597), .C2(new_n637), .ZN(new_n815));
  INV_X1    g629(.A(new_n603), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n432), .A2(new_n434), .A3(new_n444), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n616), .A2(new_n817), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n358), .A2(new_n598), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n813), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n559), .A2(new_n596), .A3(new_n636), .A4(new_n648), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n643), .A3(new_n750), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n724), .A2(new_n725), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n752), .B(new_n822), .C1(new_n823), .C2(new_n738), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n694), .A2(new_n698), .A3(new_n703), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n717), .B2(new_n718), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n827), .A3(new_n748), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n791), .B1(new_n809), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT101), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(KEYINPUT101), .B(new_n791), .C1(new_n809), .C2(new_n828), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n799), .A2(new_n804), .A3(KEYINPUT52), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n748), .A3(new_n827), .A4(new_n825), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(new_n799), .B2(new_n804), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(KEYINPUT102), .A3(KEYINPUT53), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT102), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n747), .A2(KEYINPUT42), .ZN(new_n840));
  INV_X1    g654(.A(new_n740), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n694), .A2(new_n698), .A3(new_n703), .ZN(new_n843));
  INV_X1    g657(.A(new_n718), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n844), .B2(new_n716), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n807), .A2(new_n846), .A3(new_n825), .A4(new_n834), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n839), .B1(new_n847), .B2(new_n791), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n838), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n790), .B1(new_n833), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n791), .B1(new_n835), .B2(new_n836), .ZN(new_n851));
  INV_X1    g665(.A(new_n808), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n805), .B2(new_n806), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT103), .B1(new_n842), .B2(new_n845), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT103), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n827), .A2(new_n748), .A3(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n820), .A2(new_n824), .A3(new_n791), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n853), .A2(new_n854), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n851), .A2(new_n790), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT104), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n851), .A2(new_n858), .A3(KEYINPUT104), .A4(new_n790), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n850), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n765), .A2(new_n436), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT105), .Z(new_n866));
  NOR3_X1   g680(.A1(new_n788), .A2(new_n442), .A3(new_n692), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n713), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT50), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT106), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n736), .A2(new_n692), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n871), .B1(new_n866), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n726), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n866), .A2(new_n713), .A3(new_n750), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n783), .A2(new_n560), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n777), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n872), .A2(new_n237), .A3(new_n436), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n665), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n614), .A2(new_n615), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n876), .A2(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n870), .A2(new_n875), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n866), .A2(new_n702), .A3(new_n713), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n615), .A3(new_n614), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n435), .B(KEYINPUT107), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n743), .A2(new_n746), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n873), .B2(new_n874), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT48), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT48), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n893), .B(new_n890), .C1(new_n873), .C2(new_n874), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n889), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n870), .A2(KEYINPUT51), .A3(new_n875), .A4(new_n882), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n885), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n864), .A2(new_n897), .A3(KEYINPUT108), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(G952), .B2(G953), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT108), .B1(new_n864), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n789), .B1(new_n899), .B2(new_n900), .ZN(G75));
  OR2_X1    g715(.A1(new_n223), .A2(G952), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT111), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n422), .A2(new_n423), .A3(new_n365), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n400), .ZN(new_n906));
  XOR2_X1   g720(.A(KEYINPUT109), .B(KEYINPUT55), .Z(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n188), .B1(new_n851), .B2(new_n858), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(G210), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(KEYINPUT110), .B(KEYINPUT56), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n904), .B(new_n912), .C1(new_n910), .C2(new_n914), .ZN(G51));
  XNOR2_X1  g729(.A(new_n589), .B(KEYINPUT57), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n851), .A2(new_n790), .A3(new_n858), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n790), .B1(new_n851), .B2(new_n858), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT112), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n586), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n909), .A2(new_n756), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n920), .B1(new_n919), .B2(new_n586), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n903), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT113), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(KEYINPUT113), .B(new_n903), .C1(new_n923), .C2(new_n924), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(G54));
  NAND3_X1  g743(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n552), .A2(new_n524), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n930), .A2(KEYINPUT114), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT114), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n904), .B1(new_n930), .B2(new_n931), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G60));
  NAND2_X1  g749(.A1(new_n609), .A2(new_n610), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n612), .B(KEYINPUT59), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n864), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n917), .B2(new_n918), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT115), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT115), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n943), .B(new_n940), .C1(new_n917), .C2(new_n918), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n904), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n939), .B1(KEYINPUT116), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n945), .A2(KEYINPUT116), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(G63));
  XNOR2_X1  g762(.A(KEYINPUT117), .B(KEYINPUT60), .ZN(new_n949));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n851), .B2(new_n858), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n903), .B1(new_n952), .B2(new_n234), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n633), .B2(new_n952), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT61), .ZN(G66));
  NOR2_X1   g769(.A1(new_n845), .A2(new_n820), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(G953), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n223), .B1(new_n438), .B2(G224), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT118), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n398), .B(new_n399), .C1(G898), .C2(new_n223), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(G69));
  XOR2_X1   g776(.A(new_n307), .B(new_n544), .Z(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT119), .Z(new_n964));
  OAI21_X1  g778(.A(new_n801), .B1(new_n745), .B2(new_n650), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n727), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(KEYINPUT120), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT120), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n965), .B2(new_n727), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n671), .A3(new_n673), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT122), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT121), .ZN(new_n974));
  OR3_X1    g788(.A1(new_n971), .A2(new_n974), .A3(KEYINPUT62), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n971), .B2(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n739), .A2(new_n736), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n616), .A2(new_n627), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT123), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n656), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n779), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(new_n774), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n973), .A2(new_n977), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n964), .B1(new_n984), .B2(G953), .ZN(new_n985));
  INV_X1    g799(.A(new_n963), .ZN(new_n986));
  INV_X1    g800(.A(new_n714), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n762), .A2(new_n987), .A3(new_n890), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n779), .A2(new_n752), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(new_n774), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n990), .A2(KEYINPUT125), .A3(new_n748), .A4(new_n970), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT125), .ZN(new_n992));
  AOI22_X1  g806(.A1(new_n777), .A2(new_n778), .B1(new_n978), .B2(new_n751), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n773), .A2(new_n772), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n993), .B(new_n988), .C1(new_n994), .C2(new_n770), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n970), .A2(new_n748), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(G953), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n645), .A2(G953), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT124), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n986), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n223), .B1(G227), .B2(G900), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n985), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n985), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  NAND3_X1  g820(.A1(new_n991), .A2(new_n997), .A3(new_n956), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  AND3_X1   g823(.A1(new_n1007), .A2(KEYINPUT127), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(KEYINPUT127), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n341), .B(new_n308), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n833), .A2(new_n849), .ZN(new_n1013));
  INV_X1    g827(.A(new_n333), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1009), .B1(new_n1014), .B2(new_n344), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1012), .B(new_n903), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n973), .A2(new_n956), .A3(new_n977), .A4(new_n983), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1017), .A2(KEYINPUT126), .A3(new_n1009), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n660), .ZN(new_n1019));
  AOI21_X1  g833(.A(KEYINPUT126), .B1(new_n1017), .B2(new_n1009), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1016), .A2(new_n1021), .ZN(G57));
endmodule


