//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT4), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT81), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT81), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G101), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n202), .A2(new_n203), .A3(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT82), .B1(new_n199), .B2(new_n208), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n201), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n213), .B(new_n214), .C1(new_n216), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n215), .B2(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(KEYINPUT64), .A3(G143), .ZN(new_n222));
  INV_X1    g036(.A(new_n213), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(G146), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n199), .A2(new_n227), .A3(G101), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT83), .B1(new_n212), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n203), .B1(new_n202), .B2(new_n209), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n199), .A2(KEYINPUT82), .A3(new_n208), .ZN(new_n232));
  OAI211_X1 g046(.A(KEYINPUT4), .B(new_n200), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT83), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n226), .A4(new_n228), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n196), .A2(G104), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n204), .B1(new_n237), .B2(new_n198), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n239), .B1(new_n231), .B2(new_n232), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT84), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n210), .B2(new_n211), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n217), .A2(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n224), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT67), .B(G128), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n246), .B1(G143), .B2(new_n217), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n251), .B(KEYINPUT68), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT1), .B1(new_n215), .B2(G146), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G128), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n256), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT68), .B1(new_n261), .B2(new_n251), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n249), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n241), .A2(new_n244), .A3(KEYINPUT10), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI22_X1  g080(.A1(new_n265), .A2(KEYINPUT11), .B1(new_n266), .B2(G137), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT65), .A4(G134), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT66), .A2(G131), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n265), .A2(KEYINPUT11), .B1(new_n266), .B2(G137), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n245), .B1(new_n259), .B2(new_n253), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n249), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n242), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT10), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n236), .A2(new_n264), .A3(new_n276), .A4(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT73), .B(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G227), .ZN(new_n284));
  XOR2_X1   g098(.A(G110), .B(G140), .Z(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT85), .B1(new_n263), .B2(new_n242), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n248), .B1(new_n293), .B2(new_n254), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n240), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n289), .A2(new_n279), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n276), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(KEYINPUT12), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT12), .B1(new_n296), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(KEYINPUT86), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT86), .ZN(new_n301));
  AOI211_X1 g115(.A(new_n301), .B(KEYINPUT12), .C1(new_n296), .C2(new_n297), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n288), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n236), .A2(new_n264), .A3(new_n281), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n297), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n282), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n286), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n192), .B1(new_n308), .B2(new_n190), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n282), .B1(new_n300), .B2(new_n302), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n286), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n288), .A2(new_n305), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(G469), .A3(new_n312), .ZN(new_n313));
  AOI211_X1 g127(.A(KEYINPUT87), .B(new_n189), .C1(new_n309), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT87), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n303), .A2(new_n307), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n190), .A3(new_n191), .ZN(new_n317));
  INV_X1    g131(.A(new_n192), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n315), .B1(new_n319), .B2(new_n188), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G116), .ZN(new_n323));
  INV_X1    g137(.A(G116), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G119), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT5), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n326), .B(G113), .C1(KEYINPUT5), .C2(new_n323), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n325), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT2), .B(G113), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n241), .A2(new_n244), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n329), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n233), .A2(new_n334), .A3(new_n228), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G122), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n332), .A2(new_n337), .A3(new_n335), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(KEYINPUT6), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n342), .A3(new_n338), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n219), .A2(new_n225), .ZN(new_n344));
  INV_X1    g158(.A(G125), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n294), .B2(G125), .ZN(new_n348));
  INV_X1    g162(.A(G224), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(G953), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n348), .B(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n341), .A2(new_n343), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n346), .B1(new_n263), .B2(new_n345), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT88), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT7), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI22_X1  g171(.A1(new_n354), .A2(new_n357), .B1(new_n356), .B2(new_n350), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n337), .B(KEYINPUT8), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n242), .A2(new_n331), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n242), .A2(new_n331), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n348), .A2(new_n355), .A3(KEYINPUT7), .A4(new_n351), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n358), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n364), .B2(new_n340), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n353), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G210), .B1(G237), .B2(G902), .ZN(new_n367));
  XOR2_X1   g181(.A(new_n367), .B(KEYINPUT89), .Z(new_n368));
  XOR2_X1   g182(.A(new_n368), .B(KEYINPUT90), .Z(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n368), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n353), .A2(new_n365), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G214), .B1(G237), .B2(G902), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G475), .ZN(new_n378));
  NAND2_X1  g192(.A1(KEYINPUT18), .A2(G131), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT72), .B(G237), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n283), .A2(new_n380), .A3(G214), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n215), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n283), .A2(new_n380), .A3(G143), .A4(G214), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n379), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n379), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n382), .A2(KEYINPUT91), .A3(new_n387), .A4(new_n383), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G140), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G125), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n345), .A2(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT78), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n397), .A3(new_n217), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  OAI22_X1  g215(.A1(new_n400), .A2(new_n401), .B1(new_n217), .B2(new_n396), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n389), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT16), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n390), .A3(G125), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n393), .B2(new_n404), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n217), .ZN(new_n407));
  OAI211_X1 g221(.A(G146), .B(new_n405), .C1(new_n393), .C2(new_n404), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G131), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n382), .B2(new_n383), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n411), .B2(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n384), .A2(G131), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n382), .A2(new_n410), .A3(new_n383), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n415), .B2(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n403), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n193), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n403), .A2(new_n416), .A3(new_n419), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n378), .B1(new_n423), .B2(new_n191), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n403), .A2(new_n416), .A3(new_n419), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT19), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n395), .A2(new_n397), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n393), .A2(KEYINPUT19), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n217), .A3(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n429), .A2(new_n408), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n389), .A2(new_n402), .B1(new_n415), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT92), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n419), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n415), .A2(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n403), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT92), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n425), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(G475), .A2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT20), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n403), .A2(new_n432), .A3(new_n434), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n420), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n431), .A2(new_n432), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n422), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n438), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n424), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(G234), .A2(G237), .ZN(new_n449));
  INV_X1    g263(.A(G953), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n449), .A2(G952), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n283), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n452), .A2(G902), .A3(new_n449), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(G898), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT93), .ZN(new_n456));
  INV_X1    g270(.A(G122), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(G116), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n324), .A2(KEYINPUT93), .A3(G122), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(G116), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G107), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n196), .A3(new_n461), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n257), .A2(G128), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n467), .A3(G143), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n259), .A2(G143), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n266), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT95), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n266), .B1(new_n474), .B2(new_n469), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n468), .A2(new_n470), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n474), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n471), .A2(new_n472), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n465), .A2(new_n473), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(G134), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n471), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n460), .A2(KEYINPUT14), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT14), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n458), .A2(new_n483), .A3(new_n459), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n482), .A2(new_n484), .A3(new_n461), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n481), .B(new_n464), .C1(new_n485), .C2(new_n196), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G217), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n187), .A2(new_n488), .A3(G953), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n489), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n479), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n490), .A2(KEYINPUT96), .A3(new_n191), .A4(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G478), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n494), .A2(KEYINPUT15), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n493), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n448), .A2(new_n455), .A3(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n377), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n321), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n252), .A2(G119), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(G119), .B2(new_n259), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT24), .B(G110), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT23), .B1(new_n259), .B2(G119), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(new_n322), .B2(G128), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT77), .B(G110), .Z(new_n507));
  INV_X1    g321(.A(KEYINPUT23), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n506), .B(new_n507), .C1(new_n501), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n510), .B(new_n408), .C1(new_n400), .C2(new_n401), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n506), .B1(new_n501), .B2(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G110), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n409), .B(new_n513), .C1(new_n502), .C2(new_n503), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT22), .B(G137), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n511), .A2(new_n514), .A3(new_n518), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(G217), .A2(G902), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n488), .B2(G234), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT75), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(G902), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n520), .A2(new_n191), .A3(new_n521), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n528), .A2(KEYINPUT25), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n525), .B(KEYINPUT76), .Z(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n528), .B2(KEYINPUT25), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n527), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT80), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n226), .B1(new_n274), .B2(new_n275), .ZN(new_n537));
  INV_X1    g351(.A(new_n334), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n269), .A2(G134), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n266), .A2(G137), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n410), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AND4_X1   g356(.A1(KEYINPUT65), .A2(new_n268), .A3(new_n269), .A4(G134), .ZN(new_n543));
  AOI22_X1  g357(.A1(KEYINPUT65), .A2(new_n268), .B1(new_n269), .B2(G134), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n273), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n542), .B1(new_n545), .B2(G131), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n537), .B(new_n538), .C1(new_n294), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT71), .ZN(new_n548));
  INV_X1    g362(.A(new_n546), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n263), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT71), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n550), .A2(new_n551), .A3(new_n538), .A4(new_n537), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n293), .A2(new_n254), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n546), .B1(new_n553), .B2(new_n249), .ZN(new_n554));
  INV_X1    g368(.A(new_n275), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n344), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n334), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n548), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT28), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n283), .A2(new_n380), .A3(G210), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT27), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT26), .B(G101), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT28), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n547), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n560), .A2(KEYINPUT29), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n191), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n548), .A2(new_n552), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT70), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT30), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n572), .A2(KEYINPUT69), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(KEYINPUT69), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n573), .B(new_n574), .C1(new_n554), .C2(new_n557), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n550), .A2(KEYINPUT69), .A3(new_n572), .A4(new_n537), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n571), .B1(new_n577), .B2(new_n334), .ZN(new_n578));
  AOI211_X1 g392(.A(KEYINPUT70), .B(new_n538), .C1(new_n575), .C2(new_n576), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n570), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n564), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n566), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n559), .B2(KEYINPUT28), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT29), .B1(new_n584), .B2(new_n564), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n568), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G472), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT74), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n560), .A2(new_n564), .A3(new_n566), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT29), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n581), .B2(new_n580), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n589), .B(G472), .C1(new_n593), .C2(new_n568), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n564), .B(new_n570), .C1(new_n578), .C2(new_n579), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n560), .A2(new_n566), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n581), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT31), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n577), .A2(new_n334), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT70), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n577), .A2(new_n571), .A3(new_n334), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n604), .A2(KEYINPUT31), .A3(new_n564), .A4(new_n570), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n600), .A2(new_n605), .A3(new_n587), .A4(new_n191), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT32), .ZN(new_n607));
  INV_X1    g421(.A(new_n596), .ZN(new_n608));
  AOI21_X1  g422(.A(G902), .B1(new_n608), .B2(KEYINPUT31), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT32), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n587), .A4(new_n600), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n536), .B1(new_n595), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n500), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n209), .ZN(G3));
  NAND2_X1  g430(.A1(new_n319), .A2(new_n188), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT87), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n189), .B1(new_n309), .B2(new_n313), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n315), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n191), .B1(new_n596), .B2(new_n599), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n606), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n536), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n618), .A2(new_n620), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n618), .A2(new_n620), .A3(KEYINPUT97), .A4(new_n625), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n490), .A2(new_n191), .A3(new_n492), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n494), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(KEYINPUT100), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(KEYINPUT100), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n489), .A2(KEYINPUT98), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n487), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n487), .B2(new_n635), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT99), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n490), .A2(new_n637), .A3(new_n492), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT99), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n494), .A2(G902), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n634), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n448), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n455), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n353), .A2(new_n365), .A3(new_n371), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n371), .B1(new_n353), .B2(new_n365), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n648), .B(new_n375), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n628), .A2(new_n629), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n447), .A2(new_n497), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n656), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n366), .A2(new_n368), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n376), .B1(new_n659), .B2(new_n372), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n496), .B(new_n424), .C1(new_n440), .C2(new_n446), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n660), .A2(new_n661), .A3(KEYINPUT101), .A4(new_n648), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n628), .A2(new_n629), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n519), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n515), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n526), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n529), .B2(new_n531), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n624), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n321), .A2(new_n499), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  AOI21_X1  g489(.A(new_n671), .B1(new_n595), .B2(new_n612), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n451), .B1(new_n453), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n657), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n321), .A2(new_n676), .A3(new_n660), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  XOR2_X1   g495(.A(new_n678), .B(KEYINPUT39), .Z(new_n682));
  NAND2_X1  g496(.A1(new_n321), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT40), .Z(new_n684));
  NOR2_X1   g498(.A1(new_n447), .A2(new_n496), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n375), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n580), .A2(new_n564), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n191), .B1(new_n559), .B2(new_n564), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n686), .B1(new_n612), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n373), .B(KEYINPUT38), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n671), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT102), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n684), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NOR2_X1   g510(.A1(new_n647), .A2(new_n678), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n321), .A2(new_n676), .A3(new_n660), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NAND3_X1  g513(.A1(new_n612), .A2(new_n594), .A3(new_n588), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n287), .B1(new_n305), .B2(new_n282), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n296), .A2(new_n297), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n301), .B1(new_n702), .B2(KEYINPUT12), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n299), .A2(KEYINPUT86), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(new_n298), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n701), .B1(new_n705), .B2(new_n288), .ZN(new_n706));
  OAI21_X1  g520(.A(G469), .B1(new_n706), .B2(G902), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n317), .ZN(new_n709));
  OAI211_X1 g523(.A(KEYINPUT103), .B(G469), .C1(new_n706), .C2(G902), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n189), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n536), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n700), .A2(new_n711), .A3(new_n712), .A4(new_n652), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n700), .A2(new_n663), .A3(new_n711), .A4(new_n712), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  AND2_X1   g531(.A1(new_n711), .A2(new_n660), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n498), .A3(new_n676), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  XOR2_X1   g534(.A(new_n532), .B(KEYINPUT104), .Z(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n624), .ZN(new_n722));
  INV_X1    g536(.A(new_n651), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n711), .A2(new_n722), .A3(new_n723), .A4(new_n685), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NAND4_X1  g539(.A1(new_n711), .A2(new_n672), .A3(new_n660), .A4(new_n697), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  AND2_X1   g541(.A1(new_n607), .A2(new_n611), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n588), .A2(new_n594), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n721), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n370), .A2(new_n375), .A3(new_n372), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n319), .A2(new_n188), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n619), .A2(KEYINPUT105), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND4_X1   g551(.A1(KEYINPUT42), .A2(new_n731), .A3(new_n697), .A4(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(KEYINPUT106), .A3(new_n613), .A4(new_n697), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n737), .A2(new_n613), .A3(new_n697), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n738), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n410), .ZN(G33));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n679), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n737), .A2(new_n748), .A3(new_n613), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n311), .A2(new_n312), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(G469), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n751), .B1(new_n756), .B2(new_n192), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n318), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n317), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n188), .ZN(new_n760));
  INV_X1    g574(.A(new_n682), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n760), .A2(KEYINPUT108), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT108), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n646), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n448), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT43), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n624), .A3(new_n670), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n732), .B1(new_n768), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n764), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  XNOR2_X1  g588(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n760), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n730), .A2(new_n536), .A3(new_n697), .A4(new_n732), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT110), .Z(new_n779));
  NAND3_X1  g593(.A1(new_n759), .A2(new_n188), .A3(new_n775), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT111), .Z(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT112), .B(G140), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G42));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n767), .A2(new_n451), .A3(new_n722), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n777), .A2(new_n780), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n188), .B1(new_n709), .B2(new_n710), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n732), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n692), .A2(new_n375), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n786), .A2(new_n711), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT50), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n711), .A2(new_n732), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT117), .Z(new_n796));
  NAND2_X1  g610(.A1(new_n767), .A2(new_n451), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n794), .B1(new_n672), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n612), .A2(new_n690), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n712), .A2(new_n451), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n796), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n447), .A3(new_n765), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n789), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n791), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n798), .A2(new_n731), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT48), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n786), .A2(new_n718), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(G952), .A3(new_n450), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n765), .A2(new_n447), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n802), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n805), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n672), .A2(new_n697), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n737), .A2(new_n813), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n448), .A2(new_n497), .A3(new_n671), .A4(new_n678), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n321), .A2(new_n700), .A3(new_n732), .A4(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n749), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n700), .A2(new_n498), .A3(new_n670), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n711), .A2(new_n660), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n716), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n713), .A2(new_n724), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n377), .A2(new_n648), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n810), .B1(new_n824), .B2(new_n657), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n661), .A2(KEYINPUT113), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n628), .A2(new_n629), .A3(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n321), .B(new_n499), .C1(new_n613), .C2(new_n672), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n817), .A2(new_n822), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n745), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n618), .A2(new_n620), .A3(new_n660), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n670), .B(new_n679), .C1(new_n728), .C2(new_n729), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n726), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n670), .B(new_n697), .C1(new_n728), .C2(new_n729), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n659), .A2(new_n372), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n670), .A2(new_n678), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT114), .B1(new_n619), .B2(new_n840), .ZN(new_n841));
  AND4_X1   g655(.A1(KEYINPUT114), .A2(new_n319), .A3(new_n188), .A4(new_n840), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n838), .B(new_n691), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n680), .A2(new_n698), .A3(new_n726), .A4(new_n843), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT115), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  INV_X1    g663(.A(new_n834), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(KEYINPUT52), .A3(new_n698), .A4(new_n843), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n831), .A2(new_n848), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n828), .A2(new_n829), .ZN(new_n858));
  AND4_X1   g672(.A1(KEYINPUT53), .A2(new_n749), .A3(new_n814), .A4(new_n816), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n820), .B2(new_n821), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n713), .A2(new_n724), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(KEYINPUT116), .A3(new_n716), .A4(new_n719), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n858), .A2(new_n859), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n745), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n849), .A2(new_n851), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n856), .A2(new_n857), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n831), .A2(new_n855), .A3(new_n866), .ZN(new_n869));
  INV_X1    g683(.A(new_n854), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n869), .B1(new_n870), .B2(new_n855), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n868), .B1(new_n871), .B2(new_n857), .ZN(new_n872));
  OAI22_X1  g686(.A1(new_n812), .A2(new_n872), .B1(G952), .B2(G953), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n709), .A2(new_n710), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT49), .Z(new_n875));
  NOR3_X1   g689(.A1(new_n721), .A2(new_n189), .A3(new_n376), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n766), .ZN(new_n877));
  OR4_X1    g691(.A1(new_n800), .A2(new_n875), .A3(new_n692), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n873), .A2(new_n878), .ZN(G75));
  NOR2_X1   g693(.A1(new_n283), .A2(G952), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n341), .A2(new_n343), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n352), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n856), .A2(new_n867), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(G902), .A3(new_n368), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(G902), .A3(new_n369), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n884), .A2(new_n890), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT56), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n880), .B(new_n888), .C1(new_n889), .C2(new_n893), .ZN(G51));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n755), .B(KEYINPUT121), .ZN(new_n896));
  AOI211_X1 g710(.A(new_n191), .B(new_n896), .C1(new_n856), .C2(new_n867), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n192), .B(KEYINPUT57), .ZN(new_n898));
  AOI221_X4 g712(.A(KEYINPUT54), .B1(new_n865), .B2(new_n866), .C1(new_n854), .C2(new_n855), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n857), .B1(new_n856), .B2(new_n867), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n897), .B1(new_n901), .B2(new_n316), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n895), .B1(new_n902), .B2(new_n880), .ZN(new_n903));
  INV_X1    g717(.A(new_n880), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n852), .B1(new_n849), .B2(new_n851), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT53), .B1(new_n907), .B2(new_n831), .ZN(new_n908));
  INV_X1    g722(.A(new_n867), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT54), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n868), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n706), .B1(new_n911), .B2(new_n898), .ZN(new_n912));
  OAI211_X1 g726(.A(KEYINPUT122), .B(new_n904), .C1(new_n912), .C2(new_n897), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n903), .A2(new_n913), .ZN(G54));
  NAND2_X1  g728(.A1(KEYINPUT58), .A2(G475), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n885), .A2(G902), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n437), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n885), .A2(G902), .A3(new_n444), .A4(new_n916), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n904), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G60));
  INV_X1    g736(.A(new_n643), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT59), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n911), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n872), .B2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n880), .ZN(G63));
  XOR2_X1   g742(.A(new_n523), .B(KEYINPUT60), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n885), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n522), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n885), .A2(new_n668), .A3(new_n929), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n904), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n935), .A2(KEYINPUT124), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(KEYINPUT124), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n880), .B1(new_n930), .B2(new_n931), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(KEYINPUT124), .A3(new_n935), .A4(new_n933), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(G66));
  OAI21_X1  g755(.A(G953), .B1(new_n454), .B2(new_n349), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n858), .A2(new_n822), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n452), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n881), .B1(G898), .B2(new_n283), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT125), .Z(new_n946));
  XNOR2_X1  g760(.A(new_n944), .B(new_n946), .ZN(G69));
  NAND3_X1  g761(.A1(new_n731), .A2(new_n660), .A3(new_n685), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n770), .B2(new_n771), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n764), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n749), .A3(new_n837), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n781), .B(KEYINPUT111), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n951), .A2(new_n745), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n283), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n427), .A2(new_n428), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n577), .B(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n954), .B(new_n957), .C1(G227), .C2(new_n283), .ZN(new_n958));
  OAI21_X1  g772(.A(G900), .B1(new_n957), .B2(G227), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n452), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n695), .A2(KEYINPUT62), .A3(new_n837), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT62), .B1(new_n695), .B2(new_n837), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n825), .A2(new_n826), .ZN(new_n964));
  INV_X1    g778(.A(new_n732), .ZN(new_n965));
  NOR4_X1   g779(.A1(new_n683), .A2(new_n964), .A3(new_n614), .A4(new_n965), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT126), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n782), .A2(new_n963), .A3(new_n773), .A4(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(new_n283), .A3(new_n956), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n958), .A2(new_n960), .A3(new_n969), .ZN(G72));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  INV_X1    g786(.A(new_n943), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n953), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n604), .A2(new_n581), .A3(new_n570), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT127), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n687), .A3(new_n972), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n871), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n972), .B1(new_n968), .B2(new_n973), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n880), .B1(new_n980), .B2(new_n688), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n977), .A2(new_n979), .A3(new_n981), .ZN(G57));
endmodule


