//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT15), .B1(new_n203), .B2(G43gat), .ZN(new_n204));
  INV_X1    g003(.A(G43gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G50gat), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n204), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(G50gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT89), .B(G43gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(G50gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT88), .B(KEYINPUT15), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n216), .A2(KEYINPUT90), .A3(new_n208), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT90), .B1(new_n216), .B2(new_n208), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n215), .ZN(new_n220));
  NOR3_X1   g019(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n221));
  OAI22_X1  g020(.A1(new_n220), .A2(new_n221), .B1(new_n207), .B2(new_n208), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n204), .A2(new_n206), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(KEYINPUT87), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT87), .ZN(new_n225));
  AND2_X1   g024(.A1(G29gat), .A2(G36gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT14), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n207), .A3(new_n208), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n226), .B1(new_n228), .B2(new_n215), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n203), .A2(G43gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n210), .A2(new_n230), .A3(KEYINPUT15), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n225), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n214), .A2(new_n219), .B1(new_n224), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G15gat), .B(G22gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT16), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G1gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G8gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT91), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n239), .B1(new_n234), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G22gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G15gat), .ZN(new_n243));
  INV_X1    g042(.A(G15gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G22gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n245), .A3(new_n240), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(G8gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n238), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(G8gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n240), .A3(new_n239), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n237), .A4(new_n236), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n202), .B1(new_n233), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n224), .A2(new_n232), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n205), .A2(KEYINPUT89), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT89), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G43gat), .ZN(new_n257));
  AOI21_X1  g056(.A(G50gat), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n210), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n213), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n209), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n219), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n262), .A3(KEYINPUT17), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT92), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n254), .A2(new_n262), .A3(KEYINPUT92), .A4(KEYINPUT17), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n248), .A2(new_n251), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT17), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n262), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n253), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n202), .B(KEYINPUT13), .Z(new_n273));
  INV_X1    g072(.A(KEYINPUT95), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(new_n268), .B2(new_n270), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n268), .A2(new_n270), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n233), .A2(KEYINPUT95), .A3(new_n252), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n272), .A2(KEYINPUT18), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT94), .ZN(new_n280));
  XOR2_X1   g079(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n281));
  OAI21_X1  g080(.A(new_n280), .B1(new_n272), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n252), .B1(new_n233), .B2(KEYINPUT17), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n284), .B1(new_n265), .B2(new_n266), .ZN(new_n285));
  OAI211_X1 g084(.A(KEYINPUT94), .B(new_n283), .C1(new_n285), .C2(new_n253), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n279), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n288));
  XNOR2_X1  g087(.A(G113gat), .B(G141gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G169gat), .B(G197gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT12), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT96), .B1(new_n272), .B2(new_n281), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT96), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n297), .B(new_n283), .C1(new_n285), .C2(new_n253), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n279), .A2(new_n296), .A3(new_n298), .A4(new_n293), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT28), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT27), .B(G183gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(KEYINPUT65), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT27), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT65), .B1(new_n305), .B2(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n302), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n303), .A2(KEYINPUT28), .A3(new_n307), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G169gat), .ZN(new_n312));
  INV_X1    g111(.A(G176gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n314), .A2(KEYINPUT26), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n315), .A2(KEYINPUT26), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n311), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n315), .B(KEYINPUT23), .Z(new_n322));
  OR2_X1    g121(.A1(new_n317), .A2(KEYINPUT24), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT64), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n324), .A2(new_n325), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n324), .A2(new_n325), .ZN(new_n328));
  INV_X1    g127(.A(G183gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n307), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(KEYINPUT24), .A3(new_n317), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n322), .A2(new_n327), .A3(new_n328), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n323), .A3(new_n326), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n315), .B(KEYINPUT23), .ZN(new_n334));
  OAI22_X1  g133(.A1(new_n333), .A2(new_n334), .B1(new_n324), .B2(new_n325), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G113gat), .ZN(new_n337));
  INV_X1    g136(.A(G120gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(G113gat), .B2(G120gat), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT66), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G127gat), .B(G134gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n343), .B(KEYINPUT66), .C1(new_n339), .C2(new_n341), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n321), .A2(new_n336), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT67), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n321), .A2(new_n336), .ZN(new_n351));
  INV_X1    g150(.A(new_n347), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n311), .A2(new_n320), .B1(new_n332), .B2(new_n335), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT67), .A3(new_n347), .ZN(new_n355));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n350), .A2(new_n353), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT69), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT34), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n357), .B2(new_n358), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT32), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n350), .A2(new_n355), .A3(new_n353), .ZN(new_n365));
  INV_X1    g164(.A(new_n356), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT33), .B1(new_n365), .B2(new_n366), .ZN(new_n368));
  XOR2_X1   g167(.A(G15gat), .B(G43gat), .Z(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT68), .ZN(new_n370));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n367), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  AOI221_X4 g173(.A(new_n364), .B1(KEYINPUT33), .B2(new_n372), .C1(new_n365), .C2(new_n366), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n363), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT70), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT70), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(new_n363), .C1(new_n374), .C2(new_n375), .ZN(new_n379));
  INV_X1    g178(.A(new_n362), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n360), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT32), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n385), .A3(new_n372), .ZN(new_n386));
  INV_X1    g185(.A(new_n375), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n381), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n377), .A2(KEYINPUT36), .A3(new_n379), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n376), .A2(new_n388), .ZN(new_n390));
  XOR2_X1   g189(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G211gat), .B(G218gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT22), .B1(new_n398), .B2(G218gat), .ZN(new_n399));
  XOR2_X1   g198(.A(G197gat), .B(G204gat), .Z(new_n400));
  OAI21_X1  g199(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  INV_X1    g201(.A(G218gat), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n396), .B2(new_n397), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n402), .B(new_n394), .C1(new_n404), .C2(KEYINPUT22), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G226gat), .ZN(new_n408));
  INV_X1    g207(.A(G233gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(new_n351), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n410), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n354), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n407), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n354), .B2(KEYINPUT29), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT73), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n351), .A2(new_n417), .A3(new_n410), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT73), .B1(new_n354), .B2(new_n413), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n416), .A2(new_n418), .A3(new_n419), .A4(new_n406), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT74), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G92gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT75), .B(G64gat), .ZN(new_n425));
  XOR2_X1   g224(.A(new_n424), .B(new_n425), .Z(new_n426));
  INV_X1    g225(.A(KEYINPUT74), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n415), .A2(new_n420), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n426), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n420), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT30), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n431), .A2(new_n432), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n437));
  INV_X1    g236(.A(G155gat), .ZN(new_n438));
  INV_X1    g237(.A(G162gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G155gat), .A2(G162gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT76), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(KEYINPUT76), .A3(new_n441), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(KEYINPUT2), .ZN(new_n446));
  INV_X1    g245(.A(G141gat), .ZN(new_n447));
  INV_X1    g246(.A(G148gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G141gat), .A2(G148gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n442), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n449), .A2(new_n450), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT76), .A4(new_n446), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(new_n347), .ZN(new_n457));
  NAND2_X1  g256(.A1(G225gat), .A2(G233gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n437), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n352), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n458), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n456), .A2(new_n347), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT4), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n456), .A2(new_n468), .A3(new_n347), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n460), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n464), .A2(new_n458), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT78), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n466), .A2(new_n473), .A3(KEYINPUT4), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n467), .A2(KEYINPUT78), .A3(new_n469), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n472), .A2(new_n437), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G1gat), .B(G29gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT0), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(G57gat), .ZN(new_n479));
  INV_X1    g278(.A(G85gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n471), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT79), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n471), .A2(new_n476), .ZN(new_n485));
  INV_X1    g284(.A(new_n481), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n471), .A2(new_n476), .A3(KEYINPUT79), .A4(new_n481), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n484), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n487), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT6), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n436), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G78gat), .B(G106gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n406), .A2(new_n411), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n456), .B1(new_n496), .B2(new_n461), .ZN(new_n497));
  NAND2_X1  g296(.A1(G228gat), .A2(G233gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT29), .B1(new_n456), .B2(new_n461), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(new_n406), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT81), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n500), .A2(new_n406), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT29), .B1(new_n401), .B2(new_n405), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n455), .B(new_n452), .C1(new_n504), .C2(KEYINPUT3), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n503), .A2(new_n505), .A3(new_n506), .A4(new_n499), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n500), .A2(new_n406), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT80), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n497), .A2(KEYINPUT80), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n499), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n508), .A2(new_n513), .A3(G22gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n512), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n498), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n502), .A2(new_n507), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n242), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n495), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT31), .B(G50gat), .ZN(new_n520));
  OAI21_X1  g319(.A(G22gat), .B1(new_n508), .B2(new_n513), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n242), .A3(new_n517), .ZN(new_n522));
  INV_X1    g321(.A(new_n495), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n520), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n523), .B1(new_n521), .B2(new_n522), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n494), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n393), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT82), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT82), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n393), .A2(new_n533), .A3(new_n530), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n416), .B1(new_n413), .B2(new_n354), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n406), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n416), .A2(new_n418), .A3(new_n419), .A4(new_n407), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT38), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n415), .A2(new_n420), .A3(new_n535), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n426), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT85), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT38), .B1(new_n537), .B2(new_n538), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT85), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n546), .A3(new_n426), .A4(new_n542), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n490), .A2(new_n492), .A3(new_n431), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n422), .A2(KEYINPUT37), .A3(new_n428), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT38), .B1(new_n551), .B2(new_n543), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n550), .A2(new_n552), .B1(new_n525), .B2(new_n529), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n475), .A2(new_n464), .A3(new_n474), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n459), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(KEYINPUT39), .C1(new_n459), .C2(new_n457), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT39), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n557), .A3(new_n459), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n558), .A2(KEYINPUT83), .A3(new_n481), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT83), .B1(new_n558), .B2(new_n481), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT40), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(KEYINPUT40), .B(new_n556), .C1(new_n559), .C2(new_n560), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n563), .A2(new_n435), .A3(new_n487), .A4(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT84), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n431), .B(KEYINPUT30), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n491), .B1(new_n568), .B2(new_n429), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n569), .A2(KEYINPUT84), .A3(new_n564), .A4(new_n563), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n532), .A2(new_n534), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n379), .A2(new_n388), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n386), .A2(new_n387), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n378), .B1(new_n575), .B2(new_n363), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n529), .A2(new_n525), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n490), .A2(new_n492), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(new_n435), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT35), .ZN(new_n583));
  INV_X1    g382(.A(new_n390), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n578), .A2(new_n580), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n301), .B1(new_n573), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(G211gat), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT21), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G71gat), .ZN(new_n596));
  INV_X1    g395(.A(G78gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G57gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G64gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(KEYINPUT98), .A2(G64gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(KEYINPUT98), .A2(G64gat), .ZN(new_n605));
  OAI21_X1  g404(.A(G57gat), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(KEYINPUT99), .B(G57gat), .C1(new_n604), .C2(new_n605), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n600), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n598), .A2(new_n599), .ZN(new_n611));
  INV_X1    g410(.A(G64gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(G57gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n594), .B1(new_n614), .B2(KEYINPUT97), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n602), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n611), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n593), .B1(new_n610), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT100), .Z(new_n620));
  XOR2_X1   g419(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT101), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n607), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n609), .A3(new_n602), .ZN(new_n625));
  INV_X1    g424(.A(new_n600), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n614), .A2(KEYINPUT97), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n595), .A3(new_n617), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n598), .A2(new_n599), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n625), .A2(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT21), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n252), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n329), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n620), .A2(new_n622), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n623), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n634), .B1(new_n623), .B2(new_n635), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n592), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n633), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n636), .A3(new_n591), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(G232gat), .A2(G233gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(KEYINPUT41), .ZN(new_n645));
  XNOR2_X1  g444(.A(G190gat), .B(G218gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G85gat), .A2(G92gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT7), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT7), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(G85gat), .A3(G92gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G99gat), .A2(G106gat), .ZN(new_n654));
  INV_X1    g453(.A(G92gat), .ZN(new_n655));
  AOI22_X1  g454(.A1(KEYINPUT8), .A2(new_n654), .B1(new_n480), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G99gat), .B(G106gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n653), .B2(new_n656), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n270), .B2(new_n269), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n267), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n270), .A2(new_n661), .B1(KEYINPUT41), .B2(new_n644), .ZN(new_n664));
  XNOR2_X1  g463(.A(G134gat), .B(G162gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT102), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n663), .B2(new_n664), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n648), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n668), .A3(new_n647), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT10), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n659), .A2(new_n660), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n630), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT104), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n630), .A2(new_n681), .A3(new_n678), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n612), .ZN(new_n684));
  NAND2_X1  g483(.A1(KEYINPUT98), .A2(G64gat), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n601), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n602), .B1(new_n686), .B2(KEYINPUT99), .ZN(new_n687));
  INV_X1    g486(.A(new_n609), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n626), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n653), .A2(new_n656), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n657), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G57gat), .B(G64gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n595), .B1(new_n695), .B2(new_n616), .ZN(new_n696));
  INV_X1    g495(.A(new_n617), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n629), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n690), .A2(new_n691), .A3(new_n657), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n689), .A2(new_n694), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n661), .B1(new_n610), .B2(new_n618), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n680), .A2(new_n682), .B1(new_n702), .B2(new_n677), .ZN(new_n703));
  INV_X1    g502(.A(G230gat), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n409), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n676), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n705), .ZN(new_n707));
  INV_X1    g506(.A(new_n660), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(KEYINPUT10), .A3(new_n658), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n709), .A2(new_n610), .A3(new_n618), .A4(KEYINPUT104), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n681), .B1(new_n630), .B2(new_n678), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT10), .B1(new_n700), .B2(new_n701), .ZN(new_n713));
  OAI211_X1 g512(.A(KEYINPUT105), .B(new_n707), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n702), .A2(new_n707), .ZN(new_n715));
  XNOR2_X1  g514(.A(G120gat), .B(G148gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G176gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G204gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n706), .A2(new_n714), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n703), .A2(new_n705), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n718), .B1(new_n721), .B2(new_n715), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n643), .A2(new_n675), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n587), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n493), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n237), .ZN(G1324gat));
  NOR2_X1   g528(.A1(new_n727), .A2(new_n436), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT16), .B(G8gat), .Z(new_n731));
  AND2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n732), .A2(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(KEYINPUT42), .ZN(new_n734));
  OAI21_X1  g533(.A(G8gat), .B1(new_n727), .B2(new_n436), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(G1325gat));
  OAI21_X1  g535(.A(G15gat), .B1(new_n727), .B2(new_n393), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n584), .A2(new_n244), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n727), .B2(new_n738), .ZN(G1326gat));
  NOR2_X1   g538(.A1(new_n727), .A2(new_n578), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT43), .B(G22gat), .Z(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1327gat));
  INV_X1    g541(.A(new_n643), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n724), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n675), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n587), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n207), .A3(new_n579), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT45), .ZN(new_n748));
  INV_X1    g547(.A(new_n578), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n749), .A2(new_n494), .B1(new_n389), .B2(new_n392), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n572), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n586), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT44), .B1(new_n752), .B2(new_n674), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n675), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n573), .B2(new_n586), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n744), .A2(new_n301), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G29gat), .B1(new_n760), .B2(new_n493), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n748), .A2(new_n761), .ZN(G1328gat));
  AND3_X1   g561(.A1(new_n746), .A2(new_n208), .A3(new_n435), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(G36gat), .B1(new_n760), .B2(new_n436), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(G1329gat));
  INV_X1    g567(.A(KEYINPUT106), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n573), .A2(new_n586), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n755), .ZN(new_n774));
  INV_X1    g573(.A(new_n393), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n750), .A2(new_n572), .B1(new_n582), .B2(new_n585), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n754), .B1(new_n776), .B2(new_n675), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .A4(new_n759), .ZN(new_n778));
  INV_X1    g577(.A(new_n211), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n746), .A2(new_n211), .A3(new_n584), .ZN(new_n781));
  AOI211_X1 g580(.A(new_n771), .B(new_n772), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  AND4_X1   g581(.A1(new_n769), .A2(new_n780), .A3(new_n770), .A4(new_n781), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(G1330gat));
  NAND4_X1  g583(.A1(new_n587), .A2(new_n203), .A3(new_n749), .A4(new_n745), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT48), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(KEYINPUT107), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n774), .A2(new_n749), .A3(new_n777), .A4(new_n759), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n203), .A2(KEYINPUT48), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n758), .A2(KEYINPUT108), .A3(new_n749), .A4(new_n759), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n793), .A3(G50gat), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n790), .B1(new_n796), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g596(.A1(new_n723), .A2(new_n299), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n643), .A2(new_n295), .A3(new_n675), .A4(new_n798), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT109), .Z(new_n800));
  NOR2_X1   g599(.A1(new_n776), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n579), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g602(.A(new_n436), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT110), .Z(new_n806));
  NOR2_X1   g605(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(G1333gat));
  AOI21_X1  g607(.A(new_n596), .B1(new_n801), .B2(new_n775), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n390), .A2(G71gat), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n801), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g611(.A1(new_n801), .A2(new_n749), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g613(.A1(new_n643), .A2(new_n300), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n723), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT111), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n758), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G85gat), .B1(new_n818), .B2(new_n493), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n675), .B1(new_n751), .B2(new_n586), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n820), .A2(KEYINPUT51), .A3(new_n815), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT51), .B1(new_n820), .B2(new_n815), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n723), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n579), .A2(new_n480), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n819), .B1(new_n823), .B2(new_n824), .ZN(G1336gat));
  NAND4_X1  g624(.A1(new_n774), .A2(new_n435), .A3(new_n777), .A4(new_n817), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G92gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n436), .A2(G92gat), .A3(new_n724), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT112), .Z(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n821), .B2(new_n822), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n827), .A2(new_n830), .A3(KEYINPUT52), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n758), .A2(KEYINPUT113), .A3(new_n435), .A4(new_n817), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n834), .A3(G92gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n828), .B1(new_n821), .B2(new_n822), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n831), .B1(new_n837), .B2(new_n838), .ZN(G1337gat));
  NOR2_X1   g638(.A1(new_n818), .A2(new_n393), .ZN(new_n840));
  XNOR2_X1  g639(.A(KEYINPUT114), .B(G99gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n584), .A2(new_n841), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n840), .A2(new_n841), .B1(new_n823), .B2(new_n842), .ZN(G1338gat));
  NAND4_X1  g642(.A1(new_n774), .A2(new_n749), .A3(new_n777), .A4(new_n817), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(G106gat), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n578), .A2(G106gat), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n723), .B(new_n846), .C1(new_n821), .C2(new_n822), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g648(.A1(new_n725), .A2(new_n300), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n267), .A2(new_n271), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n202), .B1(new_n852), .B2(new_n276), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n278), .A2(new_n273), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n292), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT115), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n267), .A2(new_n271), .B1(new_n270), .B2(new_n268), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n857), .A2(new_n202), .B1(new_n273), .B2(new_n278), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n859), .A3(new_n292), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n674), .A2(new_n861), .A3(new_n299), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n863), .B1(new_n703), .B2(new_n705), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n706), .A2(new_n864), .A3(new_n714), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n863), .B(new_n707), .C1(new_n712), .C2(new_n713), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(new_n718), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT55), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n866), .A2(KEYINPUT55), .A3(new_n718), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n720), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n862), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n858), .A2(new_n859), .A3(new_n292), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n859), .B1(new_n858), .B2(new_n292), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n723), .B(new_n299), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT116), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n706), .A2(new_n714), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n877), .A2(new_n719), .B1(new_n865), .B2(new_n869), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n865), .A2(new_n867), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT55), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n300), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n861), .A2(new_n883), .A3(new_n299), .A4(new_n723), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n876), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n872), .B1(new_n675), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n851), .B1(new_n886), .B2(new_n643), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(new_n579), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n577), .A2(new_n578), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n436), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n337), .B1(new_n891), .B2(new_n301), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n887), .A2(new_n578), .A3(new_n584), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n493), .A2(new_n435), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(G113gat), .A3(new_n300), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT117), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT117), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n892), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1340gat));
  NAND2_X1  g699(.A1(new_n893), .A2(new_n894), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(new_n338), .A3(new_n724), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n890), .A2(new_n436), .A3(new_n723), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n338), .ZN(G1341gat));
  OAI21_X1  g703(.A(G127gat), .B1(new_n901), .B2(new_n743), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n743), .A2(G127gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n891), .B2(new_n906), .ZN(G1342gat));
  INV_X1    g706(.A(G134gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n436), .A2(new_n674), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT118), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n890), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT56), .Z(new_n913));
  OAI21_X1  g712(.A(G134gat), .B1(new_n901), .B2(new_n675), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT119), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1343gat));
  AND3_X1   g715(.A1(new_n393), .A2(KEYINPUT121), .A3(new_n749), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT121), .B1(new_n393), .B2(new_n749), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n919), .A2(new_n579), .A3(new_n436), .A4(new_n887), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n300), .A2(new_n447), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n871), .A2(new_n868), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n924), .A2(new_n299), .A3(new_n674), .A4(new_n861), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n924), .A2(new_n300), .B1(new_n798), .B2(new_n861), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n674), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n850), .B1(new_n927), .B2(new_n743), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT57), .B1(new_n928), .B2(new_n578), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT57), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n885), .A2(new_n675), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n643), .B1(new_n931), .B2(new_n925), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n930), .B(new_n749), .C1(new_n932), .C2(new_n850), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n393), .A2(new_n894), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n929), .A2(new_n933), .A3(new_n300), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G141gat), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n923), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n922), .B1(new_n936), .B2(KEYINPUT120), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n935), .A2(new_n940), .A3(G141gat), .ZN(new_n941));
  AOI211_X1 g740(.A(KEYINPUT122), .B(new_n937), .C1(new_n939), .C2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n936), .A2(KEYINPUT120), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n941), .A3(new_n923), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n943), .B1(new_n945), .B2(KEYINPUT58), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n938), .B1(new_n942), .B2(new_n946), .ZN(G1344gat));
  INV_X1    g746(.A(new_n920), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n448), .A3(new_n723), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT59), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n930), .B1(new_n887), .B2(new_n749), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n928), .A2(KEYINPUT57), .A3(new_n578), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n723), .A3(new_n934), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n950), .B1(new_n954), .B2(G148gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n929), .A2(new_n933), .A3(new_n934), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(new_n724), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n957), .A2(KEYINPUT59), .A3(new_n448), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n949), .B1(new_n955), .B2(new_n958), .ZN(G1345gat));
  NAND3_X1  g758(.A1(new_n948), .A2(new_n438), .A3(new_n643), .ZN(new_n960));
  OAI21_X1  g759(.A(G155gat), .B1(new_n956), .B2(new_n743), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1346gat));
  OAI21_X1  g761(.A(G162gat), .B1(new_n956), .B2(new_n675), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n888), .A2(new_n439), .A3(new_n911), .A4(new_n919), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1347gat));
  NOR2_X1   g764(.A1(new_n579), .A2(new_n436), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n893), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n967), .A2(new_n312), .A3(new_n301), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n969), .B1(new_n887), .B2(new_n493), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n970), .A2(new_n436), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n887), .A2(new_n969), .A3(new_n493), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n971), .A2(new_n889), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT124), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n971), .A2(new_n975), .A3(new_n889), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(new_n300), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n968), .B1(new_n978), .B2(new_n312), .ZN(G1348gat));
  NAND3_X1  g778(.A1(new_n977), .A2(new_n313), .A3(new_n723), .ZN(new_n980));
  OAI21_X1  g779(.A(G176gat), .B1(new_n967), .B2(new_n724), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1349gat));
  OAI21_X1  g781(.A(G183gat), .B1(new_n967), .B2(new_n743), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n643), .A2(new_n303), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n973), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g785(.A(G190gat), .B1(new_n967), .B2(new_n675), .ZN(new_n987));
  XNOR2_X1  g786(.A(new_n987), .B(KEYINPUT61), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n675), .A2(G190gat), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n989), .B1(new_n977), .B2(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(new_n990), .ZN(new_n992));
  AOI211_X1 g791(.A(KEYINPUT125), .B(new_n992), .C1(new_n974), .C2(new_n976), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n988), .B1(new_n991), .B2(new_n993), .ZN(G1351gat));
  INV_X1    g793(.A(new_n972), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n995), .A2(new_n970), .A3(new_n436), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n775), .A2(new_n578), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(G197gat), .B1(new_n998), .B2(new_n300), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT126), .ZN(new_n1000));
  AND2_X1   g799(.A1(new_n927), .A2(new_n743), .ZN(new_n1001));
  OAI211_X1 g800(.A(new_n930), .B(new_n749), .C1(new_n1001), .C2(new_n850), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n887), .A2(new_n749), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n1000), .B(new_n1002), .C1(new_n1003), .C2(new_n930), .ZN(new_n1004));
  OAI21_X1  g803(.A(KEYINPUT126), .B1(new_n951), .B2(new_n952), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n393), .A2(new_n966), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AND2_X1   g806(.A1(new_n300), .A2(G197gat), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n999), .B1(new_n1007), .B2(new_n1008), .ZN(G1352gat));
  NAND4_X1  g808(.A1(new_n1004), .A2(new_n1005), .A3(new_n723), .A4(new_n1006), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(G204gat), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n724), .A2(G204gat), .ZN(new_n1012));
  NAND4_X1  g811(.A1(new_n971), .A2(new_n997), .A3(new_n972), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT62), .ZN(new_n1015));
  NAND4_X1  g814(.A1(new_n996), .A2(new_n1015), .A3(new_n997), .A4(new_n1012), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1011), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g818(.A1(new_n1011), .A2(KEYINPUT127), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1019), .A2(new_n1020), .ZN(G1353gat));
  NAND3_X1  g820(.A1(new_n953), .A2(new_n643), .A3(new_n1006), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1022), .A2(G211gat), .ZN(new_n1023));
  INV_X1    g822(.A(KEYINPUT63), .ZN(new_n1024));
  XNOR2_X1  g823(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  NAND4_X1  g824(.A1(new_n998), .A2(new_n396), .A3(new_n397), .A4(new_n643), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1025), .A2(new_n1026), .ZN(G1354gat));
  AOI21_X1  g826(.A(G218gat), .B1(new_n998), .B2(new_n674), .ZN(new_n1028));
  NOR2_X1   g827(.A1(new_n675), .A2(new_n403), .ZN(new_n1029));
  AOI21_X1  g828(.A(new_n1028), .B1(new_n1007), .B2(new_n1029), .ZN(G1355gat));
endmodule


