

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U320 ( .A(G99GAT), .B(G85GAT), .Z(n357) );
  NAND2_X1 U321 ( .A1(n418), .A2(n536), .ZN(n419) );
  XOR2_X1 U322 ( .A(G43GAT), .B(KEYINPUT7), .Z(n288) );
  XOR2_X1 U323 ( .A(n440), .B(n375), .Z(n289) );
  INV_X1 U324 ( .A(n554), .ZN(n418) );
  OR2_X1 U325 ( .A1(n420), .A2(n419), .ZN(n421) );
  XNOR2_X1 U326 ( .A(n364), .B(KEYINPUT78), .ZN(n365) );
  XNOR2_X1 U327 ( .A(n366), .B(n365), .ZN(n369) );
  OR2_X1 U328 ( .A1(n580), .A2(n424), .ZN(n462) );
  XNOR2_X1 U329 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U330 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(G127GAT), .B(KEYINPUT95), .Z(n291) );
  XNOR2_X1 U332 ( .A(G71GAT), .B(KEYINPUT65), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n291), .B(n290), .ZN(n304) );
  XOR2_X1 U334 ( .A(G190GAT), .B(G99GAT), .Z(n293) );
  XNOR2_X1 U335 ( .A(G43GAT), .B(G134GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U337 ( .A(G176GAT), .B(G183GAT), .Z(n295) );
  XNOR2_X1 U338 ( .A(KEYINPUT93), .B(KEYINPUT20), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U340 ( .A(n297), .B(n296), .Z(n302) );
  XOR2_X1 U341 ( .A(G113GAT), .B(KEYINPUT0), .Z(n447) );
  XOR2_X1 U342 ( .A(G120GAT), .B(n447), .Z(n299) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U345 ( .A(G15GAT), .B(n300), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT94), .Z(n306) );
  XNOR2_X1 U349 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U351 ( .A(G169GAT), .B(n307), .ZN(n352) );
  XOR2_X1 U352 ( .A(n308), .B(n352), .Z(n559) );
  XOR2_X1 U353 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n310) );
  XNOR2_X1 U354 ( .A(KEYINPUT10), .B(KEYINPUT85), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n310), .B(n309), .ZN(n323) );
  XOR2_X1 U356 ( .A(KEYINPUT11), .B(n357), .Z(n312) );
  XOR2_X1 U357 ( .A(G36GAT), .B(G190GAT), .Z(n347) );
  XNOR2_X1 U358 ( .A(G218GAT), .B(n347), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U360 ( .A(G29GAT), .B(G134GAT), .Z(n440) );
  XNOR2_X1 U361 ( .A(KEYINPUT73), .B(KEYINPUT8), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n288), .B(n313), .ZN(n375) );
  NAND2_X1 U363 ( .A1(G232GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n289), .B(n314), .ZN(n315) );
  XOR2_X1 U365 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U366 ( .A(G50GAT), .B(KEYINPUT83), .Z(n336) );
  XOR2_X1 U367 ( .A(KEYINPUT84), .B(G92GAT), .Z(n318) );
  XNOR2_X1 U368 ( .A(G162GAT), .B(G106GAT), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n336), .B(n319), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X2 U372 ( .A(n323), .B(n322), .Z(n554) );
  NAND2_X1 U373 ( .A1(n559), .A2(n554), .ZN(n455) );
  XOR2_X1 U374 ( .A(KEYINPUT98), .B(KEYINPUT100), .Z(n325) );
  XNOR2_X1 U375 ( .A(KEYINPUT24), .B(KEYINPUT96), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U377 ( .A(KEYINPUT22), .B(KEYINPUT99), .Z(n327) );
  XNOR2_X1 U378 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U380 ( .A(n329), .B(n328), .Z(n341) );
  XNOR2_X1 U381 ( .A(G211GAT), .B(G218GAT), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n330), .B(KEYINPUT21), .ZN(n331) );
  XOR2_X1 U383 ( .A(n331), .B(KEYINPUT97), .Z(n333) );
  XNOR2_X1 U384 ( .A(G197GAT), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n346) );
  XOR2_X1 U386 ( .A(G78GAT), .B(G148GAT), .Z(n335) );
  XNOR2_X1 U387 ( .A(G106GAT), .B(KEYINPUT79), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n367) );
  XOR2_X1 U389 ( .A(n336), .B(n367), .Z(n338) );
  NAND2_X1 U390 ( .A1(G228GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n346), .B(n339), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U394 ( .A(KEYINPUT3), .B(G162GAT), .Z(n343) );
  XNOR2_X1 U395 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U397 ( .A(G141GAT), .B(n344), .ZN(n445) );
  XNOR2_X1 U398 ( .A(n345), .B(n445), .ZN(n473) );
  XOR2_X1 U399 ( .A(n347), .B(n346), .Z(n349) );
  NAND2_X1 U400 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n351) );
  XNOR2_X1 U402 ( .A(G176GAT), .B(G92GAT), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n350), .B(G64GAT), .ZN(n370) );
  XOR2_X1 U404 ( .A(n351), .B(n370), .Z(n356) );
  INV_X1 U405 ( .A(n352), .ZN(n354) );
  XNOR2_X1 U406 ( .A(G8GAT), .B(G183GAT), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n353), .B(KEYINPUT86), .ZN(n415) );
  XNOR2_X1 U408 ( .A(n354), .B(n415), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n520) );
  XOR2_X1 U410 ( .A(KEYINPUT77), .B(n357), .Z(n359) );
  XOR2_X1 U411 ( .A(G120GAT), .B(G57GAT), .Z(n439) );
  XNOR2_X1 U412 ( .A(G204GAT), .B(n439), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U414 ( .A(KEYINPUT81), .B(KEYINPUT33), .Z(n361) );
  XNOR2_X1 U415 ( .A(KEYINPUT80), .B(KEYINPUT31), .ZN(n360) );
  XOR2_X1 U416 ( .A(n361), .B(n360), .Z(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n366) );
  NAND2_X1 U418 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XOR2_X1 U419 ( .A(n367), .B(KEYINPUT32), .Z(n368) );
  XNOR2_X1 U420 ( .A(n369), .B(n368), .ZN(n371) );
  XNOR2_X1 U421 ( .A(n371), .B(n370), .ZN(n373) );
  XNOR2_X1 U422 ( .A(G71GAT), .B(KEYINPUT76), .ZN(n372) );
  XOR2_X1 U423 ( .A(n372), .B(KEYINPUT13), .Z(n414) );
  XNOR2_X1 U424 ( .A(n373), .B(n414), .ZN(n424) );
  INV_X1 U425 ( .A(KEYINPUT41), .ZN(n374) );
  XNOR2_X1 U426 ( .A(n424), .B(n374), .ZN(n506) );
  INV_X1 U427 ( .A(n506), .ZN(n532) );
  XOR2_X1 U428 ( .A(n375), .B(KEYINPUT70), .Z(n377) );
  NAND2_X1 U429 ( .A1(G229GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U431 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n379) );
  XNOR2_X1 U432 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U435 ( .A(G1GAT), .B(G197GAT), .Z(n383) );
  XNOR2_X1 U436 ( .A(G113GAT), .B(G141GAT), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U439 ( .A(G50GAT), .B(G29GAT), .Z(n388) );
  XNOR2_X1 U440 ( .A(G15GAT), .B(G22GAT), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n386), .B(KEYINPUT74), .ZN(n409) );
  XNOR2_X1 U442 ( .A(G36GAT), .B(n409), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U444 ( .A(n390), .B(n389), .Z(n395) );
  XOR2_X1 U445 ( .A(KEYINPUT68), .B(KEYINPUT75), .Z(n392) );
  XNOR2_X1 U446 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U448 ( .A(G169GAT), .B(n393), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n570) );
  NAND2_X1 U450 ( .A1(n532), .A2(n570), .ZN(n397) );
  XOR2_X1 U451 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n420) );
  XOR2_X1 U453 ( .A(KEYINPUT15), .B(G64GAT), .Z(n399) );
  XNOR2_X1 U454 ( .A(G78GAT), .B(G57GAT), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U456 ( .A(KEYINPUT90), .B(KEYINPUT87), .Z(n401) );
  XNOR2_X1 U457 ( .A(KEYINPUT91), .B(KEYINPUT14), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U459 ( .A(n403), .B(n402), .Z(n408) );
  XOR2_X1 U460 ( .A(KEYINPUT89), .B(KEYINPUT12), .Z(n405) );
  NAND2_X1 U461 ( .A1(G231GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U463 ( .A(KEYINPUT88), .B(n406), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n413) );
  XOR2_X1 U465 ( .A(G1GAT), .B(G127GAT), .Z(n436) );
  XOR2_X1 U466 ( .A(n436), .B(G211GAT), .Z(n411) );
  XNOR2_X1 U467 ( .A(n409), .B(G155GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U469 ( .A(n413), .B(n412), .Z(n417) );
  XOR2_X1 U470 ( .A(n415), .B(n414), .Z(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n536) );
  XNOR2_X1 U472 ( .A(n421), .B(KEYINPUT47), .ZN(n428) );
  XNOR2_X1 U473 ( .A(n554), .B(KEYINPUT109), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n422), .B(KEYINPUT36), .ZN(n581) );
  NOR2_X1 U475 ( .A1(n581), .A2(n536), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n423), .B(KEYINPUT45), .ZN(n425) );
  NAND2_X1 U477 ( .A1(n425), .A2(n424), .ZN(n426) );
  NOR2_X1 U478 ( .A1(n426), .A2(n570), .ZN(n427) );
  NOR2_X1 U479 ( .A1(n428), .A2(n427), .ZN(n429) );
  XNOR2_X1 U480 ( .A(KEYINPUT48), .B(n429), .ZN(n527) );
  NOR2_X1 U481 ( .A1(n520), .A2(n527), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n430), .B(KEYINPUT54), .ZN(n452) );
  XOR2_X1 U483 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n432) );
  XNOR2_X1 U484 ( .A(KEYINPUT102), .B(KEYINPUT1), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n451) );
  XOR2_X1 U486 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n434) );
  XNOR2_X1 U487 ( .A(KEYINPUT101), .B(KEYINPUT4), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U489 ( .A(n435), .B(G85GAT), .Z(n438) );
  XNOR2_X1 U490 ( .A(G148GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n444) );
  XOR2_X1 U492 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U493 ( .A1(G225GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U495 ( .A(n444), .B(n443), .Z(n449) );
  INV_X1 U496 ( .A(n445), .ZN(n446) );
  XNOR2_X1 U497 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U498 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U499 ( .A(n451), .B(n450), .Z(n472) );
  XNOR2_X1 U500 ( .A(KEYINPUT105), .B(n472), .ZN(n545) );
  NAND2_X1 U501 ( .A1(n452), .A2(n545), .ZN(n453) );
  XNOR2_X1 U502 ( .A(n453), .B(KEYINPUT64), .ZN(n461) );
  NOR2_X1 U503 ( .A1(n473), .A2(n461), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n454), .B(KEYINPUT55), .ZN(n561) );
  OR2_X1 U505 ( .A1(n455), .A2(n561), .ZN(n459) );
  XOR2_X1 U506 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n457) );
  INV_X1 U507 ( .A(G190GAT), .ZN(n456) );
  INV_X1 U508 ( .A(G204GAT), .ZN(n465) );
  XOR2_X1 U509 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n463) );
  INV_X1 U510 ( .A(n559), .ZN(n557) );
  NAND2_X1 U511 ( .A1(n557), .A2(n473), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT26), .ZN(n466) );
  NOR2_X1 U513 ( .A1(n461), .A2(n466), .ZN(n577) );
  INV_X1 U514 ( .A(n577), .ZN(n580) );
  XNOR2_X1 U515 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U516 ( .A(n465), .B(n464), .ZN(G1353GAT) );
  XNOR2_X1 U517 ( .A(n520), .B(KEYINPUT27), .ZN(n475) );
  NOR2_X1 U518 ( .A1(n466), .A2(n475), .ZN(n546) );
  NOR2_X1 U519 ( .A1(n520), .A2(n557), .ZN(n467) );
  NOR2_X1 U520 ( .A1(n473), .A2(n467), .ZN(n468) );
  XOR2_X1 U521 ( .A(n468), .B(KEYINPUT25), .Z(n469) );
  XNOR2_X1 U522 ( .A(KEYINPUT106), .B(n469), .ZN(n470) );
  NOR2_X1 U523 ( .A1(n546), .A2(n470), .ZN(n471) );
  NOR2_X1 U524 ( .A1(n472), .A2(n471), .ZN(n478) );
  XNOR2_X1 U525 ( .A(n473), .B(KEYINPUT67), .ZN(n474) );
  XNOR2_X1 U526 ( .A(n474), .B(KEYINPUT28), .ZN(n524) );
  NOR2_X1 U527 ( .A1(n545), .A2(n475), .ZN(n476) );
  NAND2_X1 U528 ( .A1(n524), .A2(n476), .ZN(n529) );
  NOR2_X1 U529 ( .A1(n559), .A2(n529), .ZN(n477) );
  NOR2_X1 U530 ( .A1(n478), .A2(n477), .ZN(n492) );
  NOR2_X1 U531 ( .A1(n554), .A2(n536), .ZN(n479) );
  XOR2_X1 U532 ( .A(KEYINPUT92), .B(n479), .Z(n480) );
  XNOR2_X1 U533 ( .A(n480), .B(KEYINPUT16), .ZN(n481) );
  NOR2_X1 U534 ( .A1(n492), .A2(n481), .ZN(n507) );
  NAND2_X1 U535 ( .A1(n424), .A2(n570), .ZN(n482) );
  XOR2_X1 U536 ( .A(KEYINPUT82), .B(n482), .Z(n496) );
  NAND2_X1 U537 ( .A1(n507), .A2(n496), .ZN(n490) );
  NOR2_X1 U538 ( .A1(n545), .A2(n490), .ZN(n483) );
  XOR2_X1 U539 ( .A(KEYINPUT34), .B(n483), .Z(n484) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NOR2_X1 U541 ( .A1(n520), .A2(n490), .ZN(n485) );
  XOR2_X1 U542 ( .A(G8GAT), .B(n485), .Z(G1325GAT) );
  NOR2_X1 U543 ( .A1(n490), .A2(n557), .ZN(n489) );
  XOR2_X1 U544 ( .A(KEYINPUT107), .B(KEYINPUT35), .Z(n487) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT108), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n524), .A2(n490), .ZN(n491) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n491), .Z(G1327GAT) );
  NOR2_X1 U550 ( .A1(n581), .A2(n492), .ZN(n493) );
  NAND2_X1 U551 ( .A1(n536), .A2(n493), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT37), .B(n494), .ZN(n495) );
  XNOR2_X1 U553 ( .A(KEYINPUT110), .B(n495), .ZN(n517) );
  NAND2_X1 U554 ( .A1(n496), .A2(n517), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(KEYINPUT38), .ZN(n503) );
  NOR2_X1 U556 ( .A1(n503), .A2(n545), .ZN(n499) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n520), .A2(n503), .ZN(n500) );
  XOR2_X1 U560 ( .A(G36GAT), .B(n500), .Z(G1329GAT) );
  NOR2_X1 U561 ( .A1(n503), .A2(n557), .ZN(n501) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(n501), .Z(n502) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT111), .ZN(n505) );
  NOR2_X1 U565 ( .A1(n524), .A2(n503), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  NOR2_X1 U567 ( .A1(n570), .A2(n506), .ZN(n518) );
  NAND2_X1 U568 ( .A1(n518), .A2(n507), .ZN(n513) );
  NOR2_X1 U569 ( .A1(n545), .A2(n513), .ZN(n508) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n508), .Z(n509) );
  XNOR2_X1 U571 ( .A(KEYINPUT42), .B(n509), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n520), .A2(n513), .ZN(n510) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n510), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n557), .A2(n513), .ZN(n511) );
  XOR2_X1 U575 ( .A(KEYINPUT112), .B(n511), .Z(n512) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n512), .ZN(G1334GAT) );
  NOR2_X1 U577 ( .A1(n524), .A2(n513), .ZN(n515) );
  XNOR2_X1 U578 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U580 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  NAND2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n523) );
  NOR2_X1 U582 ( .A1(n545), .A2(n523), .ZN(n519) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n519), .Z(G1336GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n523), .ZN(n521) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n521), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n557), .A2(n523), .ZN(n522) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n522), .Z(G1338GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(n525), .Z(n526) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U591 ( .A(G113GAT), .B(KEYINPUT115), .Z(n531) );
  OR2_X1 U592 ( .A1(n557), .A2(n527), .ZN(n528) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n540), .A2(n570), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U597 ( .A1(n540), .A2(n532), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(n535), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n538) );
  INV_X1 U601 ( .A(n536), .ZN(n578) );
  NAND2_X1 U602 ( .A1(n540), .A2(n578), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U606 ( .A1(n540), .A2(n554), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT119), .Z(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NOR2_X1 U610 ( .A1(n545), .A2(n527), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U612 ( .A(KEYINPUT120), .B(n548), .Z(n555) );
  NAND2_X1 U613 ( .A1(n555), .A2(n570), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U616 ( .A1(n532), .A2(n555), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n555), .A2(n578), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n561), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n570), .A2(n568), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n559), .A2(n532), .ZN(n560) );
  OR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n567) );
  XOR2_X1 U630 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n578), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n574) );
  INV_X1 U639 ( .A(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U645 ( .A(KEYINPUT62), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

