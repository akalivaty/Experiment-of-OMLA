//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(G107), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n194), .A2(new_n197), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n196), .A2(G104), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n193), .A2(G107), .ZN(new_n202));
  OAI21_X1  g016(.A(G101), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  AND4_X1   g022(.A1(new_n204), .A2(new_n206), .A3(new_n208), .A4(G128), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n207), .B(G146), .C1(new_n210), .C2(KEYINPUT1), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n205), .A3(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n200), .B(new_n203), .C1(new_n209), .C2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n204), .A3(G128), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n211), .A2(KEYINPUT66), .A3(new_n212), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT66), .B1(new_n211), .B2(new_n212), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n200), .A2(new_n203), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n214), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT11), .ZN(new_n223));
  INV_X1    g037(.A(G137), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(G134), .ZN(new_n225));
  INV_X1    g039(.A(G134), .ZN(new_n226));
  OAI22_X1  g040(.A1(new_n226), .A2(G137), .B1(KEYINPUT65), .B2(KEYINPUT11), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n224), .B2(G134), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n229), .B1(new_n228), .B2(new_n232), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n221), .A2(KEYINPUT12), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT12), .B1(new_n221), .B2(new_n235), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n194), .A2(new_n197), .A3(new_n199), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(G101), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT79), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n239), .A2(KEYINPUT79), .A3(new_n240), .A4(G101), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n215), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n206), .A2(new_n208), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT0), .B(G128), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT64), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n239), .A2(G101), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT4), .A3(new_n200), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n245), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n235), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT10), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n214), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n219), .A2(KEYINPUT10), .A3(new_n220), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n255), .A2(new_n256), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n192), .B1(new_n238), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n255), .A2(new_n258), .A3(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n235), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n260), .A3(new_n191), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G902), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n187), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n260), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n192), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n260), .A2(new_n191), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n271), .A2(new_n238), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT80), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n273), .A2(new_n274), .A3(new_n187), .A4(new_n267), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n191), .B1(new_n264), .B2(new_n260), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n271), .A2(new_n238), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n187), .B(new_n267), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT80), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n268), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G221), .ZN(new_n281));
  XOR2_X1   g095(.A(KEYINPUT9), .B(G234), .Z(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(new_n267), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n189), .A2(G952), .ZN(new_n285));
  NAND2_X1  g099(.A1(G234), .A2(G237), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT21), .B(G898), .Z(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(G902), .A3(G953), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G214), .B1(G237), .B2(G902), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(G110), .B(G122), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT82), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT84), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n294), .B(KEYINPUT82), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT84), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT8), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n297), .A3(KEYINPUT8), .ZN(new_n304));
  XNOR2_X1  g118(.A(G116), .B(G119), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT5), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT5), .ZN(new_n307));
  INV_X1    g121(.A(G119), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(G116), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(G113), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G113), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT2), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G113), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n315), .A2(new_n305), .A3(KEYINPUT67), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT67), .B1(new_n315), .B2(new_n305), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n310), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n220), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n317), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n315), .A2(new_n305), .A3(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n220), .B1(new_n323), .B2(new_n310), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n303), .B(new_n304), .C1(new_n320), .C2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n219), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n252), .A2(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G224), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G953), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT85), .ZN(new_n334));
  OAI22_X1  g148(.A1(new_n316), .A2(new_n317), .B1(new_n305), .B2(new_n315), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n245), .A2(new_n335), .A3(new_n254), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT81), .B1(new_n318), .B2(new_n319), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n323), .A2(new_n338), .A3(new_n220), .A4(new_n310), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n336), .A2(new_n337), .A3(new_n296), .A4(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT85), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n329), .A2(new_n341), .A3(KEYINPUT7), .A4(new_n332), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n325), .A2(new_n334), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n329), .B1(KEYINPUT7), .B2(new_n332), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n267), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n298), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT6), .A4(new_n340), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n347), .A2(KEYINPUT6), .A3(new_n340), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n346), .A2(new_n351), .A3(new_n298), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT83), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n349), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n329), .B(new_n331), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n345), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT86), .ZN(new_n358));
  OAI21_X1  g172(.A(G210), .B1(G237), .B2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n347), .A2(KEYINPUT6), .A3(new_n340), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT83), .A3(new_n352), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n355), .B1(new_n363), .B2(new_n349), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n361), .B1(new_n364), .B2(new_n345), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n358), .A2(new_n360), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n357), .A2(new_n359), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT87), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n354), .A2(new_n356), .ZN(new_n370));
  INV_X1    g184(.A(new_n345), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n359), .B1(new_n372), .B2(new_n361), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n369), .B1(new_n373), .B2(new_n358), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n284), .B(new_n293), .C1(new_n368), .C2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n252), .B1(new_n233), .B2(new_n234), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n226), .A2(G137), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n224), .A2(G134), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n229), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n231), .B1(new_n227), .B2(new_n225), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n381), .B2(new_n229), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n219), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n377), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n384), .B1(new_n377), .B2(new_n383), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n335), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n315), .A2(new_n305), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n321), .B2(new_n322), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n377), .A2(new_n383), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(G101), .ZN(new_n392));
  INV_X1    g206(.A(G237), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n189), .A3(G210), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n392), .B(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n387), .A2(KEYINPUT31), .A3(new_n390), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n267), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n387), .A2(new_n390), .A3(new_n395), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n377), .A2(new_n383), .A3(new_n389), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n389), .B1(new_n377), .B2(new_n383), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT28), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT28), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n390), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n395), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT31), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n397), .B1(new_n398), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT32), .ZN(new_n408));
  INV_X1    g222(.A(G472), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n396), .A2(new_n267), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n377), .A2(new_n383), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n335), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n402), .B1(new_n413), .B2(new_n390), .ZN(new_n414));
  INV_X1    g228(.A(new_n403), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n405), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT31), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n398), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n411), .A2(new_n418), .A3(new_n409), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT32), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n410), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n387), .A2(new_n390), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(new_n395), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n401), .A2(new_n395), .A3(new_n403), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n267), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n425), .A2(new_n426), .ZN(new_n429));
  OAI21_X1  g243(.A(G472), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n421), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(KEYINPUT72), .A2(G125), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT73), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n433), .A3(G140), .ZN(new_n434));
  INV_X1    g248(.A(G140), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT73), .B1(new_n435), .B2(G125), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(KEYINPUT72), .A3(G125), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT16), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT16), .B1(new_n435), .B2(G125), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n205), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(KEYINPUT24), .A2(G110), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT24), .A2(G110), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(KEYINPUT69), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT69), .ZN(new_n447));
  INV_X1    g261(.A(new_n445), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n448), .B2(new_n443), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G119), .B(G128), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT71), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT23), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n308), .B2(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n308), .A2(G128), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT71), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n457), .A2(new_n210), .A3(KEYINPUT23), .A4(G119), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n453), .A2(new_n455), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  OAI22_X1  g273(.A1(new_n450), .A2(new_n451), .B1(new_n459), .B2(G110), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT75), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n442), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n326), .A2(G140), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n435), .A2(G125), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n205), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT76), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n462), .B(new_n466), .C1(new_n461), .C2(new_n460), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n439), .A2(new_n441), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G146), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n440), .B1(new_n438), .B2(KEYINPUT16), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n205), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n469), .A2(new_n471), .B1(G110), .B2(new_n459), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n446), .A2(new_n449), .A3(new_n451), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n446), .A2(new_n449), .A3(KEYINPUT70), .A4(new_n451), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT74), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n459), .A2(G110), .ZN(new_n479));
  AOI211_X1 g293(.A(G146), .B(new_n440), .C1(new_n438), .C2(KEYINPUT16), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n442), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n477), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n467), .B1(new_n478), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT22), .B(G137), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT77), .ZN(new_n487));
  INV_X1    g301(.A(G234), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n281), .A2(new_n488), .A3(G953), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n487), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n467), .B(new_n490), .C1(new_n478), .C2(new_n484), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n267), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n497));
  INV_X1    g311(.A(new_n495), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n492), .A2(new_n267), .A3(new_n493), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G217), .B1(new_n488), .B2(G902), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT68), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n492), .A2(new_n493), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(G902), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n500), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n431), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G122), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT94), .B1(new_n507), .B2(G116), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n509));
  INV_X1    g323(.A(G116), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(G122), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n510), .A2(G122), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n512), .A2(G107), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n513), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT14), .ZN(new_n516));
  OAI211_X1 g330(.A(KEYINPUT96), .B(new_n515), .C1(new_n512), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n512), .A2(new_n516), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT96), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n516), .B1(new_n508), .B2(new_n511), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n519), .B1(new_n520), .B2(new_n513), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n514), .B1(new_n522), .B2(G107), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n207), .A2(G128), .ZN(new_n524));
  OR3_X1    g338(.A1(new_n210), .A2(KEYINPUT95), .A3(G143), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT95), .B1(new_n210), .B2(G143), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n226), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n524), .A2(KEYINPUT13), .ZN(new_n530));
  OR3_X1    g344(.A1(new_n527), .A2(new_n226), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n527), .B1(new_n226), .B2(new_n530), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n512), .A2(new_n513), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(new_n196), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n531), .B(new_n532), .C1(new_n514), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n282), .ZN(new_n536));
  INV_X1    g350(.A(G217), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n536), .A2(new_n537), .A3(G953), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n529), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n538), .B1(new_n529), .B2(new_n535), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n267), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G478), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n542), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT20), .ZN(new_n547));
  XNOR2_X1  g361(.A(G113), .B(G122), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(new_n193), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n438), .A2(KEYINPUT19), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT19), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n463), .A2(new_n464), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n550), .A2(new_n205), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT91), .B1(new_n553), .B2(new_n442), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n393), .A2(new_n189), .A3(G214), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n207), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n393), .A2(new_n189), .A3(G143), .A4(G214), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n555), .B1(new_n559), .B2(new_n229), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT89), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n561), .A3(new_n229), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n557), .A2(new_n558), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT90), .A3(G131), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT89), .B1(new_n563), .B2(G131), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n560), .A2(new_n562), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n550), .A2(new_n205), .A3(new_n552), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n567), .B(new_n568), .C1(new_n205), .C2(new_n470), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n554), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n438), .A2(G146), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n466), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n563), .A2(KEYINPUT88), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT18), .A3(G131), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(KEYINPUT18), .B2(G131), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT92), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n549), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n570), .A2(new_n577), .A3(KEYINPUT92), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n469), .A2(KEYINPUT93), .A3(new_n471), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT93), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n442), .B2(new_n480), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT90), .B1(new_n563), .B2(G131), .ZN(new_n585));
  AOI211_X1 g399(.A(new_n555), .B(new_n229), .C1(new_n557), .C2(new_n558), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT17), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n582), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n585), .A2(new_n586), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n565), .A4(new_n562), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n575), .A2(new_n576), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n588), .A2(new_n591), .B1(new_n572), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n580), .A2(new_n581), .B1(new_n593), .B2(new_n549), .ZN(new_n594));
  NOR2_X1   g408(.A1(G475), .A2(G902), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n547), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n591), .A2(new_n584), .A3(new_n582), .A4(new_n587), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n598), .A2(new_n549), .A3(new_n577), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n549), .B1(new_n598), .B2(new_n577), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n267), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G475), .ZN(new_n602));
  INV_X1    g416(.A(new_n581), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT92), .B1(new_n570), .B2(new_n577), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n603), .A2(new_n604), .A3(new_n549), .ZN(new_n605));
  OAI211_X1 g419(.A(KEYINPUT20), .B(new_n595), .C1(new_n605), .C2(new_n599), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n546), .A2(new_n597), .A3(new_n602), .A4(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n376), .A2(new_n506), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  NAND2_X1  g424(.A1(new_n411), .A2(new_n418), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G472), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n612), .A2(new_n419), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n505), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n614), .A2(new_n283), .A3(new_n280), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n360), .B1(new_n364), .B2(new_n345), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n292), .B1(new_n367), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n597), .A2(new_n602), .A3(new_n606), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT33), .B1(new_n540), .B2(new_n541), .ZN(new_n620));
  INV_X1    g434(.A(new_n541), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n539), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n620), .A2(new_n623), .A3(G478), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n543), .B(new_n267), .C1(new_n540), .C2(new_n541), .ZN(new_n625));
  NAND2_X1  g439(.A1(G478), .A2(G902), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n618), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n615), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  NOR2_X1   g446(.A1(new_n619), .A2(new_n546), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n615), .A2(new_n617), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT35), .B(G107), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT97), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n634), .B(new_n636), .ZN(G9));
  NAND2_X1  g451(.A1(new_n612), .A2(new_n419), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n500), .A2(new_n502), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n485), .A2(KEYINPUT98), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n491), .A2(KEYINPUT36), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n485), .A2(KEYINPUT98), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n504), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n638), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n376), .A2(new_n608), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G110), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT99), .B(KEYINPUT37), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  NAND2_X1  g464(.A1(new_n639), .A2(new_n645), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n651), .A2(new_n431), .A3(new_n284), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n289), .A2(G900), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n287), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n619), .A2(new_n546), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n291), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n367), .B2(new_n616), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n659), .B1(new_n656), .B2(new_n658), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n652), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  NAND2_X1  g477(.A1(new_n366), .A2(KEYINPUT87), .ZN(new_n664));
  INV_X1    g478(.A(new_n367), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n373), .B2(new_n358), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n664), .B1(new_n666), .B2(KEYINPUT87), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT38), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT38), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n423), .A2(new_n405), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n399), .A2(new_n400), .ZN(new_n672));
  AOI21_X1  g486(.A(G902), .B1(new_n672), .B2(new_n405), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n421), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n542), .B(new_n544), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n619), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n654), .B(KEYINPUT39), .Z(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n284), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n657), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n670), .A2(new_n676), .A3(new_n679), .A4(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n651), .B1(new_n682), .B2(KEYINPUT40), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n207), .ZN(G45));
  AND3_X1   g504(.A1(new_n619), .A2(new_n627), .A3(new_n654), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n652), .A2(new_n658), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  NAND2_X1  g507(.A1(new_n275), .A2(new_n279), .ZN(new_n694));
  INV_X1    g508(.A(new_n283), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n273), .A2(new_n267), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n431), .A2(new_n698), .A3(new_n505), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n629), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  AND4_X1   g516(.A1(new_n431), .A2(new_n698), .A3(new_n505), .A4(new_n633), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n617), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT101), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n510), .ZN(G18));
  AND3_X1   g520(.A1(new_n651), .A2(new_n698), .A3(new_n658), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n431), .A2(new_n608), .A3(new_n290), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  NAND3_X1  g524(.A1(new_n617), .A2(new_n505), .A3(new_n613), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n275), .A2(new_n279), .B1(new_n696), .B2(G469), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n677), .A3(new_n619), .A4(new_n695), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT102), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n503), .A2(new_n504), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n613), .A2(new_n639), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n678), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n718), .A3(new_n719), .A4(new_n617), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  AND2_X1   g536(.A1(new_n646), .A2(new_n691), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n367), .A2(new_n616), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n291), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n717), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  INV_X1    g542(.A(new_n268), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n694), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT103), .B1(new_n730), .B2(new_n695), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT103), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n280), .A2(new_n732), .A3(new_n283), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n408), .B1(new_n407), .B2(new_n409), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n408), .A2(new_n411), .A3(new_n418), .A4(new_n409), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT104), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n410), .A2(new_n420), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n430), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n734), .A2(KEYINPUT42), .A3(new_n505), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n366), .A2(new_n367), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n369), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n291), .A3(new_n664), .A4(new_n691), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT105), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n740), .A2(new_n505), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n730), .A2(KEYINPUT103), .A3(new_n695), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n732), .B1(new_n280), .B2(new_n283), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n748), .A3(KEYINPUT42), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n368), .A2(new_n374), .A3(new_n657), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n691), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n506), .A3(new_n691), .A4(new_n734), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n745), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n229), .ZN(G33));
  AND4_X1   g571(.A1(new_n506), .A2(new_n752), .A3(new_n656), .A4(new_n734), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT106), .B(G134), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G36));
  AND3_X1   g574(.A1(new_n597), .A2(new_n602), .A3(new_n606), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n627), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(KEYINPUT44), .A3(new_n638), .A4(new_n651), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT109), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n766), .A2(new_n657), .A3(new_n667), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n266), .B(KEYINPUT45), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(G469), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n187), .A2(new_n267), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT46), .ZN(new_n775));
  INV_X1    g589(.A(new_n769), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n776), .B2(new_n770), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n769), .A2(KEYINPUT107), .A3(KEYINPUT46), .A4(new_n771), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n777), .A3(new_n694), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n695), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n780), .A2(KEYINPUT108), .A3(new_n680), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n764), .A2(new_n638), .A3(new_n651), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT108), .B1(new_n780), .B2(new_n680), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n767), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n779), .A2(new_n695), .B1(KEYINPUT110), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(KEYINPUT110), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n744), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n780), .A2(new_n791), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n431), .A2(new_n505), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NOR2_X1   g612(.A1(new_n762), .A2(new_n657), .ZN(new_n799));
  INV_X1    g613(.A(new_n712), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT49), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n799), .A2(new_n505), .A3(new_n695), .A4(new_n801), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT111), .Z(new_n803));
  NOR2_X1   g617(.A1(new_n800), .A2(KEYINPUT49), .ZN(new_n804));
  OR4_X1    g618(.A1(new_n676), .A2(new_n803), .A3(new_n670), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n628), .A2(KEYINPUT112), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n619), .A2(new_n627), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n809), .B(new_n293), .C1(new_n368), .C2(new_n374), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT113), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n667), .A2(new_n812), .A3(new_n293), .A4(new_n809), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n813), .A3(new_n615), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n667), .A2(new_n615), .A3(new_n293), .A4(new_n633), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n609), .A2(new_n814), .A3(new_n647), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n607), .B2(new_n655), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n761), .A2(KEYINPUT114), .A3(new_n546), .A4(new_n654), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n651), .A2(new_n431), .A3(new_n284), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n646), .A2(new_n747), .A3(new_n748), .A4(new_n691), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n752), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n714), .A2(new_n720), .B1(new_n703), .B2(new_n617), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n629), .A2(new_n699), .B1(new_n707), .B2(new_n708), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n725), .A2(new_n678), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n654), .A2(KEYINPUT115), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n651), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n654), .A2(KEYINPUT115), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n280), .A2(new_n283), .A3(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n828), .A2(new_n676), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n662), .A2(new_n692), .A3(new_n727), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n821), .A2(new_n725), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n837), .A2(new_n691), .B1(new_n723), .B2(new_n726), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(KEYINPUT52), .A3(new_n662), .A4(new_n833), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n827), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n745), .A2(new_n753), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n754), .A2(new_n755), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n758), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n816), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n816), .A2(new_n840), .A3(new_n843), .A4(KEYINPUT53), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n846), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT54), .B1(new_n846), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n668), .A2(new_n669), .A3(new_n698), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n287), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n764), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n764), .A2(KEYINPUT116), .A3(new_n854), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n614), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n853), .A2(new_n859), .A3(new_n657), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT50), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n853), .A2(new_n859), .A3(KEYINPUT50), .A4(new_n657), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n752), .A2(new_n698), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n857), .B2(new_n858), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n646), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n505), .A2(new_n854), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n865), .A2(new_n676), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n627), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n761), .A3(new_n870), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n792), .A2(new_n794), .B1(new_n283), .B2(new_n712), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n859), .A2(new_n752), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n867), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n851), .B1(new_n864), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n869), .A2(new_n619), .A3(new_n627), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT48), .ZN(new_n877));
  INV_X1    g691(.A(new_n746), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n866), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n866), .B2(new_n878), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n285), .B(new_n876), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n726), .B2(new_n859), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n872), .A2(new_n873), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n862), .A2(new_n863), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n867), .A2(new_n871), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT51), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n875), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n850), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n805), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(KEYINPUT117), .B(new_n805), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(G75));
  AOI21_X1  g708(.A(new_n267), .B1(new_n846), .B2(new_n847), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(G210), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n354), .B(new_n355), .ZN(new_n898));
  XNOR2_X1  g712(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n189), .A2(G952), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G51));
  XNOR2_X1  g718(.A(new_n770), .B(KEYINPUT57), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n850), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n273), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n895), .A2(new_n776), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(G54));
  NAND3_X1  g723(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n910), .A2(new_n594), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n594), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n911), .A2(new_n912), .A3(new_n903), .ZN(G60));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n620), .A2(new_n623), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n626), .B(KEYINPUT59), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n850), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n814), .A2(new_n609), .A3(new_n647), .A4(new_n815), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n919), .A2(new_n756), .A3(new_n758), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT53), .B1(new_n920), .B2(new_n840), .ZN(new_n921));
  AND4_X1   g735(.A1(KEYINPUT53), .A2(new_n816), .A3(new_n840), .A4(new_n843), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n846), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n924), .A3(new_n916), .ZN(new_n925));
  INV_X1    g739(.A(new_n915), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n903), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n923), .A2(new_n915), .A3(new_n924), .A4(new_n916), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT119), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n917), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n917), .A2(new_n927), .A3(KEYINPUT120), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(G63));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n643), .A2(new_n644), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n537), .A2(new_n267), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n936), .B(new_n939), .C1(new_n921), .C2(new_n922), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n939), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n846), .B2(new_n847), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(KEYINPUT122), .A3(new_n936), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n935), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n903), .B1(new_n942), .B2(new_n945), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n944), .A2(new_n503), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n949), .B(new_n948), .C1(new_n946), .C2(KEYINPUT61), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(G66));
  AOI21_X1  g767(.A(new_n189), .B1(new_n288), .B2(G224), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n825), .A2(new_n826), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n816), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n954), .B1(new_n956), .B2(new_n189), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n363), .B(new_n349), .C1(G898), .C2(new_n189), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n957), .B(new_n958), .Z(G69));
  NOR2_X1   g773(.A1(new_n385), .A2(new_n386), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n550), .A2(new_n552), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(G900), .A2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n838), .A2(new_n662), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT124), .Z(new_n965));
  AND2_X1   g779(.A1(new_n965), .A2(new_n843), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n781), .A2(new_n878), .A3(new_n785), .A4(new_n828), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n966), .A2(new_n787), .A3(new_n797), .A4(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n962), .B(new_n963), .C1(new_n968), .C2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n787), .A2(new_n797), .ZN(new_n970));
  INV_X1    g784(.A(new_n689), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n965), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n971), .A2(new_n965), .A3(KEYINPUT62), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n809), .A2(new_n633), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n752), .A3(new_n506), .A4(new_n683), .ZN(new_n978));
  AOI21_X1  g792(.A(G953), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n969), .B1(new_n979), .B2(new_n962), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n969), .B2(KEYINPUT125), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  OAI221_X1 g797(.A(new_n969), .B1(KEYINPUT125), .B2(new_n981), .C1(new_n979), .C2(new_n962), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(G72));
  INV_X1    g799(.A(new_n671), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n976), .A2(new_n955), .A3(new_n816), .A4(new_n978), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  AOI21_X1  g803(.A(new_n986), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n989), .B1(new_n968), .B2(new_n956), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n423), .A2(new_n405), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT126), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n986), .A2(new_n992), .A3(new_n989), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n846), .B2(new_n847), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n990), .A2(new_n994), .A3(new_n903), .A4(new_n997), .ZN(G57));
endmodule


