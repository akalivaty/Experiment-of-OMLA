//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1135, new_n1136;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(G234));
  NAND2_X1  g027(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(new_n457), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT69), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT70), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  OAI211_X1 g054(.A(G137), .B(new_n476), .C1(new_n467), .C2(new_n468), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n472), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OR3_X1    g057(.A1(new_n469), .A2(KEYINPUT71), .A3(new_n476), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT71), .B1(new_n469), .B2(new_n476), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n469), .A2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G136), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n469), .A2(new_n476), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G126), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n467), .B2(new_n468), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n501), .B(KEYINPUT72), .C1(new_n468), .C2(new_n467), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT4), .A4(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT74), .A2(KEYINPUT4), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT74), .A2(KEYINPUT4), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT75), .B1(new_n502), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n476), .A2(G138), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n507), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n520), .B1(new_n502), .B2(new_n503), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n505), .B1(new_n521), .B2(new_n506), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n499), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(G164));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(new_n527), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT5), .B(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n529), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n534), .A2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n531), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G51), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT5), .B(G543), .Z(new_n545));
  NAND2_X1  g120(.A1(new_n531), .A2(G89), .ZN(new_n546));
  NAND2_X1  g121(.A1(G63), .A2(G651), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n544), .A2(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  NAND2_X1  g125(.A1(new_n528), .A2(G52), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(new_n533), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n536), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n553), .A2(new_n555), .ZN(G171));
  NAND2_X1  g131(.A1(new_n528), .A2(G43), .ZN(new_n557));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n558), .B2(new_n533), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n532), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n536), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(KEYINPUT9), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n528), .A2(new_n573), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n574), .A2(new_n572), .A3(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n545), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n533), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n578), .A2(G651), .B1(new_n579), .B2(G91), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n574), .B1(new_n572), .B2(KEYINPUT9), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  OAI21_X1  g158(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n579), .A2(G87), .B1(G49), .B2(new_n528), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n545), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G48), .B2(new_n528), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n533), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n533), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT79), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n592), .A2(new_n595), .A3(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n579), .A2(G85), .B1(G47), .B2(new_n528), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n536), .B2(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n531), .A2(new_n532), .A3(G92), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n532), .A2(G66), .ZN(new_n605));
  INV_X1    g180(.A(G79), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT80), .B1(new_n606), .B2(new_n525), .ZN(new_n607));
  OR3_X1    g182(.A1(new_n606), .A2(new_n525), .A3(KEYINPUT80), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n602), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n602), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT81), .ZN(G148));
  NAND2_X1  g196(.A1(new_n612), .A2(new_n619), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n486), .A2(G123), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT83), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n491), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n476), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2096), .ZN(new_n633));
  INV_X1    g208(.A(new_n469), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(new_n478), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT13), .B(G2100), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n632), .A2(new_n633), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT84), .Z(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT85), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n660), .A2(new_n661), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2096), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n665), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n676), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  AOI211_X1 g255(.A(new_n678), .B(new_n680), .C1(new_n673), .C2(new_n677), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT86), .ZN(new_n682));
  XOR2_X1   g257(.A(G1981), .B(G1986), .Z(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n682), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1971), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n689), .A2(G6), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G305), .B2(G16), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT32), .B(G1981), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G288), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(new_n689), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n689), .B2(G23), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT33), .B(G1976), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n694), .A2(new_n696), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n701), .A2(new_n703), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n698), .A2(new_n704), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT90), .B(KEYINPUT34), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n709), .ZN(new_n711));
  MUX2_X1   g286(.A(G24), .B(G290), .S(G16), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT89), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1986), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n715), .A2(G25), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n491), .A2(G131), .ZN(new_n717));
  NOR2_X1   g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT87), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(new_n476), .B2(G107), .ZN(new_n720));
  INV_X1    g295(.A(G119), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n717), .B1(new_n719), .B2(new_n720), .C1(new_n485), .C2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(G29), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT88), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n723), .A2(new_n725), .ZN(new_n727));
  NOR3_X1   g302(.A1(new_n726), .A2(new_n727), .A3(KEYINPUT91), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n710), .A2(new_n711), .A3(new_n714), .A4(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n689), .A2(G4), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n612), .B2(new_n689), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT92), .ZN(new_n734));
  INV_X1    g309(.A(G1348), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT30), .B(G28), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(new_n715), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT31), .B(G11), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n738), .B(new_n739), .C1(new_n631), .C2(new_n715), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT96), .ZN(new_n741));
  INV_X1    g316(.A(G2078), .ZN(new_n742));
  NAND2_X1  g317(.A1(G164), .A2(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G27), .B2(G29), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n736), .B(new_n741), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n729), .A2(new_n730), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n689), .A2(G5), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G171), .B2(new_n689), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1961), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n689), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n689), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n715), .A2(G33), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n491), .A2(G139), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT95), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT25), .Z(new_n758));
  AOI22_X1  g333(.A1(new_n634), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n476), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n754), .B1(new_n761), .B2(new_n715), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n753), .B1(new_n762), .B2(G2072), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT24), .ZN(new_n764));
  INV_X1    g339(.A(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n764), .B2(new_n765), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G160), .B2(new_n715), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n749), .B(new_n763), .C1(G2084), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n689), .A2(G19), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n565), .B2(new_n689), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1341), .Z(new_n772));
  NOR2_X1   g347(.A1(new_n768), .A2(G2084), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT97), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n715), .A2(G26), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT94), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT28), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n486), .A2(G128), .ZN(new_n778));
  NOR2_X1   g353(.A1(G104), .A2(G2105), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT93), .Z(new_n780));
  INV_X1    g355(.A(G116), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n473), .B1(new_n781), .B2(G2105), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n780), .A2(new_n782), .B1(new_n491), .B2(G140), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(G29), .ZN(new_n785));
  INV_X1    g360(.A(G2067), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n774), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n689), .A2(G20), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT23), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n616), .B2(new_n689), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G1956), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n791), .A2(G1956), .ZN(new_n793));
  AOI211_X1 g368(.A(new_n792), .B(new_n793), .C1(G2072), .C2(new_n762), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n769), .A2(new_n772), .A3(new_n788), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n715), .A2(G35), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G162), .B2(new_n715), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT29), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT98), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(G2090), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(G2090), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n715), .A2(G32), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n491), .A2(G141), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n478), .A2(G105), .ZN(new_n805));
  NAND3_X1  g380(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT26), .Z(new_n807));
  NAND3_X1  g382(.A1(new_n804), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n486), .B2(G129), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n803), .B1(new_n809), .B2(new_n715), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT27), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1996), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n742), .B2(new_n744), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n795), .A2(new_n802), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n731), .A2(new_n745), .A3(new_n746), .A4(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  XOR2_X1   g391(.A(KEYINPUT100), .B(G93), .Z(new_n817));
  AOI22_X1  g392(.A1(new_n579), .A2(new_n817), .B1(G55), .B2(new_n528), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n532), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n536), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n818), .B1(new_n820), .B2(KEYINPUT99), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n820), .A2(KEYINPUT99), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n564), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n562), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n612), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n831));
  AOI21_X1  g406(.A(G860), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n831), .B2(new_n830), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT101), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n824), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(new_n631), .B(new_n481), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n493), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n784), .B(new_n523), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n761), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n809), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n491), .A2(G142), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n476), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n486), .B2(G130), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(new_n637), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n722), .B(KEYINPUT102), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n849), .B(new_n850), .Z(new_n851));
  AND2_X1   g426(.A1(new_n851), .A2(KEYINPUT103), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n843), .A2(new_n852), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n840), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n851), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n843), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n843), .A2(new_n856), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n839), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n855), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(G395));
  NOR2_X1   g438(.A1(new_n823), .A2(G868), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n827), .B(new_n622), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n616), .A2(new_n612), .ZN(new_n867));
  NAND2_X1  g442(.A1(G299), .A2(new_n611), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT105), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT106), .B1(new_n869), .B2(KEYINPUT41), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(KEYINPUT41), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(new_n873), .A3(new_n868), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n871), .B1(new_n875), .B2(KEYINPUT106), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(new_n865), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n878));
  INV_X1    g453(.A(new_n869), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n865), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n870), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(G290), .B(G303), .Z(new_n882));
  XNOR2_X1  g457(.A(G288), .B(G305), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT42), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n870), .A2(new_n877), .A3(new_n880), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n864), .B1(new_n889), .B2(G868), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT107), .ZN(G295));
  NAND2_X1  g466(.A1(new_n889), .A2(G868), .ZN(new_n892));
  INV_X1    g467(.A(new_n864), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(G331));
  XNOR2_X1  g469(.A(G286), .B(G171), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n827), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n827), .A2(new_n896), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT108), .B1(new_n827), .B2(new_n896), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n899), .A2(new_n879), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n900), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(new_n897), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n876), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(new_n884), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n905), .B2(new_n884), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n907), .B2(KEYINPUT109), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n909));
  INV_X1    g484(.A(new_n884), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n904), .A2(new_n876), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(new_n902), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n909), .B1(new_n912), .B2(G37), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT43), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n860), .B1(new_n905), .B2(new_n884), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n875), .ZN(new_n918));
  OR3_X1    g493(.A1(new_n903), .A2(new_n869), .A3(new_n897), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n910), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n915), .A2(new_n916), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT44), .B1(new_n914), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n916), .B1(new_n908), .B2(new_n913), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n915), .A2(KEYINPUT43), .A3(new_n920), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(G397));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT45), .B1(new_n523), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g504(.A(KEYINPUT110), .B(G40), .Z(new_n930));
  NOR2_X1   g505(.A1(new_n481), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n784), .B(new_n786), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(new_n809), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n932), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT46), .B1(new_n932), .B2(G1996), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n937), .B(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n932), .ZN(new_n940));
  INV_X1    g515(.A(G1996), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(new_n809), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n942), .A2(KEYINPUT111), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(KEYINPUT111), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n933), .B1(new_n941), .B2(new_n809), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n943), .A2(new_n944), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n724), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n778), .A2(new_n786), .A3(new_n783), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n932), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n722), .A2(new_n947), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n940), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n946), .A2(new_n953), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n932), .A2(G1986), .A3(G290), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT48), .Z(new_n956));
  AOI211_X1 g531(.A(new_n939), .B(new_n951), .C1(new_n954), .C2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G8), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n523), .A2(new_n928), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT4), .B1(new_n515), .B2(KEYINPUT72), .ZN(new_n962));
  INV_X1    g537(.A(new_n506), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT73), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n511), .A2(new_n518), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n965), .A3(new_n507), .ZN(new_n966));
  AOI21_X1  g541(.A(G1384), .B1(new_n966), .B2(new_n499), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n961), .A2(new_n931), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n752), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n959), .A2(KEYINPUT50), .ZN(new_n971));
  INV_X1    g546(.A(new_n931), .ZN(new_n972));
  NOR2_X1   g547(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n523), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G2084), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n958), .B1(new_n970), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g552(.A(KEYINPUT113), .B(G8), .Z(new_n978));
  NOR2_X1   g553(.A1(G168), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT51), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AOI211_X1 g555(.A(G168), .B(new_n978), .C1(new_n970), .C2(new_n976), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n978), .B1(new_n970), .B2(new_n976), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n979), .A2(KEYINPUT51), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n980), .A2(new_n981), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI221_X1 g562(.A(KEYINPUT62), .B1(new_n982), .B2(new_n984), .C1(new_n980), .C2(new_n981), .ZN(new_n988));
  NAND2_X1  g563(.A1(G303), .A2(G8), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT55), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n523), .A2(new_n973), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n991), .B(new_n931), .C1(new_n967), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G2090), .ZN(new_n995));
  INV_X1    g570(.A(G1971), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n994), .A2(new_n995), .B1(new_n969), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n990), .B1(new_n997), .B2(new_n978), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n978), .B1(new_n967), .B2(new_n931), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n699), .A2(G1976), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT52), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n523), .A2(new_n931), .A3(new_n928), .ZN(new_n1003));
  INV_X1    g578(.A(new_n978), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(G288), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1003), .A2(new_n1000), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1981), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n592), .A2(new_n597), .A3(new_n1008), .A4(new_n595), .ZN(new_n1009));
  OR2_X1    g584(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n528), .A2(G48), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n532), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n1012), .B2(new_n536), .ZN(new_n1013));
  OAI21_X1  g588(.A(G1981), .B1(new_n1013), .B2(new_n596), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1009), .A2(new_n1010), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1009), .A2(KEYINPUT114), .A3(KEYINPUT49), .A4(new_n1014), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n1003), .A3(new_n1004), .A4(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1002), .A2(KEYINPUT116), .A3(new_n1007), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1007), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n999), .B2(new_n1000), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n961), .A2(new_n931), .A3(new_n968), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1027), .A2(G1971), .B1(G2090), .B2(new_n993), .ZN(new_n1028));
  INV_X1    g603(.A(new_n990), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(G8), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n998), .A2(new_n1026), .A3(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n961), .A2(new_n968), .A3(new_n742), .A4(new_n931), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n1033));
  INV_X1    g608(.A(G1961), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1032), .A2(new_n1033), .B1(new_n1034), .B2(new_n993), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1033), .A2(G2078), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1027), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G171), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1031), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n987), .A2(new_n988), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1019), .A2(new_n1005), .A3(new_n699), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1009), .B(KEYINPUT115), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n999), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1002), .A2(new_n1007), .A3(new_n1019), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n1030), .B2(new_n1045), .ZN(new_n1046));
  AOI211_X1 g621(.A(G286), .B(new_n978), .C1(new_n970), .C2(new_n976), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n998), .A2(new_n1026), .A3(new_n1030), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT63), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n990), .B1(new_n997), .B2(new_n958), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1052), .A3(new_n1030), .A4(new_n1047), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1046), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1041), .A2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT56), .B(G2072), .Z(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT118), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n961), .A2(new_n968), .A3(new_n931), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n1059), .B(G1956), .C1(new_n971), .C2(new_n974), .ZN(new_n1060));
  INV_X1    g635(.A(G1956), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT117), .B1(new_n993), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1058), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  XOR2_X1   g638(.A(G299), .B(KEYINPUT57), .Z(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1003), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n993), .A2(new_n735), .B1(new_n1067), .B2(new_n786), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n611), .B2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1064), .B(new_n1058), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n993), .A2(new_n735), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1067), .A2(new_n786), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(KEYINPUT60), .A3(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1074), .A2(KEYINPUT121), .A3(new_n611), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n611), .B1(new_n1074), .B2(KEYINPUT121), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n1075), .A2(new_n1076), .B1(KEYINPUT121), .B2(new_n1074), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1068), .A2(KEYINPUT60), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1066), .A2(KEYINPUT61), .A3(new_n1070), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT120), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n969), .A2(G1996), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT58), .B(G1341), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1067), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n565), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT59), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1066), .A2(new_n1087), .A3(KEYINPUT61), .A4(new_n1070), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1079), .A2(new_n1081), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT61), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT119), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n1093));
  AOI211_X1 g668(.A(new_n1093), .B(KEYINPUT61), .C1(new_n1066), .C2(new_n1070), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1071), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n480), .ZN(new_n1097));
  INV_X1    g672(.A(G101), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n474), .B2(new_n477), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT122), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n479), .A2(new_n1101), .A3(new_n480), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1100), .A2(new_n1102), .A3(G40), .A4(new_n472), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT123), .Z(new_n1104));
  NAND3_X1  g679(.A1(new_n961), .A2(new_n1104), .A3(KEYINPUT124), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1103), .B(KEYINPUT123), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n929), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1105), .A2(new_n1108), .A3(new_n968), .A4(new_n1036), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1112));
  OAI211_X1 g687(.A(G301), .B(new_n1035), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1038), .B2(G171), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1109), .B(new_n1110), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1118), .A2(new_n1114), .A3(G301), .A4(new_n1035), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1035), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G171), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1038), .A2(G171), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(new_n1117), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1031), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n985), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1120), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1055), .B1(new_n1096), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(G290), .B(G1986), .Z(new_n1129));
  OAI21_X1  g704(.A(new_n954), .B1(new_n932), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT112), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1130), .B(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n957), .B1(new_n1128), .B2(new_n1132), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g708(.A1(G229), .A2(new_n464), .A3(G227), .ZN(new_n1135));
  AND2_X1   g709(.A1(new_n1135), .A2(new_n657), .ZN(new_n1136));
  OAI211_X1 g710(.A(new_n1136), .B(new_n861), .C1(new_n924), .C2(new_n925), .ZN(G225));
  INV_X1    g711(.A(G225), .ZN(G308));
endmodule


