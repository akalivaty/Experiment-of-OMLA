//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n464), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n470), .A2(G2105), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n464), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n476), .B1(new_n466), .B2(G2104), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n474), .A2(G137), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n477), .A2(new_n473), .A3(G2105), .A4(new_n467), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  OAI221_X1 g061(.A(new_n482), .B1(new_n483), .B2(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n475), .B2(G114), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(new_n484), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n477), .A2(new_n473), .A3(new_n502), .A4(new_n467), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT3), .B(G2104), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n501), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(KEYINPUT4), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n500), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT70), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(G88), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n514), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(KEYINPUT71), .A3(new_n515), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n510), .A2(new_n512), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n520), .A2(new_n523), .B1(G651), .B2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n514), .A2(G51), .A3(G543), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n513), .A2(G89), .A3(new_n514), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n513), .A2(new_n514), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n539), .A2(new_n540), .B1(new_n517), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n538), .A2(new_n542), .ZN(G171));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n539), .A2(new_n544), .B1(new_n517), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n513), .A2(G56), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n537), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n510), .B2(new_n512), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n558));
  AND2_X1   g133(.A1(G78), .A2(G543), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(G651), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n517), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n514), .A2(new_n565), .A3(G53), .A4(G543), .ZN(new_n566));
  INV_X1    g141(.A(new_n539), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n564), .A2(new_n566), .B1(new_n567), .B2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n562), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  NAND2_X1  g146(.A1(new_n527), .A2(G651), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n518), .A2(new_n519), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT71), .B1(new_n522), .B2(new_n515), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(G303));
  OR2_X1    g150(.A1(new_n513), .A2(G74), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G49), .B2(new_n521), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT73), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n567), .B2(G87), .ZN(new_n579));
  INV_X1    g154(.A(G87), .ZN(new_n580));
  NOR3_X1   g155(.A1(new_n539), .A2(KEYINPUT73), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n577), .B1(new_n579), .B2(new_n581), .ZN(G288));
  AOI22_X1  g157(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n537), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n539), .A2(new_n585), .B1(new_n517), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n567), .A2(G85), .B1(new_n521), .B2(G47), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n537), .B2(new_n591), .ZN(G290));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT10), .B1(new_n539), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n510), .B2(new_n512), .ZN(new_n596));
  AND2_X1   g171(.A1(G79), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n521), .A2(G54), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n513), .A2(new_n600), .A3(G92), .A4(new_n514), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n594), .A2(new_n598), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n603), .B2(G171), .ZN(G321));
  XNOR2_X1  g180(.A(G321), .B(KEYINPUT74), .ZN(G284));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n562), .A2(new_n568), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(new_n602), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  NOR2_X1   g188(.A1(new_n602), .A2(G559), .ZN(new_n614));
  OR3_X1    g189(.A1(new_n614), .A2(KEYINPUT75), .A3(new_n603), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT75), .B1(new_n614), .B2(new_n603), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n615), .B(new_n616), .C1(G868), .C2(new_n550), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n504), .A2(new_n471), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  OR2_X1    g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n624));
  INV_X1    g199(.A(G123), .ZN(new_n625));
  INV_X1    g200(.A(G135), .ZN(new_n626));
  OAI221_X1 g201(.A(new_n624), .B1(new_n625), .B2(new_n484), .C1(new_n485), .C2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT76), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2430), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(G14), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n642), .B2(new_n643), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  XNOR2_X1  g223(.A(G2096), .B(G2100), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(KEYINPUT78), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(KEYINPUT78), .B2(new_n652), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n652), .B(KEYINPUT17), .Z(new_n657));
  INV_X1    g232(.A(new_n651), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n654), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT79), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT80), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n655), .A2(new_n652), .A3(new_n651), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT77), .B(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n656), .A2(new_n651), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n664), .B1(new_n657), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n660), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n661), .B1(new_n660), .B2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n650), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n671), .A2(new_n667), .A3(new_n649), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(KEYINPUT82), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT81), .B(KEYINPUT19), .Z(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(KEYINPUT82), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n679), .A2(new_n680), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n681), .A2(new_n689), .ZN(new_n690));
  MUX2_X1   g265(.A(new_n690), .B(new_n689), .S(new_n685), .Z(new_n691));
  AOI21_X1  g266(.A(new_n678), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n688), .A2(new_n691), .A3(new_n678), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n677), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n694), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n696), .A2(new_n676), .A3(new_n692), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n675), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n676), .B1(new_n696), .B2(new_n692), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n693), .A2(new_n677), .A3(new_n694), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n699), .A2(new_n700), .A3(new_n674), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n704), .A2(G33), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n504), .A2(G127), .ZN(new_n706));
  NAND2_X1  g281(.A1(G115), .A2(G2104), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n475), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n709), .B2(new_n708), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT25), .ZN(new_n713));
  INV_X1    g288(.A(new_n485), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G139), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n705), .B1(new_n716), .B2(G29), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G2072), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n704), .A2(G27), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G164), .B2(new_n704), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT98), .B(G2078), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n720), .B(new_n721), .Z(new_n722));
  NOR2_X1   g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT31), .B(G11), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT95), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT30), .B(G28), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n704), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n728), .A2(G5), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G301), .B2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n727), .B1(new_n704), .B2(new_n627), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n728), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n728), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT94), .B(G1966), .Z(new_n735));
  XOR2_X1   g310(.A(new_n734), .B(new_n735), .Z(new_n736));
  NOR2_X1   g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT96), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n740), .B2(KEYINPUT24), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(KEYINPUT24), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n479), .B2(new_n704), .ZN(new_n743));
  INV_X1    g318(.A(G2084), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT91), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(KEYINPUT91), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n704), .A2(G32), .ZN(new_n748));
  INV_X1    g323(.A(G141), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n485), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n471), .A2(G105), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G129), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n484), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT92), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n748), .B1(new_n760), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT27), .B(G1996), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n746), .A2(new_n747), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(KEYINPUT96), .B1(new_n732), .B2(new_n736), .ZN(new_n764));
  AND4_X1   g339(.A1(new_n723), .A2(new_n739), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n489), .A2(G29), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n704), .A2(G35), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT29), .ZN(new_n770));
  INV_X1    g345(.A(G2090), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n766), .A2(new_n772), .A3(new_n768), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n770), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n730), .A2(new_n731), .B1(new_n743), .B2(new_n744), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n761), .B2(new_n762), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT97), .Z(new_n777));
  AND3_X1   g352(.A1(new_n765), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT101), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n728), .A2(G4), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n611), .B2(new_n728), .ZN(new_n781));
  INV_X1    g356(.A(G1348), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G19), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n550), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT87), .B(G1341), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n704), .A2(G26), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(G104), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n792));
  INV_X1    g367(.A(G128), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n484), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n714), .B2(G140), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n790), .B1(new_n795), .B2(new_n704), .ZN(new_n796));
  INV_X1    g371(.A(G2067), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n783), .A2(new_n787), .A3(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT89), .Z(new_n800));
  AOI21_X1  g375(.A(new_n771), .B1(new_n770), .B2(new_n773), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n728), .A2(G20), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT99), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT23), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G299), .B2(G16), .ZN(new_n805));
  INV_X1    g380(.A(G1956), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  OR3_X1    g382(.A1(new_n801), .A2(KEYINPUT100), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT100), .B1(new_n801), .B2(new_n807), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n778), .A2(new_n779), .A3(new_n800), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n765), .A2(new_n800), .A3(new_n774), .A4(new_n777), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n808), .A2(new_n809), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT101), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n588), .A2(G16), .ZN(new_n816));
  OR2_X1    g391(.A1(G6), .A2(G16), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT32), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT32), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n816), .A2(new_n820), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G1981), .ZN(new_n823));
  INV_X1    g398(.A(G1981), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n819), .A2(new_n824), .A3(new_n821), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  MUX2_X1   g401(.A(G23), .B(G288), .S(G16), .Z(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT33), .B(G1976), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n728), .A2(G22), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G166), .B2(new_n728), .ZN(new_n831));
  INV_X1    g406(.A(G1971), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n826), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n714), .A2(G131), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(G95), .A2(G2105), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n838), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT83), .ZN(new_n840));
  INV_X1    g415(.A(new_n484), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G119), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G29), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G25), .B2(G29), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT35), .B(G1991), .Z(new_n847));
  AND2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n728), .A2(G24), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT84), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G290), .B2(G16), .ZN(new_n852));
  INV_X1    g427(.A(G1986), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  OR3_X1    g429(.A1(new_n848), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n835), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n834), .A2(KEYINPUT85), .A3(KEYINPUT34), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT85), .B1(new_n834), .B2(KEYINPUT34), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT86), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT86), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n856), .B(new_n861), .C1(new_n858), .C2(new_n857), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(KEYINPUT36), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT36), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n859), .A2(KEYINPUT86), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n815), .A2(new_n863), .A3(new_n865), .ZN(G311));
  NAND3_X1  g441(.A1(new_n815), .A2(new_n863), .A3(new_n865), .ZN(G150));
  NOR2_X1   g442(.A1(new_n602), .A2(new_n612), .ZN(new_n868));
  XNOR2_X1  g443(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n871));
  NAND2_X1  g446(.A1(G80), .A2(G543), .ZN(new_n872));
  INV_X1    g447(.A(G67), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n871), .B(new_n872), .C1(new_n525), .C2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n873), .B1(new_n510), .B2(new_n512), .ZN(new_n875));
  INV_X1    g450(.A(new_n872), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT103), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(G651), .A3(new_n877), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n567), .A2(G93), .B1(new_n521), .B2(G55), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n546), .A2(new_n549), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n550), .A2(new_n878), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n870), .B(new_n884), .Z(new_n885));
  AND2_X1   g460(.A1(new_n885), .A2(KEYINPUT39), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(KEYINPUT39), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n886), .A2(new_n887), .A3(G860), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n880), .A2(G860), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT37), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n888), .A2(new_n890), .ZN(G145));
  NOR2_X1   g466(.A1(new_n760), .A2(new_n716), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n760), .A2(new_n716), .ZN(new_n894));
  INV_X1    g469(.A(new_n620), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n837), .B2(new_n843), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n836), .A2(new_n620), .A3(new_n840), .A4(new_n842), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n894), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  INV_X1    g475(.A(new_n894), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n901), .B2(new_n892), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n504), .A2(new_n505), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n841), .A2(G126), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT104), .A4(new_n498), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n500), .B2(new_n506), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n795), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n908), .A2(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n795), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g491(.A1(G106), .A2(G2105), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n917), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n918));
  INV_X1    g493(.A(G130), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n484), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n714), .B2(G142), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n921), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n913), .A2(new_n923), .A3(new_n915), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n903), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G160), .B(new_n627), .ZN(new_n927));
  XNOR2_X1  g502(.A(G162), .B(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n899), .A2(new_n902), .A3(new_n922), .A4(new_n924), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G37), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n926), .A2(new_n929), .ZN(new_n933));
  INV_X1    g508(.A(new_n928), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n933), .A2(KEYINPUT105), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT105), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(KEYINPUT106), .B(new_n932), .C1(new_n935), .C2(new_n936), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n939), .A2(KEYINPUT40), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT40), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(G395));
  NOR2_X1   g518(.A1(G288), .A2(G290), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n946));
  NAND2_X1  g521(.A1(G288), .A2(G290), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT109), .B1(new_n949), .B2(new_n944), .ZN(new_n950));
  XNOR2_X1  g525(.A(G166), .B(new_n588), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(G166), .B(G305), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n953), .B(KEYINPUT109), .C1(new_n949), .C2(new_n944), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT42), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n562), .A2(new_n568), .A3(KEYINPUT107), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n611), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT107), .B1(new_n562), .B2(new_n568), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n608), .A2(KEYINPUT107), .A3(new_n611), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT41), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n958), .A2(new_n959), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n965));
  NAND2_X1  g540(.A1(G299), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(new_n611), .A3(new_n957), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT41), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n962), .A2(new_n963), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n884), .B(new_n614), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n964), .A2(new_n967), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(KEYINPUT108), .A3(KEYINPUT41), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n971), .B2(new_n972), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n975), .A2(KEYINPUT110), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(KEYINPUT110), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n956), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n977), .A2(new_n956), .ZN(new_n979));
  OAI21_X1  g554(.A(G868), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n880), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(G868), .B2(new_n981), .ZN(G295));
  OAI21_X1  g557(.A(new_n980), .B1(G868), .B2(new_n981), .ZN(G331));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n984));
  AOI21_X1  g559(.A(G301), .B1(G168), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(G286), .A2(KEYINPUT111), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n882), .A2(new_n987), .A3(new_n883), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n987), .B1(new_n882), .B2(new_n883), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n987), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n884), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n882), .A2(new_n987), .A3(new_n883), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n993), .A3(new_n985), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n970), .A2(new_n995), .A3(new_n973), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n990), .A2(new_n994), .A3(new_n964), .A4(new_n967), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n955), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n931), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n955), .B1(new_n996), .B2(new_n997), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT43), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT112), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1003), .B(KEYINPUT43), .C1(new_n999), .C2(new_n1000), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n962), .A2(new_n1005), .A3(new_n969), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n964), .A2(new_n967), .A3(KEYINPUT113), .A4(new_n968), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n995), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT114), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1006), .A2(new_n995), .A3(new_n1010), .A4(new_n1007), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n997), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n955), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n1015));
  INV_X1    g590(.A(new_n999), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1002), .A2(new_n1004), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1014), .A2(KEYINPUT43), .A3(new_n1016), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n999), .A2(new_n1000), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(KEYINPUT43), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT44), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(new_n1024), .ZN(G397));
  OR2_X1    g600(.A1(G288), .A2(G1976), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n588), .A2(new_n824), .ZN(new_n1027));
  OAI21_X1  g602(.A(G1981), .B1(new_n584), .B2(new_n587), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(KEYINPUT120), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n1031));
  NAND3_X1  g606(.A1(G305), .A2(new_n1031), .A3(G1981), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1029), .A2(new_n1032), .A3(KEYINPUT121), .A4(new_n1030), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n500), .B2(new_n506), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n470), .A2(G2105), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n471), .A2(G101), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1041), .A2(new_n478), .A3(G40), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n472), .A2(KEYINPUT115), .A3(G40), .A4(new_n478), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1040), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G8), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(KEYINPUT49), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1026), .B1(new_n1037), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1027), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n577), .B(G1976), .C1(new_n579), .C2(new_n581), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT52), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1976), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1058), .A2(new_n1047), .A3(G8), .A4(new_n1054), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n1037), .B2(new_n1050), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT45), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1039), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1063), .A2(G1384), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n908), .A2(new_n910), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT117), .A4(new_n1066), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1039), .A2(KEYINPUT50), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n1038), .C1(new_n500), .C2(new_n506), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1072), .A2(new_n1045), .A3(new_n1046), .A4(new_n1074), .ZN(new_n1075));
  OAI22_X1  g650(.A1(new_n1071), .A2(G1971), .B1(G2090), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n1077));
  NAND4_X1  g652(.A1(G303), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n1079));
  INV_X1    g654(.A(G8), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1079), .B1(G166), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n520), .A2(new_n523), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1080), .B1(new_n1083), .B2(new_n572), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT118), .B1(new_n1084), .B2(KEYINPUT55), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1077), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(KEYINPUT119), .A3(new_n1081), .A4(new_n1078), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1076), .A2(new_n1086), .A3(G8), .A4(new_n1090), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1053), .A2(new_n1048), .B1(new_n1062), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT122), .B1(new_n564), .B2(new_n566), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(KEYINPUT57), .ZN(new_n1094));
  XNOR2_X1  g669(.A(G299), .B(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1065), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1075), .A2(new_n806), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1095), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1099), .A2(new_n1095), .A3(new_n1100), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1075), .A2(new_n782), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(new_n797), .A3(new_n1040), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1103), .A2(new_n1105), .A3(KEYINPUT123), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n611), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1102), .B1(new_n1110), .B2(KEYINPUT124), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1108), .A2(new_n1112), .A3(new_n611), .A4(new_n1109), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1101), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1103), .A2(new_n1105), .A3(KEYINPUT123), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT123), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT60), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1108), .A2(new_n1118), .A3(new_n1109), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1119), .A3(new_n611), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1047), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1996), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n1071), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT59), .B1(new_n1125), .B2(new_n881), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1096), .A2(new_n1124), .A3(new_n1097), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1122), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n550), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1099), .A2(new_n1095), .A3(new_n1100), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1099), .A2(KEYINPUT61), .A3(new_n1095), .A4(new_n1100), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(KEYINPUT60), .B(new_n602), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1120), .A2(new_n1131), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1114), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1075), .A2(G2090), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n832), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1140), .B1(new_n1143), .B2(new_n1080), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(new_n1061), .A3(new_n1091), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1075), .A2(new_n731), .ZN(new_n1146));
  INV_X1    g721(.A(G2078), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1096), .A2(new_n1147), .A3(new_n1097), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(G171), .B(KEYINPUT54), .Z(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT45), .B1(new_n911), .B2(new_n1038), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1149), .A2(G2078), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1043), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1151), .B1(new_n1156), .B2(new_n1096), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1150), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1066), .B1(new_n500), .B2(new_n506), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1064), .A2(new_n1045), .A3(new_n1046), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1160), .A2(new_n1154), .ZN(new_n1161));
  AOI211_X1 g736(.A(new_n1161), .B(new_n1146), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1151), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1158), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1104), .A2(new_n744), .A3(new_n1074), .A4(new_n1072), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1160), .A2(new_n735), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(new_n1166), .A3(G168), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT51), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1167), .A2(new_n1168), .A3(G8), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1160), .A2(new_n735), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1075), .A2(G2084), .ZN(new_n1171));
  OAI21_X1  g746(.A(G286), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1172), .A2(G8), .A3(new_n1167), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1169), .B1(KEYINPUT51), .B2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1145), .A2(new_n1164), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1092), .B1(new_n1139), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1167), .A2(G8), .ZN(new_n1178));
  AOI21_X1  g753(.A(G168), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT51), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1167), .A2(new_n1168), .A3(G8), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1161), .ZN(new_n1184));
  AOI21_X1  g759(.A(G301), .B1(new_n1150), .B2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1185), .A2(new_n1144), .A3(new_n1091), .A4(new_n1061), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1177), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1144), .A2(new_n1061), .A3(new_n1091), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1188), .A2(KEYINPUT125), .A3(new_n1189), .A4(new_n1185), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n1174), .A2(new_n1181), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1187), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI211_X1 g767(.A(new_n1080), .B(G286), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1144), .A2(new_n1061), .A3(new_n1091), .A4(new_n1193), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT63), .Z(new_n1195));
  NAND3_X1  g770(.A1(new_n1176), .A2(new_n1192), .A3(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n844), .B(new_n847), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT116), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n912), .A2(G2067), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n795), .A2(new_n797), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(G1996), .B1(new_n755), .B2(new_n759), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n760), .A2(new_n1124), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1198), .A2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g780(.A(G290), .B(new_n853), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1152), .A2(new_n1104), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1196), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1209), .A2(new_n1124), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1212), .B(KEYINPUT46), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1201), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1209), .B1(new_n760), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  XOR2_X1   g791(.A(new_n1216), .B(KEYINPUT47), .Z(new_n1217));
  NOR3_X1   g792(.A1(new_n1208), .A2(G1986), .A3(G290), .ZN(new_n1218));
  OAI22_X1  g793(.A1(new_n1205), .A2(new_n1208), .B1(KEYINPUT48), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1219), .B1(KEYINPUT48), .B2(new_n1218), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n844), .A2(new_n847), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1200), .B1(new_n1204), .B2(new_n1221), .ZN(new_n1222));
  AND2_X1   g797(.A1(new_n1222), .A2(new_n1209), .ZN(new_n1223));
  NOR3_X1   g798(.A1(new_n1217), .A2(new_n1220), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1211), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n1227));
  NAND2_X1  g801(.A1(new_n647), .A2(G319), .ZN(new_n1228));
  OAI21_X1  g802(.A(new_n1227), .B1(G227), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g803(.A(new_n462), .B1(new_n644), .B2(new_n646), .ZN(new_n1230));
  NAND4_X1  g804(.A1(new_n1230), .A2(KEYINPUT126), .A3(new_n672), .A4(new_n670), .ZN(new_n1231));
  NAND3_X1  g805(.A1(new_n702), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g808(.A1(new_n702), .A2(new_n1229), .A3(KEYINPUT127), .A4(new_n1231), .ZN(new_n1235));
  AOI22_X1  g809(.A1(new_n939), .A2(new_n940), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AND2_X1   g810(.A1(new_n1236), .A2(new_n1018), .ZN(G308));
  NAND2_X1  g811(.A1(new_n1236), .A2(new_n1018), .ZN(G225));
endmodule


