//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1301, new_n1302, new_n1303,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n207), .B1(new_n202), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n201), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n206), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT1), .Z(new_n218));
  INV_X1    g0018(.A(KEYINPUT64), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(new_n206), .B2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G13), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n221), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n203), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n218), .A2(new_n225), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n238), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G58), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND2_X1  g0050(.A1(G33), .A2(G97), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT19), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n229), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G97), .A2(G107), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n209), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n258), .A2(new_n260), .A3(new_n229), .A4(G68), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n229), .A2(G33), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n252), .B1(new_n262), .B2(new_n214), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n256), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n265), .A2(KEYINPUT69), .A3(new_n228), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT69), .B1(new_n265), .B2(new_n228), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT15), .B(G87), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n221), .A2(new_n229), .A3(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n271), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n274), .B(new_n276), .C1(new_n266), .C2(new_n267), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT87), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(G87), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT87), .B1(new_n277), .B2(new_n209), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n273), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  OAI211_X1 g0083(.A(G1), .B(G13), .C1(new_n257), .C2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n258), .A2(new_n260), .A3(G244), .A4(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT85), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n288), .A2(KEYINPUT85), .A3(G244), .A4(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OR2_X1    g0090(.A1(KEYINPUT86), .A2(G116), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT86), .A2(G116), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n257), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n258), .A2(new_n260), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n293), .B1(new_n295), .B2(G238), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n284), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n284), .A2(G274), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G1), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(new_n210), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n298), .A2(new_n300), .B1(new_n284), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(G200), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n258), .A2(new_n260), .A3(G238), .A4(new_n294), .ZN(new_n305));
  AND2_X1   g0105(.A1(KEYINPUT86), .A2(G116), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT86), .A2(G116), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n305), .B1(new_n308), .B2(new_n257), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n287), .B2(new_n289), .ZN(new_n310));
  OAI211_X1 g0110(.A(G190), .B(new_n302), .C1(new_n310), .C2(new_n284), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n282), .A2(new_n304), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n313), .B(new_n302), .C1(new_n310), .C2(new_n284), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n269), .B(new_n272), .C1(new_n277), .C2(new_n270), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n297), .A2(new_n303), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n314), .B(new_n315), .C1(new_n316), .C2(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT82), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n295), .A2(new_n319), .A3(KEYINPUT4), .A4(G244), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n258), .A2(new_n260), .A3(G250), .A4(G1698), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G283), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n258), .A2(new_n260), .A3(G244), .A4(new_n294), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT4), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT82), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n325), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n320), .A2(new_n323), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT5), .B(G41), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n298), .A2(new_n300), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n300), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n284), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n215), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n330), .A2(G179), .A3(new_n332), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n284), .A2(G274), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  AOI211_X1 g0139(.A(new_n339), .B(new_n335), .C1(new_n328), .C2(new_n329), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G107), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT7), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n288), .B2(G20), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n258), .A2(new_n260), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G20), .A2(G33), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G77), .ZN(new_n350));
  NAND2_X1  g0150(.A1(KEYINPUT6), .A2(G97), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(G107), .ZN(new_n352));
  XNOR2_X1  g0152(.A(G97), .B(G107), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT6), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n350), .B1(new_n355), .B2(new_n229), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n268), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n277), .A2(new_n214), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n274), .A2(G97), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n357), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT84), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT84), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n357), .A2(new_n359), .A3(new_n364), .A4(new_n361), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT83), .ZN(new_n367));
  INV_X1    g0167(.A(new_n268), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT7), .B1(new_n346), .B2(new_n229), .ZN(new_n369));
  AOI211_X1 g0169(.A(new_n344), .B(G20), .C1(new_n258), .C2(new_n260), .ZN(new_n370));
  OAI21_X1  g0170(.A(G107), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(G97), .A2(G107), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n354), .B1(new_n372), .B2(new_n254), .ZN(new_n373));
  INV_X1    g0173(.A(new_n352), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(G20), .B1(G77), .B2(new_n349), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n368), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n377), .A2(new_n358), .A3(new_n360), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n330), .A2(G190), .A3(new_n332), .A4(new_n336), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G200), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n335), .B1(new_n328), .B2(new_n329), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n332), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n367), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n330), .A2(new_n332), .A3(new_n336), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G200), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n386), .A2(KEYINPUT83), .A3(new_n378), .A4(new_n379), .ZN(new_n387));
  AOI221_X4 g0187(.A(new_n318), .B1(new_n342), .B2(new_n366), .C1(new_n384), .C2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n266), .ZN(new_n389));
  INV_X1    g0189(.A(new_n267), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n271), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n229), .A2(G1), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(G50), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n349), .A2(G150), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n398), .A2(KEYINPUT70), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(KEYINPUT70), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT8), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G58), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n262), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n394), .B1(G50), .B2(new_n274), .C1(new_n405), .C2(new_n368), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT9), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT77), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n405), .A2(new_n368), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n274), .A2(G50), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT77), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT9), .A4(new_n394), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n295), .A2(G222), .ZN(new_n415));
  INV_X1    g0215(.A(G77), .ZN(new_n416));
  INV_X1    g0216(.A(G223), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n288), .A2(G1698), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n415), .B1(new_n416), .B2(new_n288), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n329), .ZN(new_n420));
  AOI21_X1  g0220(.A(G1), .B1(new_n283), .B2(new_n299), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n284), .A2(G274), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n284), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT68), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n425), .B(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n423), .B1(new_n427), .B2(G226), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n381), .B1(new_n420), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n420), .A2(new_n428), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n430), .B2(G190), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n414), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n406), .A2(new_n407), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(KEYINPUT76), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT76), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n406), .B2(new_n407), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT10), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n433), .B(KEYINPUT76), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT10), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n414), .A4(new_n431), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n391), .A2(G77), .A3(new_n393), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n271), .A2(new_n416), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT73), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n349), .B(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n398), .A2(new_n402), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT72), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT72), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n398), .A2(new_n402), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n447), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n229), .A2(new_n416), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT74), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(KEYINPUT74), .A3(new_n454), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n457), .B(new_n458), .C1(new_n262), .C2(new_n270), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n445), .B1(new_n459), .B2(new_n268), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n423), .B1(new_n427), .B2(G244), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n418), .A2(new_n208), .B1(new_n343), .B2(new_n288), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n346), .A2(new_n213), .A3(G1698), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n329), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(G169), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT75), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n458), .B1(new_n262), .B2(new_n270), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT74), .B1(new_n452), .B2(new_n454), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n268), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(new_n444), .A3(new_n443), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT75), .ZN(new_n471));
  INV_X1    g0271(.A(new_n465), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n461), .A2(new_n313), .A3(new_n464), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n466), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n461), .A2(new_n464), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G200), .ZN(new_n477));
  INV_X1    g0277(.A(G190), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n460), .B(new_n477), .C1(new_n478), .C2(new_n476), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n288), .A2(G232), .A3(G1698), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n288), .A2(new_n294), .ZN(new_n482));
  INV_X1    g0282(.A(G226), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n481), .B(new_n251), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n329), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n425), .A2(new_n426), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT68), .B1(new_n284), .B2(new_n424), .ZN(new_n487));
  OAI21_X1  g0287(.A(G238), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n422), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT13), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n485), .A2(new_n488), .A3(KEYINPUT13), .A4(new_n422), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(G169), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT14), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n423), .B1(new_n427), .B2(G238), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(new_n485), .B1(KEYINPUT79), .B2(KEYINPUT13), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT79), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(G179), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT14), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n491), .A2(new_n500), .A3(G169), .A4(new_n492), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n494), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n271), .A2(new_n202), .ZN(new_n503));
  XOR2_X1   g0303(.A(new_n503), .B(KEYINPUT12), .Z(new_n504));
  AOI22_X1  g0304(.A1(new_n349), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n416), .B2(new_n262), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT11), .B1(new_n268), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n268), .A2(new_n506), .A3(KEYINPUT11), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n391), .A2(G68), .A3(new_n393), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n491), .A2(G200), .A3(new_n492), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT78), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n491), .A2(KEYINPUT78), .A3(G200), .A4(new_n492), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n489), .B1(new_n497), .B2(new_n490), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n497), .B2(new_n492), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n511), .B1(new_n519), .B2(G190), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n442), .A2(new_n480), .A3(new_n512), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n430), .A2(new_n313), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n523), .B(KEYINPUT71), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n406), .B1(new_n430), .B2(G169), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n422), .B1(new_n425), .B2(new_n213), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n288), .A2(G223), .A3(new_n294), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G87), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(new_n529), .C1(new_n418), .C2(new_n483), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n527), .B1(new_n530), .B2(new_n329), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT81), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n532), .A3(new_n313), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n532), .B1(new_n531), .B2(new_n313), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n534), .A2(new_n535), .B1(G169), .B2(new_n531), .ZN(new_n536));
  OAI21_X1  g0336(.A(G68), .B1(new_n369), .B2(new_n370), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT80), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G58), .A2(G68), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n229), .B1(new_n203), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n349), .A2(G159), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n539), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G58), .A2(G68), .ZN(new_n545));
  OAI21_X1  g0345(.A(G20), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(KEYINPUT80), .A3(new_n541), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n537), .A2(KEYINPUT16), .A3(new_n543), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT16), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n543), .A2(new_n547), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n202), .B1(new_n345), .B2(new_n347), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(new_n552), .A3(new_n268), .ZN(new_n553));
  INV_X1    g0353(.A(new_n403), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n392), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n391), .B1(new_n271), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT18), .B1(new_n536), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n531), .A2(G169), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n531), .A2(new_n313), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT81), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n560), .B1(new_n562), .B2(new_n533), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT18), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n557), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n531), .A2(new_n478), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G200), .B2(new_n531), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n553), .A3(new_n556), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT17), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n526), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n522), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n329), .B1(new_n300), .B2(new_n331), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G270), .ZN(new_n577));
  INV_X1    g0377(.A(G303), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n346), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G257), .A2(G1698), .ZN(new_n580));
  INV_X1    g0380(.A(G264), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(G1698), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n579), .B(new_n329), .C1(new_n346), .C2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n577), .A2(new_n332), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(new_n341), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n322), .B(new_n229), .C1(G33), .C2(new_n214), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n306), .A2(new_n307), .A3(new_n229), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n265), .A2(new_n228), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT88), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n291), .A2(G20), .A3(new_n292), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT88), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n265), .A2(new_n228), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n588), .B1(new_n591), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT89), .B1(new_n596), .B2(KEYINPUT20), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n593), .B1(new_n592), .B2(new_n594), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n587), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT20), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(G116), .ZN(new_n604));
  INV_X1    g0404(.A(new_n308), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n277), .A2(new_n604), .B1(new_n274), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n600), .A2(new_n601), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(KEYINPUT89), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n586), .B1(new_n603), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n584), .A2(new_n313), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n603), .B2(new_n609), .ZN(new_n614));
  OAI211_X1 g0414(.A(KEYINPUT21), .B(new_n586), .C1(new_n603), .C2(new_n609), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n584), .A2(new_n478), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(G200), .B2(new_n584), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n596), .A2(KEYINPUT20), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n608), .A2(new_n618), .A3(KEYINPUT89), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n596), .A2(KEYINPUT20), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT89), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n606), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n612), .A2(new_n614), .A3(new_n615), .A4(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT90), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n615), .A2(new_n614), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n627), .A2(KEYINPUT90), .A3(new_n612), .A4(new_n623), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n288), .A2(G257), .A3(G1698), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT93), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT93), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n288), .A2(new_n632), .A3(G257), .A4(G1698), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n295), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n284), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n332), .B1(new_n581), .B2(new_n334), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n313), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(G169), .B2(new_n638), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n258), .A2(new_n260), .A3(new_n229), .A4(G87), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT22), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT22), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n288), .A2(new_n643), .A3(new_n229), .A4(G87), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT23), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n229), .B2(G107), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n343), .A2(KEYINPUT23), .A3(G20), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n293), .A2(new_n229), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n645), .A2(KEYINPUT91), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT91), .B1(new_n645), .B2(new_n649), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT24), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n649), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT91), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n652), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n268), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT92), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n645), .A2(KEYINPUT91), .A3(new_n649), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(KEYINPUT24), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n368), .B1(new_n651), .B2(new_n652), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n271), .A2(new_n343), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT25), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(G107), .B2(new_n278), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n640), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(G200), .B1(new_n636), .B2(new_n637), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n339), .B1(G264), .B2(new_n576), .ZN(new_n671));
  INV_X1    g0471(.A(G294), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n482), .A2(new_n210), .B1(new_n257), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n633), .B2(new_n631), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n671), .B(G190), .C1(new_n674), .C2(new_n284), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n670), .A2(new_n675), .A3(new_n668), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n662), .B1(new_n661), .B2(new_n663), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT94), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT94), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n665), .A2(new_n681), .A3(new_n676), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n669), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AND4_X1   g0483(.A1(new_n388), .A2(new_n575), .A3(new_n629), .A4(new_n683), .ZN(G372));
  NAND3_X1  g0484(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT95), .B1(new_n685), .B2(new_n669), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n615), .A2(new_n614), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n622), .A2(new_n619), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT21), .B1(new_n688), .B2(new_n586), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n668), .B1(new_n677), .B2(new_n678), .ZN(new_n691));
  INV_X1    g0491(.A(new_n640), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT95), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n680), .A2(new_n682), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n686), .A2(new_n695), .A3(new_n388), .A4(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n312), .A2(new_n317), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n385), .A2(G169), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n378), .B1(new_n699), .B2(new_n337), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT26), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n317), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n366), .A2(new_n342), .A3(new_n317), .A4(new_n312), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(KEYINPUT26), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n575), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT96), .Z(new_n708));
  AND2_X1   g0508(.A1(new_n466), .A2(new_n474), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n473), .A3(new_n521), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n572), .B1(new_n710), .B2(new_n512), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n442), .B1(new_n711), .B2(new_n566), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n526), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n708), .A2(new_n714), .ZN(G369));
  NAND3_X1  g0515(.A1(new_n275), .A2(new_n229), .A3(G13), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT27), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(KEYINPUT27), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G213), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G343), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n688), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n629), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n690), .A2(new_n722), .ZN(new_n724));
  OAI21_X1  g0524(.A(G330), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n691), .A2(new_n721), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n683), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n721), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n728), .B1(new_n693), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n690), .A2(new_n721), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n683), .A2(new_n732), .B1(new_n669), .B2(new_n729), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(G399));
  INV_X1    g0534(.A(new_n223), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G41), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n255), .A2(G116), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n736), .A2(new_n275), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n227), .B2(new_n736), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT28), .Z(new_n741));
  NAND2_X1  g0541(.A1(new_n690), .A2(new_n693), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n388), .A2(new_n742), .A3(new_n696), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT97), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n704), .A2(new_n744), .A3(new_n701), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n698), .A2(new_n700), .A3(KEYINPUT26), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n744), .B1(new_n704), .B2(new_n701), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n317), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n729), .B1(new_n743), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT29), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT29), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n706), .A2(new_n752), .A3(new_n729), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G330), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n629), .A2(new_n388), .A3(new_n683), .A4(new_n729), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n638), .A2(new_n613), .A3(new_n382), .A4(new_n316), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT30), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR4_X1   g0559(.A1(new_n638), .A2(new_n316), .A3(G179), .A4(new_n585), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n385), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n757), .A2(new_n758), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n721), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT31), .B1(new_n763), .B2(new_n721), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n755), .B1(new_n756), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n741), .B1(new_n768), .B2(G1), .ZN(G364));
  NOR2_X1   g0569(.A1(new_n221), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n275), .B1(new_n770), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n736), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n726), .A2(new_n773), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n723), .A2(new_n724), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n774), .B1(G330), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n773), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n229), .A2(new_n313), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G190), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n778), .A2(G190), .A3(new_n381), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n780), .A2(new_n781), .B1(new_n783), .B2(G322), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT100), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n478), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n229), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n229), .A2(G179), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(new_n478), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n788), .A2(G294), .B1(new_n791), .B2(G283), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n779), .A2(new_n478), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n789), .A2(G190), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n793), .A2(G326), .B1(new_n795), .B2(G303), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G190), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n778), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G311), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n789), .A2(new_n797), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n288), .B1(new_n802), .B2(G329), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n792), .A2(new_n796), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n288), .B1(new_n782), .B2(new_n201), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G77), .B2(new_n799), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n780), .A2(G68), .B1(new_n791), .B2(G107), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n787), .A2(new_n214), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n795), .A2(G87), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n806), .A2(new_n807), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  OR3_X1    g0612(.A1(new_n801), .A2(KEYINPUT32), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT32), .B1(new_n801), .B2(new_n812), .ZN(new_n814));
  INV_X1    g0614(.A(new_n793), .ZN(new_n815));
  INV_X1    g0615(.A(G50), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n813), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n785), .A2(new_n804), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n341), .A2(KEYINPUT99), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n229), .B1(KEYINPUT99), .B2(new_n341), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n228), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n777), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n735), .A2(new_n288), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n299), .B2(new_n227), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n299), .B2(new_n249), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n735), .A2(new_n346), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(G355), .B1(new_n604), .B2(new_n735), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(KEYINPUT98), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(KEYINPUT98), .ZN(new_n832));
  NOR2_X1   g0632(.A1(G13), .A2(G33), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(G20), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n822), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n835), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n823), .B1(new_n831), .B2(new_n837), .C1(new_n775), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n776), .A2(new_n839), .ZN(G396));
  NAND2_X1  g0640(.A1(new_n480), .A2(new_n729), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n706), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n721), .B1(new_n697), .B2(new_n705), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n460), .A2(new_n729), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n475), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n845), .B1(new_n475), .B2(new_n479), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n843), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n767), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n773), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n849), .A2(new_n834), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n815), .A2(new_n578), .B1(new_n794), .B2(new_n343), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n808), .B(new_n855), .C1(G283), .C2(new_n780), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n288), .B1(new_n799), .B2(new_n605), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(new_n672), .C2(new_n782), .ZN(new_n858));
  INV_X1    g0658(.A(G311), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n790), .A2(new_n209), .B1(new_n801), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT101), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(KEYINPUT102), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n783), .A2(G143), .B1(new_n799), .B2(G159), .ZN(new_n865));
  INV_X1    g0665(.A(new_n780), .ZN(new_n866));
  INV_X1    g0666(.A(G150), .ZN(new_n867));
  INV_X1    g0667(.A(G137), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n865), .B1(new_n866), .B2(new_n867), .C1(new_n868), .C2(new_n815), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT34), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n790), .A2(new_n202), .ZN(new_n873));
  INV_X1    g0673(.A(G132), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n288), .B1(new_n801), .B2(new_n874), .C1(new_n816), .C2(new_n794), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n873), .B(new_n875), .C1(G58), .C2(new_n788), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n871), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT102), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n862), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n822), .B1(new_n864), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n822), .A2(new_n833), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n880), .B(new_n773), .C1(G77), .C2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n853), .B1(new_n854), .B2(new_n883), .ZN(G384));
  NOR2_X1   g0684(.A1(new_n770), .A2(new_n275), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n719), .B1(new_n553), .B2(new_n556), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n566), .B2(new_n572), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n563), .A2(new_n557), .ZN(new_n888));
  INV_X1    g0688(.A(new_n886), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n570), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n886), .B1(new_n558), .B2(new_n569), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(new_n888), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n887), .A2(new_n895), .A3(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n848), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n511), .A2(new_n721), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n512), .A2(new_n521), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n902), .B1(new_n512), .B2(new_n521), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n901), .B(new_n846), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n756), .A2(new_n766), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n900), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT106), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n894), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n892), .A2(KEYINPUT106), .A3(new_n893), .A4(new_n888), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n891), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n887), .ZN(new_n915));
  XNOR2_X1  g0715(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n910), .B1(new_n917), .B2(new_n899), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n906), .B1(new_n756), .B2(new_n766), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n909), .A2(new_n910), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n575), .A2(new_n908), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT108), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n923), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(G330), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT109), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n522), .A2(new_n574), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n751), .B2(new_n753), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n713), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT107), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n512), .A2(new_n521), .ZN(new_n933));
  INV_X1    g0733(.A(new_n902), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n903), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n475), .A2(new_n721), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT104), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n937), .B1(new_n843), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n900), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n566), .A2(new_n719), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT39), .ZN(new_n944));
  INV_X1    g0744(.A(new_n916), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n914), .B2(new_n887), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n887), .A2(new_n895), .A3(KEYINPUT38), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n512), .A2(new_n721), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n899), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n942), .A2(new_n943), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n932), .B(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n885), .B1(new_n928), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n928), .B2(new_n953), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n375), .A2(KEYINPUT35), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n375), .A2(KEYINPUT35), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n956), .A2(new_n957), .A3(G116), .A4(new_n230), .ZN(new_n958));
  XOR2_X1   g0758(.A(KEYINPUT103), .B(KEYINPUT36), .Z(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n227), .A2(G77), .A3(new_n539), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(G50), .B2(new_n202), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(G1), .A3(new_n221), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n955), .A2(new_n960), .A3(new_n963), .ZN(G367));
  OAI221_X1 g0764(.A(new_n836), .B1(new_n223), .B2(new_n270), .C1(new_n242), .C2(new_n825), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n777), .B1(new_n965), .B2(KEYINPUT114), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(KEYINPUT114), .B2(new_n965), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n346), .B1(new_n802), .B2(G137), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n816), .B2(new_n798), .C1(new_n867), .C2(new_n782), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n866), .A2(new_n812), .B1(new_n794), .B2(new_n201), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n791), .A2(G77), .ZN(new_n971));
  INV_X1    g0771(.A(G143), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n971), .B1(new_n815), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n787), .A2(new_n202), .ZN(new_n974));
  NOR4_X1   g0774(.A1(new_n969), .A2(new_n970), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n780), .A2(G294), .B1(new_n791), .B2(G97), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n343), .B2(new_n787), .C1(new_n859), .C2(new_n815), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT46), .B1(new_n795), .B2(new_n605), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G283), .A2(new_n799), .B1(new_n802), .B2(G317), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n979), .B(new_n346), .C1(new_n578), .C2(new_n782), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n795), .A2(KEYINPUT46), .A3(G116), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT115), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n975), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT47), .Z(new_n985));
  AOI21_X1  g0785(.A(new_n967), .B1(new_n985), .B2(new_n822), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n282), .A2(new_n729), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n698), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n317), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n835), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n986), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n771), .B(KEYINPUT113), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n384), .A2(new_n387), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n699), .A2(new_n337), .B1(new_n363), .B2(new_n365), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n995), .B(new_n997), .C1(new_n378), .C2(new_n729), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n700), .A2(new_n721), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(KEYINPUT110), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT110), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n998), .A2(new_n1002), .A3(new_n999), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT112), .B1(new_n1004), .B2(new_n733), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n733), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT112), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1006), .A2(new_n1001), .A3(new_n1007), .A4(new_n1003), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1005), .A2(KEYINPUT44), .A3(new_n1008), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1004), .A2(new_n733), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1004), .A2(KEYINPUT45), .A3(new_n733), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1011), .A2(new_n1012), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n731), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n683), .A2(new_n732), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n730), .B2(new_n732), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n726), .B(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1011), .A2(new_n731), .A3(new_n1012), .A4(new_n1017), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n768), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n768), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n736), .B(KEYINPUT41), .Z(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n994), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT43), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n991), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1004), .A2(new_n669), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n997), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT111), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT111), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1035), .A3(new_n997), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n729), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1021), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT42), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1031), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(KEYINPUT43), .B2(new_n990), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1019), .A2(new_n1004), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1037), .A2(new_n1030), .A3(new_n991), .A4(new_n1039), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1046), .B(new_n1031), .C1(new_n1037), .C2(new_n1039), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1044), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1042), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n993), .B1(new_n1029), .B2(new_n1050), .ZN(G387));
  NAND2_X1  g0851(.A1(new_n1023), .A2(new_n994), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n288), .B1(new_n802), .B2(G326), .ZN(new_n1053));
  INV_X1    g0853(.A(G283), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n787), .A2(new_n1054), .B1(new_n794), .B2(new_n672), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n783), .A2(G317), .B1(new_n799), .B2(G303), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n793), .A2(G322), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n859), .C2(new_n866), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT49), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1053), .B1(new_n308), .B2(new_n790), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1061), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n403), .A2(new_n780), .B1(G68), .B2(new_n799), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT116), .Z(new_n1066));
  OAI221_X1 g0866(.A(new_n288), .B1(new_n801), .B2(new_n867), .C1(new_n782), .C2(new_n816), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n416), .A2(new_n794), .B1(new_n790), .B2(new_n214), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n270), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n788), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n815), .B2(new_n812), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n822), .B1(new_n1064), .B2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n828), .A2(new_n738), .B1(new_n343), .B2(new_n735), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n238), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n824), .B1(new_n1075), .B2(new_n299), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n449), .A2(new_n451), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n816), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT50), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n299), .B1(new_n202), .B2(new_n416), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1079), .A2(new_n738), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1074), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n777), .B1(new_n1082), .B2(new_n836), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1073), .B(new_n1083), .C1(new_n730), .C2(new_n838), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1023), .A2(new_n768), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n736), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1023), .A2(new_n768), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1052), .B(new_n1084), .C1(new_n1086), .C2(new_n1087), .ZN(G393));
  NAND2_X1  g0888(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1085), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n736), .A3(new_n1025), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1020), .A2(new_n1024), .A3(new_n994), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n246), .A2(new_n824), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n836), .B1(new_n214), .B2(new_n223), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n773), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G317), .A2(new_n793), .B1(new_n783), .B2(G311), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n866), .A2(new_n578), .B1(new_n790), .B2(new_n343), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n288), .B1(new_n802), .B2(G322), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n672), .B2(new_n798), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n787), .A2(new_n308), .B1(new_n794), .B2(new_n1054), .ZN(new_n1101));
  OR3_X1    g0901(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n794), .A2(new_n202), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n787), .A2(new_n416), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(G50), .C2(new_n780), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1077), .A2(new_n799), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n288), .B1(new_n801), .B2(new_n972), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G87), .B2(new_n791), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G150), .A2(new_n793), .B1(new_n783), .B2(G159), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT51), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1097), .A2(new_n1102), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1095), .B1(new_n1112), .B2(new_n822), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1004), .B2(new_n838), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1092), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT117), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1091), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n1091), .B2(new_n1115), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(G390));
  NAND2_X1  g0920(.A1(new_n948), .A2(new_n950), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n941), .B2(new_n949), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n949), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n946), .B2(new_n947), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n317), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n342), .A2(new_n362), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1127), .A2(new_n318), .A3(new_n701), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT26), .B1(new_n996), .B2(new_n698), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n744), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n748), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1126), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n388), .A2(new_n742), .A3(new_n696), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n721), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n938), .B1(new_n1134), .B2(new_n849), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT118), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n936), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n935), .A2(KEYINPUT118), .A3(new_n903), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1125), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n908), .A2(G330), .A3(new_n849), .A4(new_n936), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1122), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1141), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n841), .B1(new_n697), .B2(new_n705), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n936), .B1(new_n1144), .B2(new_n939), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1145), .A2(new_n1123), .B1(new_n948), .B2(new_n950), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n729), .B(new_n849), .C1(new_n743), .C2(new_n749), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n938), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1124), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1143), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1142), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1121), .A2(new_n833), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n773), .B1(new_n403), .B2(new_n882), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n782), .A2(new_n874), .B1(new_n798), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n346), .B(new_n1158), .C1(G125), .C2(new_n802), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n794), .A2(new_n867), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n780), .A2(G137), .B1(new_n791), .B2(G50), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n787), .A2(new_n812), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G128), .B2(new_n793), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1104), .B1(G283), .B2(new_n793), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n343), .B2(new_n866), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n798), .A2(new_n214), .B1(new_n801), .B2(new_n672), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n288), .B(new_n1168), .C1(G116), .C2(new_n783), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n873), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n810), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1165), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1156), .B1(new_n1172), .B2(new_n822), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1154), .A2(new_n994), .B1(new_n1155), .B2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n575), .A2(G330), .A3(new_n908), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n930), .A2(new_n713), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1150), .B1(new_n767), .B2(new_n849), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1144), .A2(new_n939), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n908), .A2(G330), .A3(new_n849), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n937), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1180), .B1(new_n1182), .B2(new_n1141), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1176), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1153), .A2(new_n1184), .A3(KEYINPUT119), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n936), .B1(new_n767), .B2(new_n849), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n1143), .A2(new_n1186), .B1(new_n1144), .B2(new_n939), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1139), .A2(new_n1181), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n1135), .A3(new_n1141), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1190), .A2(new_n1142), .A3(new_n1152), .A4(new_n1176), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1185), .A2(new_n736), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT119), .B1(new_n1153), .B2(new_n1184), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1174), .B1(new_n1192), .B2(new_n1193), .ZN(G378));
  NAND2_X1  g0994(.A1(new_n909), .A2(new_n910), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n918), .A2(new_n919), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(G330), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n442), .A2(new_n526), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n719), .B1(new_n411), .B2(new_n394), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1197), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n920), .B2(G330), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n952), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1197), .A2(new_n1207), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n952), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n920), .A2(G330), .A3(new_n1209), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n773), .B1(G50), .B2(new_n882), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n815), .A2(new_n604), .B1(new_n790), .B2(new_n201), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G97), .B2(new_n780), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n346), .A2(new_n283), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G283), .B2(new_n802), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n783), .A2(G107), .B1(new_n799), .B2(new_n1069), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n974), .B1(G77), .B2(new_n795), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1219), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT58), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1220), .B(new_n816), .C1(G33), .C2(G41), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n793), .A2(G125), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n866), .B2(new_n874), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n783), .A2(G128), .B1(new_n799), .B2(G137), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n794), .B2(new_n1157), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(G150), .C2(new_n788), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n791), .A2(G159), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G33), .B(G41), .C1(new_n802), .C2(G124), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1228), .B1(new_n1225), .B2(new_n1224), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1217), .B1(new_n1240), .B2(new_n822), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1209), .B2(new_n834), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT120), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT120), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1216), .A2(new_n994), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1191), .A2(new_n1176), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1216), .A2(new_n1246), .A3(KEYINPUT57), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n736), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT57), .B1(new_n1216), .B2(new_n1246), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1245), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT121), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(KEYINPUT121), .B(new_n1245), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1253), .A2(new_n1255), .ZN(G375));
  NAND2_X1  g1056(.A1(new_n754), .A2(new_n575), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1175), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n714), .A3(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1184), .A3(new_n1028), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1139), .A2(new_n833), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n773), .B1(G68), .B2(new_n882), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n787), .A2(new_n816), .B1(new_n794), .B2(new_n812), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G132), .B2(new_n793), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n346), .B1(new_n802), .B2(G128), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n783), .A2(G137), .B1(new_n799), .B2(G150), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1157), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n780), .A2(new_n1268), .B1(new_n791), .B2(G58), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n346), .B1(new_n782), .B2(new_n1054), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G107), .B2(new_n799), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n605), .A2(new_n780), .B1(new_n793), .B2(G294), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n971), .A4(new_n1070), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n794), .A2(new_n214), .B1(new_n801), .B2(new_n578), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(KEYINPUT122), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1270), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1263), .B1(new_n1277), .B2(new_n822), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1190), .A2(new_n994), .B1(new_n1262), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1261), .A2(new_n1279), .ZN(G381));
  AND2_X1   g1080(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1027), .B1(new_n1025), .B2(new_n768), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n994), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1091), .A2(new_n1115), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT117), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1091), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n1285), .A3(new_n993), .A4(new_n1286), .ZN(new_n1287));
  OR2_X1    g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  OR3_X1    g1088(.A1(new_n1288), .A2(G384), .A3(G381), .ZN(new_n1289));
  OR3_X1    g1089(.A1(new_n1287), .A2(new_n1289), .A3(KEYINPUT123), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT123), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G375), .A2(KEYINPUT125), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G378), .A2(KEYINPUT124), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT124), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1295), .B(new_n1174), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1292), .A2(new_n1293), .A3(new_n1297), .A4(new_n1299), .ZN(G407));
  NAND2_X1  g1100(.A1(new_n720), .A2(G213), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1293), .A2(new_n1297), .A3(new_n1299), .A4(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(G407), .A2(new_n1303), .A3(G213), .ZN(G409));
  NAND3_X1  g1104(.A1(new_n1216), .A2(new_n1246), .A3(new_n1028), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1245), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1294), .A2(new_n1296), .A3(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G378), .B(new_n1245), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1260), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1259), .A2(new_n1187), .A3(KEYINPUT60), .A4(new_n1189), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1311), .A2(new_n736), .A3(new_n1184), .A4(new_n1312), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1313), .A2(G384), .A3(new_n1279), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G384), .B1(new_n1313), .B2(new_n1279), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1309), .A2(new_n1301), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1309), .A2(new_n1301), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT126), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1314), .A2(new_n1315), .A3(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1320), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1322));
  INV_X1    g1122(.A(G2897), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1301), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  OAI221_X1 g1125(.A(new_n1320), .B1(new_n1323), .B2(new_n1301), .C1(new_n1314), .C2(new_n1315), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1321), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1319), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1309), .A2(new_n1330), .A3(new_n1301), .A4(new_n1316), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1318), .A2(new_n1328), .A3(new_n1329), .A4(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(G396), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(G393), .B(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1334), .A2(KEYINPUT127), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n993), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1029), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1336), .B1(new_n1337), .B2(new_n1281), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1335), .B1(new_n1119), .B2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(G387), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1334), .A2(KEYINPUT127), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1339), .A2(new_n1342), .A3(new_n1340), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1332), .A2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1342), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1335), .ZN(new_n1349));
  AND4_X1   g1149(.A1(new_n1287), .A2(new_n1340), .A3(new_n1349), .A4(new_n1342), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1348), .A2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(KEYINPUT61), .B1(new_n1319), .B2(new_n1327), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1309), .A2(KEYINPUT63), .A3(new_n1301), .A4(new_n1316), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT63), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1317), .A2(new_n1354), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1351), .A2(new_n1352), .A3(new_n1353), .A4(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1347), .A2(new_n1356), .ZN(G405));
  NAND3_X1  g1157(.A1(new_n1252), .A2(new_n1297), .A3(new_n1254), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1316), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1358), .A2(new_n1308), .A3(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1359), .B1(new_n1358), .B2(new_n1308), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1346), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1362), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1351), .A2(new_n1364), .A3(new_n1360), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1363), .A2(new_n1365), .ZN(G402));
endmodule


