//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(new_n464), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n472), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G101), .A2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n478), .B1(new_n469), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(KEYINPUT70), .A3(new_n481), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n477), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  NOR2_X1   g063(.A1(new_n469), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n469), .A2(new_n481), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  OR3_X1    g067(.A1(KEYINPUT71), .A2(G100), .A3(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n481), .A2(G112), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT71), .B1(G100), .B2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n493), .A2(new_n494), .A3(G2104), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n490), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  NAND3_X1  g073(.A1(new_n465), .A2(KEYINPUT4), .A3(G138), .ZN(new_n499));
  NAND2_X1  g074(.A1(G102), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(G2105), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n462), .A2(new_n464), .A3(G126), .ZN(new_n502));
  NAND2_X1  g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n481), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n489), .A2(G138), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(G164));
  AND2_X1   g083(.A1(KEYINPUT72), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT72), .A2(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT6), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT73), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(KEYINPUT73), .A3(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n514), .A2(G88), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n516), .A2(new_n518), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT72), .B(G651), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n511), .A2(G50), .A3(G543), .A4(new_n513), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n520), .A2(new_n527), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n511), .A2(new_n513), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n514), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n534), .B(new_n536), .C1(new_n537), .C2(new_n522), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  AOI22_X1  g114(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n525), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n531), .A2(new_n522), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n533), .A2(G52), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n522), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(new_n526), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n511), .A2(G43), .A3(G543), .A4(new_n513), .ZN(new_n551));
  XNOR2_X1  g126(.A(KEYINPUT74), .B(G81), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n519), .A2(new_n511), .A3(new_n513), .A4(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n542), .A2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n522), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n511), .A2(G53), .A3(G543), .A4(new_n513), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n562), .B(new_n566), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT75), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n567), .B(KEYINPUT9), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n572), .A2(new_n573), .A3(new_n562), .A4(new_n566), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G299));
  OAI21_X1  g150(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n519), .A2(G87), .A3(new_n511), .A4(new_n513), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n511), .A2(G49), .A3(G543), .A4(new_n513), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  INV_X1    g155(.A(G73), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n531), .A2(new_n580), .B1(new_n581), .B2(new_n525), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n531), .A2(new_n584), .B1(new_n585), .B2(new_n525), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(new_n519), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n525), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n542), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n533), .A2(G47), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT76), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n516), .A2(new_n518), .A3(G66), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n512), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G54), .ZN(new_n599));
  NOR3_X1   g174(.A1(new_n531), .A2(new_n599), .A3(new_n532), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n519), .A2(new_n511), .A3(new_n513), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n514), .A2(KEYINPUT10), .A3(G92), .A4(new_n519), .ZN(new_n605));
  AOI211_X1 g180(.A(new_n598), .B(new_n600), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n594), .B1(new_n606), .B2(G868), .ZN(G321));
  XOR2_X1   g182(.A(G321), .B(KEYINPUT77), .Z(G284));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT78), .Z(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g194(.A1(new_n481), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT79), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT80), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G2100), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n624), .A2(G2100), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n481), .A2(G111), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n461), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI221_X1 g205(.A(new_n630), .B1(new_n629), .B2(new_n628), .C1(G99), .C2(G2105), .ZN(new_n631));
  AOI22_X1  g206(.A1(G123), .A2(new_n491), .B1(new_n489), .B2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT82), .B(G2096), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n627), .B(new_n635), .C1(new_n625), .C2(new_n623), .ZN(G156));
  INV_X1    g211(.A(G14), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT83), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n647), .A2(new_n651), .A3(new_n648), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n637), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n647), .A2(new_n648), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT17), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n664), .C2(new_n660), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT20), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  OR3_X1    g256(.A1(new_n674), .A2(new_n677), .A3(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT85), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1981), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(G229));
  AOI22_X1  g265(.A1(G129), .A2(new_n491), .B1(new_n489), .B2(G141), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n481), .A2(G105), .A3(G2104), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT97), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT98), .B(KEYINPUT26), .ZN(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  AND3_X1   g271(.A1(new_n691), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G29), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G29), .B2(G32), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT27), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G26), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n491), .A2(G128), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT90), .ZN(new_n705));
  OR2_X1    g280(.A1(G104), .A2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n706), .B(G2104), .C1(G116), .C2(new_n481), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n489), .A2(G140), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n703), .B1(new_n710), .B2(new_n702), .ZN(new_n711));
  MUX2_X1   g286(.A(new_n703), .B(new_n711), .S(KEYINPUT28), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT91), .B(G2067), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G4), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n606), .B2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1348), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n715), .A2(G19), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n719), .B(new_n720), .C1(new_n554), .C2(G16), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n719), .B2(new_n720), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT89), .B(G1341), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n715), .A2(G21), .ZN(new_n725));
  INV_X1    g300(.A(G1966), .ZN(new_n726));
  OAI221_X1 g301(.A(new_n725), .B1(KEYINPUT101), .B2(new_n726), .C1(G168), .C2(new_n715), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT101), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n727), .A2(new_n728), .A3(G1966), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n715), .A2(G5), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G171), .B2(new_n715), .ZN(new_n731));
  INV_X1    g306(.A(G1961), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n728), .B2(G1966), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n724), .A2(new_n729), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT31), .B(G11), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT99), .ZN(new_n737));
  INV_X1    g312(.A(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT30), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(KEYINPUT30), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n739), .A2(new_n740), .A3(new_n702), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n737), .B(new_n741), .C1(new_n633), .C2(new_n702), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT100), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n702), .A2(G35), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G162), .B2(new_n702), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT29), .B(G2090), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n702), .A2(G27), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G164), .B2(new_n702), .ZN(new_n750));
  INV_X1    g325(.A(G2078), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT24), .B(G34), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(G29), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n487), .B2(G29), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n748), .B(new_n752), .C1(new_n753), .C2(new_n756), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n714), .A2(new_n718), .A3(new_n735), .A4(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(new_n481), .ZN(new_n760));
  AND3_X1   g335(.A1(new_n465), .A2(G139), .A3(new_n481), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT92), .B(KEYINPUT93), .Z(new_n764));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(KEYINPUT25), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n763), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n764), .A2(new_n765), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n767), .A2(KEYINPUT25), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n770), .A2(new_n762), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n761), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(KEYINPUT94), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n775), .B(new_n761), .C1(new_n769), .C2(new_n772), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n760), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(KEYINPUT95), .ZN(new_n778));
  INV_X1    g353(.A(new_n761), .ZN(new_n779));
  INV_X1    g354(.A(new_n772), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n762), .B1(new_n770), .B2(new_n771), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(new_n775), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n773), .A2(KEYINPUT94), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n785), .A2(new_n786), .A3(new_n760), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n702), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n702), .B2(G33), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT96), .B(G2072), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n715), .A2(G20), .ZN(new_n792));
  OAI211_X1 g367(.A(KEYINPUT23), .B(new_n792), .C1(new_n610), .C2(new_n715), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(KEYINPUT23), .B2(new_n792), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1956), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n756), .A2(new_n753), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT102), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n758), .A2(new_n791), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n715), .A2(G23), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n715), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT86), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n715), .A2(G6), .ZN(new_n805));
  INV_X1    g380(.A(G305), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n715), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n802), .A2(new_n803), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n715), .A2(G22), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G166), .B2(new_n715), .ZN(new_n812));
  INV_X1    g387(.A(G1971), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n804), .A2(new_n809), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT87), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n817));
  INV_X1    g392(.A(G290), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n715), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n715), .B2(G24), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(G1986), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n491), .A2(G119), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n489), .A2(G131), .ZN(new_n825));
  NOR2_X1   g400(.A1(G95), .A2(G2105), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(new_n481), .B2(G107), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  MUX2_X1   g403(.A(G25), .B(new_n828), .S(G29), .Z(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT35), .B(G1991), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n821), .B2(G1986), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n817), .A2(new_n822), .A3(new_n823), .A4(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(KEYINPUT36), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(KEYINPUT36), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n701), .B(new_n798), .C1(new_n834), .C2(new_n835), .ZN(G311));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  INV_X1    g412(.A(new_n701), .ZN(new_n838));
  INV_X1    g413(.A(new_n798), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(G150));
  NAND3_X1  g415(.A1(new_n514), .A2(G93), .A3(new_n519), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n514), .A2(G55), .A3(G543), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n516), .A2(new_n518), .A3(G67), .ZN(new_n844));
  NAND2_X1  g419(.A1(G80), .A2(G543), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n843), .B1(new_n846), .B2(new_n526), .ZN(new_n847));
  AOI211_X1 g422(.A(KEYINPUT103), .B(new_n525), .C1(new_n844), .C2(new_n845), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n841), .B(new_n842), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  AOI21_X1  g426(.A(new_n525), .B1(new_n844), .B2(new_n845), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n843), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n853), .A2(new_n554), .A3(new_n841), .A4(new_n842), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n849), .A2(new_n555), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT39), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n606), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n851), .B1(new_n860), .B2(G860), .ZN(G145));
  XNOR2_X1  g436(.A(new_n697), .B(KEYINPUT105), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n487), .B(new_n497), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n828), .B(KEYINPUT106), .Z(new_n864));
  INV_X1    g439(.A(G164), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n778), .A2(new_n787), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n778), .B2(new_n787), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n481), .A2(G118), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n461), .B1(new_n869), .B2(KEYINPUT104), .ZN(new_n870));
  OAI221_X1 g445(.A(new_n870), .B1(KEYINPUT104), .B2(new_n869), .C1(G106), .C2(G2105), .ZN(new_n871));
  AOI22_X1  g446(.A1(G130), .A2(new_n491), .B1(new_n489), .B2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n709), .B(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n777), .A2(KEYINPUT95), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n786), .B1(new_n785), .B2(new_n760), .ZN(new_n876));
  OAI21_X1  g451(.A(G164), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n864), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n778), .A2(new_n787), .A3(new_n865), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n868), .A2(new_n874), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n874), .B1(new_n868), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n863), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n633), .B(new_n621), .ZN(new_n884));
  INV_X1    g459(.A(new_n874), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n866), .A2(new_n867), .A3(new_n864), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n868), .A2(new_n880), .A3(new_n874), .ZN(new_n889));
  INV_X1    g464(.A(new_n863), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n883), .A2(new_n884), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n884), .B1(new_n883), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n862), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  INV_X1    g470(.A(new_n884), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n881), .A2(new_n882), .A3(new_n863), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n890), .B1(new_n888), .B2(new_n889), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n862), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n883), .A2(new_n884), .A3(new_n891), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n894), .A2(new_n895), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT40), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n894), .A2(new_n905), .A3(new_n902), .A4(new_n895), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(G395));
  NOR2_X1   g482(.A1(new_n849), .A2(G868), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n616), .B(new_n856), .ZN(new_n909));
  INV_X1    g484(.A(new_n606), .ZN(new_n910));
  NAND2_X1  g485(.A1(G299), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n571), .A2(new_n574), .A3(new_n606), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n911), .A2(KEYINPUT107), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT107), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n912), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n571), .A2(new_n574), .A3(new_n606), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n606), .B1(new_n571), .B2(new_n574), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n909), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n916), .A2(KEYINPUT108), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(G303), .A2(new_n800), .ZN(new_n924));
  NAND4_X1  g499(.A1(G288), .A2(new_n527), .A3(new_n520), .A4(new_n528), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(G305), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G305), .B1(new_n924), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g503(.A(G290), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(new_n818), .A3(new_n926), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT42), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n923), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT108), .B1(new_n916), .B2(new_n922), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n935), .B(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n908), .B1(new_n937), .B2(G868), .ZN(G295));
  AOI21_X1  g513(.A(new_n908), .B1(new_n937), .B2(G868), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n854), .A2(new_n855), .A3(G301), .ZN(new_n941));
  AOI21_X1  g516(.A(G301), .B1(new_n854), .B2(new_n855), .ZN(new_n942));
  OAI21_X1  g517(.A(G286), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n849), .A2(new_n555), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n849), .A2(new_n555), .ZN(new_n945));
  OAI21_X1  g520(.A(G171), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n854), .A2(new_n855), .A3(G301), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(G168), .A3(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n943), .A2(new_n948), .A3(new_n911), .A4(new_n912), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n941), .A2(new_n942), .A3(G286), .ZN(new_n950));
  AOI21_X1  g525(.A(G168), .B1(new_n946), .B2(new_n947), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n921), .A2(new_n917), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n932), .B(new_n949), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT110), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n917), .B(new_n921), .C1(new_n950), .C2(new_n951), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n956), .A2(new_n957), .A3(new_n932), .A4(new_n949), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n943), .A2(new_n948), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n915), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n932), .B(KEYINPUT109), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n940), .B1(new_n964), .B2(KEYINPUT43), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  AOI211_X1 g541(.A(KEYINPUT111), .B(new_n966), .C1(new_n959), .C2(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n956), .A2(new_n949), .ZN(new_n968));
  AOI21_X1  g543(.A(G37), .B1(new_n962), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n959), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT44), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n965), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n959), .A2(new_n969), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n959), .A2(new_n966), .A3(new_n963), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT44), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT112), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n975), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT111), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n964), .A2(new_n940), .A3(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n978), .B(new_n981), .C1(new_n985), .C2(new_n971), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n977), .A2(new_n986), .ZN(G397));
  NAND3_X1  g562(.A1(new_n484), .A2(G40), .A3(new_n485), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n475), .B2(new_n476), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n499), .A2(new_n500), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n481), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n507), .B1(new_n505), .B2(new_n504), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(G1996), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT113), .ZN(new_n997));
  INV_X1    g572(.A(new_n995), .ZN(new_n998));
  INV_X1    g573(.A(G2067), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n710), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n709), .A2(G2067), .ZN(new_n1001));
  INV_X1    g576(.A(G1996), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1000), .B(new_n1001), .C1(new_n1002), .C2(new_n697), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n997), .A2(new_n697), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n828), .A2(new_n830), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n828), .A2(new_n830), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n998), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(G290), .B(G1986), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n998), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(G305), .A2(G1981), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G305), .A2(G1981), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1013), .A2(KEYINPUT49), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n484), .A2(G40), .A3(new_n485), .ZN(new_n1015));
  INV_X1    g590(.A(new_n476), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT69), .B1(new_n472), .B2(G2105), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1015), .B(new_n993), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(KEYINPUT49), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1014), .A2(G8), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(G8), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(G1976), .B2(new_n800), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1022), .B(new_n1023), .C1(G1976), .C2(new_n800), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1020), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n993), .A2(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1028), .A2(new_n989), .A3(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT114), .B(G2090), .Z(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(G164), .B2(G1384), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n993), .A2(KEYINPUT45), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n989), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n813), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1027), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G303), .A2(G8), .ZN(new_n1040));
  XOR2_X1   g615(.A(new_n1040), .B(KEYINPUT55), .Z(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1026), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1035), .A2(new_n989), .A3(new_n751), .A4(new_n1036), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1046));
  NAND3_X1  g621(.A1(new_n1028), .A2(new_n989), .A3(new_n1030), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1045), .A2(new_n1046), .B1(new_n1047), .B2(new_n732), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G171), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1015), .B(new_n473), .C1(new_n993), .C2(KEYINPUT45), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT123), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT123), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1035), .A2(new_n1056), .A3(new_n473), .A4(new_n1015), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1049), .B1(KEYINPUT124), .B2(new_n751), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n751), .A2(KEYINPUT124), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n993), .B2(KEYINPUT45), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1048), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1052), .B(new_n1053), .C1(G171), .C2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT125), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1062), .B2(G171), .ZN(new_n1065));
  AOI211_X1 g640(.A(KEYINPUT125), .B(G301), .C1(new_n1048), .C2(new_n1061), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1048), .A2(new_n1050), .A3(G301), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1063), .B1(new_n1068), .B2(new_n1053), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G286), .A2(G8), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT121), .ZN(new_n1071));
  AND2_X1   g646(.A1(KEYINPUT116), .A2(G2084), .ZN(new_n1072));
  NOR2_X1   g647(.A1(KEYINPUT116), .A2(G2084), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1031), .A2(new_n1074), .B1(new_n1037), .B2(new_n726), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1071), .B1(new_n1075), .B2(new_n1027), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1071), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1047), .A2(new_n1073), .A3(new_n1072), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1037), .A2(new_n726), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1077), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1079), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1035), .A2(new_n989), .A3(new_n1002), .A4(new_n1036), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT58), .B(G1341), .Z(new_n1088));
  NAND2_X1  g663(.A1(new_n1018), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n554), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1086), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n1091), .B2(new_n1090), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT61), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT118), .B(G1956), .Z(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1047), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n570), .B(KEYINPUT57), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1035), .A2(new_n989), .A3(new_n1036), .A4(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1099), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1094), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1098), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1108));
  OR3_X1    g683(.A1(new_n1090), .A2(new_n1091), .A3(KEYINPUT59), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1093), .A2(new_n1105), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1348), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1047), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1018), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n999), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT120), .B1(new_n1115), .B2(new_n910), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1111), .A2(new_n1047), .B1(new_n1113), .B2(new_n999), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1117), .A2(KEYINPUT60), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1119), .B(new_n606), .C1(new_n1117), .C2(KEYINPUT60), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1116), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1110), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1117), .A2(new_n910), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1103), .B1(new_n1124), .B2(new_n1107), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1069), .B(new_n1085), .C1(new_n1123), .C2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1084), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT126), .ZN(new_n1128));
  OR3_X1    g703(.A1(new_n1079), .A2(new_n1084), .A3(KEYINPUT62), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1052), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1131), .B(KEYINPUT62), .C1(new_n1079), .C2(new_n1084), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1044), .B1(new_n1126), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1075), .A2(new_n1027), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1026), .A2(new_n1043), .A3(new_n1042), .A4(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(KEYINPUT117), .A2(KEYINPUT63), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  OR3_X1    g713(.A1(new_n1136), .A2(G286), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(KEYINPUT117), .A2(KEYINPUT63), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1140), .B(new_n1138), .C1(new_n1136), .C2(G286), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1026), .A2(new_n1041), .A3(new_n1039), .ZN(new_n1142));
  INV_X1    g717(.A(G1976), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1020), .A2(new_n1143), .A3(new_n800), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1011), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1021), .B(KEYINPUT115), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .A4(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1010), .B1(new_n1134), .B2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1004), .A2(new_n1005), .B1(new_n999), .B2(new_n710), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n995), .A2(G1986), .A3(G290), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT48), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1150), .A2(new_n995), .B1(new_n1008), .B2(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n997), .B(KEYINPUT46), .Z(new_n1154));
  AND3_X1   g729(.A1(new_n1000), .A2(new_n1001), .A3(new_n697), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n995), .B2(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1156), .A2(KEYINPUT47), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(KEYINPUT47), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1153), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1149), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g735(.A(new_n459), .B1(new_n653), .B2(new_n654), .ZN(new_n1162));
  INV_X1    g736(.A(G227), .ZN(new_n1163));
  AND3_X1   g737(.A1(new_n1162), .A2(KEYINPUT127), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g738(.A(KEYINPUT127), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1165));
  NOR3_X1   g739(.A1(new_n1164), .A2(new_n1165), .A3(G229), .ZN(new_n1166));
  AND3_X1   g740(.A1(new_n1166), .A2(new_n903), .A3(new_n979), .ZN(G308));
  NAND3_X1  g741(.A1(new_n1166), .A2(new_n903), .A3(new_n979), .ZN(G225));
endmodule


