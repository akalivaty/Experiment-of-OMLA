//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(G116), .B(G119), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n191));
  INV_X1    g005(.A(G113), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n191), .A2(new_n192), .A3(KEYINPUT70), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT70), .B1(new_n191), .B2(new_n192), .ZN(new_n194));
  OR2_X1    g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT2), .A2(G113), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n190), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n190), .B(new_n196), .C1(new_n193), .C2(new_n194), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(G104), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n205), .A2(G107), .B1(KEYINPUT78), .B2(KEYINPUT3), .ZN(new_n206));
  OAI22_X1  g020(.A1(new_n205), .A2(G107), .B1(KEYINPUT78), .B2(KEYINPUT3), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT4), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(G101), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n204), .A2(new_n206), .A3(new_n207), .A4(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(KEYINPUT4), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n201), .A2(new_n210), .A3(new_n214), .ZN(new_n215));
  XOR2_X1   g029(.A(G110), .B(G122), .Z(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n218));
  INV_X1    g032(.A(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G116), .ZN(new_n220));
  OAI21_X1  g034(.A(G113), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G116), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G119), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT5), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT83), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT83), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT5), .ZN(new_n227));
  AND4_X1   g041(.A1(new_n220), .A2(new_n223), .A3(new_n225), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT84), .B1(new_n221), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n227), .ZN(new_n230));
  INV_X1    g044(.A(new_n220), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n192), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT84), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n190), .A2(new_n218), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n229), .A2(new_n198), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n203), .A2(G104), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n205), .A2(G107), .ZN(new_n238));
  OAI21_X1  g052(.A(G101), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n213), .A2(new_n239), .ZN(new_n240));
  OR2_X1    g054(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n215), .A2(new_n217), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n240), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT88), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n220), .A2(new_n223), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT87), .B1(new_n245), .B2(new_n224), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT87), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n190), .A2(new_n247), .A3(KEYINPUT5), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n246), .A2(new_n232), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n198), .A2(new_n213), .A3(new_n239), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n232), .A3(new_n248), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n213), .A2(new_n239), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT88), .A4(new_n198), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n243), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n216), .B(KEYINPUT8), .Z(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  XNOR2_X1  g071(.A(G143), .B(G146), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(KEYINPUT65), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  INV_X1    g075(.A(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT0), .B(G128), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT75), .B(G125), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n259), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(KEYINPUT1), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n261), .A3(new_n263), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT69), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n260), .A2(G146), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n262), .A2(G143), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G128), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n270), .A2(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n271), .A2(new_n261), .A3(new_n263), .A4(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n269), .B1(new_n281), .B2(new_n268), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT85), .B(G224), .ZN(new_n283));
  INV_X1    g097(.A(G953), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(KEYINPUT7), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n282), .A2(KEYINPUT89), .A3(KEYINPUT7), .A4(new_n285), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n255), .A2(new_n256), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT90), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n242), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n255), .A2(new_n256), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n291), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n295), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n189), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT91), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n215), .A2(new_n241), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n216), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT6), .A3(new_n242), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT6), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n304), .A3(new_n216), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n285), .B(KEYINPUT86), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n282), .B(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(KEYINPUT91), .B(new_n189), .C1(new_n294), .C2(new_n297), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n300), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n300), .A2(new_n311), .A3(new_n308), .A4(new_n309), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n188), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT23), .B1(new_n270), .B2(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n270), .A2(G119), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(KEYINPUT74), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT74), .B1(new_n219), .B2(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n219), .A2(G128), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(KEYINPUT23), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G110), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n320), .A2(new_n317), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT24), .B(G110), .Z(new_n325));
  OAI21_X1  g139(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(G140), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n268), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(G125), .A2(G140), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(new_n268), .B2(G140), .ZN(new_n331));
  OAI211_X1 g145(.A(G146), .B(new_n329), .C1(new_n331), .C2(new_n327), .ZN(new_n332));
  XNOR2_X1  g146(.A(G125), .B(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n262), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n326), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n322), .B1(new_n318), .B2(new_n321), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n324), .B2(new_n325), .ZN(new_n339));
  INV_X1    g153(.A(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT75), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G125), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n343), .A3(G140), .ZN(new_n344));
  INV_X1    g158(.A(new_n330), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n327), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(G146), .B1(new_n347), .B2(new_n329), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n341), .A2(new_n343), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n349), .A2(KEYINPUT16), .A3(G140), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n346), .A2(new_n350), .A3(new_n262), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n339), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n326), .A2(new_n332), .A3(KEYINPUT76), .A4(new_n334), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n337), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n284), .A2(G221), .A3(G234), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT22), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(G137), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n337), .A2(new_n352), .A3(new_n353), .A4(new_n357), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n189), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT25), .ZN(new_n362));
  INV_X1    g176(.A(G217), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(G234), .B2(new_n189), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n359), .A2(new_n365), .A3(new_n189), .A4(new_n360), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n359), .A2(new_n360), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n364), .A2(G902), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n259), .A2(new_n267), .ZN(new_n373));
  INV_X1    g187(.A(G131), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT11), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT66), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT66), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT11), .ZN(new_n378));
  INV_X1    g192(.A(G137), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n376), .A2(new_n378), .B1(G134), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n377), .A2(KEYINPUT11), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(G134), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT67), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n379), .B2(G134), .ZN(new_n386));
  INV_X1    g200(.A(G134), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT67), .A3(G137), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n374), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n375), .A2(KEYINPUT66), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n382), .B1(new_n381), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n376), .A2(G134), .A3(new_n379), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n392), .A2(new_n374), .A3(new_n389), .A4(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n373), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n379), .A2(KEYINPUT68), .A3(G134), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(G134), .B2(new_n379), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT68), .B1(new_n379), .B2(G134), .ZN(new_n399));
  OAI21_X1  g213(.A(G131), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n281), .A2(new_n394), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT71), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT71), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n281), .A2(new_n403), .A3(new_n394), .A4(new_n400), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n396), .A2(new_n402), .A3(KEYINPUT30), .A4(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n392), .A2(new_n389), .A3(new_n393), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G131), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n408), .A2(new_n394), .B1(new_n267), .B2(new_n259), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n281), .A2(new_n394), .A3(new_n400), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n405), .A2(new_n201), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G237), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT72), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT72), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G237), .ZN(new_n416));
  AOI21_X1  g230(.A(G953), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G210), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT26), .B(G101), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n396), .A2(new_n402), .A3(new_n200), .A4(new_n404), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n412), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT31), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n396), .A2(new_n200), .A3(new_n401), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n201), .B1(new_n409), .B2(new_n410), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n428), .B(new_n429), .C1(new_n427), .C2(new_n423), .ZN(new_n430));
  INV_X1    g244(.A(new_n422), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT31), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n412), .A2(new_n433), .A3(new_n422), .A4(new_n423), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n425), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(G472), .A2(G902), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT32), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT32), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n439), .A3(new_n436), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n428), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n396), .A2(new_n402), .A3(new_n404), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n201), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n423), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n442), .B1(new_n445), .B2(KEYINPUT28), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n431), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(G902), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n412), .A2(new_n423), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n431), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n423), .A2(new_n427), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n452), .A2(new_n422), .A3(new_n429), .A4(new_n428), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n453), .A3(new_n447), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G472), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n372), .B1(new_n441), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G113), .B(G122), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(G104), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT95), .ZN(new_n462));
  AOI21_X1  g276(.A(G143), .B1(new_n417), .B2(G214), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n417), .A2(G143), .A3(G214), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT18), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n374), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n331), .A2(G146), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n334), .ZN(new_n469));
  INV_X1    g283(.A(new_n465), .ZN(new_n470));
  OAI21_X1  g284(.A(G131), .B1(new_n470), .B2(new_n463), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n467), .B(new_n469), .C1(new_n466), .C2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n348), .A2(new_n351), .ZN(new_n473));
  OAI211_X1 g287(.A(KEYINPUT17), .B(G131), .C1(new_n470), .C2(new_n463), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n464), .A2(new_n374), .A3(new_n465), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n473), .B(new_n474), .C1(new_n476), .C2(KEYINPUT17), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n462), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n344), .A2(KEYINPUT19), .A3(new_n345), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT19), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n333), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n479), .A2(new_n262), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT92), .B1(new_n351), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n481), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n332), .B(new_n484), .C1(G146), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n476), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n472), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT94), .B1(new_n488), .B2(new_n461), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT94), .ZN(new_n490));
  INV_X1    g304(.A(new_n461), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n490), .B(new_n491), .C1(new_n487), .C2(new_n472), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n478), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G475), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n189), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT20), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G478), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(KEYINPUT15), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n222), .A2(G122), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n222), .A2(G122), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n503), .A2(new_n203), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n203), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT97), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT98), .B1(new_n270), .B2(G143), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT98), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n260), .A3(G128), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n270), .A2(G143), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT13), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n387), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n515), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT97), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n504), .A2(new_n518), .A3(new_n505), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n507), .A2(new_n516), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT99), .B1(new_n502), .B2(KEYINPUT14), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n502), .A2(KEYINPUT14), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT99), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n222), .A4(G122), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n521), .A2(new_n501), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G107), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n513), .A2(G134), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n387), .B1(new_n511), .B2(new_n512), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n527), .B(new_n505), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n530), .A2(KEYINPUT100), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(KEYINPUT100), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n520), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT9), .B(G234), .Z(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(G217), .A3(new_n284), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n520), .B(new_n537), .C1(new_n531), .C2(new_n532), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n500), .B1(new_n539), .B2(new_n189), .ZN(new_n540));
  AOI211_X1 g354(.A(G902), .B(new_n499), .C1(new_n536), .C2(new_n538), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n493), .A2(KEYINPUT20), .A3(new_n494), .A4(new_n189), .ZN(new_n543));
  INV_X1    g357(.A(new_n478), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n491), .B1(new_n477), .B2(new_n472), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n189), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT96), .B(G475), .Z(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n497), .A2(new_n542), .A3(new_n543), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n284), .A2(G952), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(G234), .B2(G237), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI211_X1 g366(.A(new_n189), .B(new_n284), .C1(G234), .C2(G237), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(KEYINPUT21), .B(G898), .Z(new_n555));
  OAI21_X1  g369(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n556), .B(KEYINPUT101), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n549), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT82), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n253), .A2(new_n281), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n240), .A2(new_n278), .A3(new_n273), .A4(new_n280), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n408), .A2(new_n394), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT12), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT12), .B1(new_n563), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT81), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(KEYINPUT79), .A2(KEYINPUT10), .ZN(new_n569));
  NOR2_X1   g383(.A1(KEYINPUT79), .A2(KEYINPUT10), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n569), .B1(new_n561), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n390), .A2(new_n395), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n214), .A2(new_n373), .A3(new_n210), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n253), .A2(new_n281), .A3(KEYINPUT79), .A4(KEYINPUT10), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(G110), .B(G140), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n284), .A2(G227), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n281), .B(new_n240), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n572), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT81), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n565), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n568), .A2(new_n575), .A3(new_n578), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n564), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n575), .ZN(new_n587));
  INV_X1    g401(.A(new_n578), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT80), .B(G469), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n586), .A2(new_n575), .A3(new_n578), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n581), .A2(new_n565), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n578), .B1(new_n593), .B2(new_n575), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n189), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n590), .A2(new_n591), .B1(new_n595), .B2(G469), .ZN(new_n596));
  INV_X1    g410(.A(G221), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n534), .B2(new_n189), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT77), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n560), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n584), .A2(new_n589), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(new_n189), .A3(new_n591), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n595), .A2(G469), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(KEYINPUT82), .A3(new_n599), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n315), .A2(new_n457), .A3(new_n559), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  AND3_X1   g423(.A1(new_n497), .A2(new_n543), .A3(new_n548), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT33), .B1(new_n537), .B2(KEYINPUT102), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n539), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n611), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n536), .A2(new_n538), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n498), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AOI211_X1 g429(.A(G478), .B(G902), .C1(new_n536), .C2(new_n538), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n498), .A2(new_n189), .ZN(new_n617));
  OR3_X1    g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n315), .A3(new_n557), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n435), .A2(new_n189), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G472), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n437), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n607), .A2(new_n371), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT34), .B(G104), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NAND3_X1  g442(.A1(new_n497), .A2(new_n543), .A3(new_n548), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n542), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n315), .A2(new_n557), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n625), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT35), .B(G107), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n358), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n354), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n369), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n367), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n623), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n315), .A2(new_n559), .A3(new_n640), .A4(new_n607), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT37), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n322), .ZN(G12));
  AOI22_X1  g457(.A1(new_n601), .A2(new_n606), .B1(new_n441), .B2(new_n456), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n554), .A2(G900), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n552), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n629), .A2(new_n542), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n644), .A2(new_n315), .A3(new_n638), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT103), .B(G128), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G30));
  XNOR2_X1  g465(.A(new_n646), .B(KEYINPUT105), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT39), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n607), .A2(new_n654), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n542), .B(new_n610), .C1(new_n655), .C2(KEYINPUT40), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n656), .B(new_n187), .C1(KEYINPUT40), .C2(new_n655), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n313), .A2(new_n314), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n658), .B(KEYINPUT38), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n445), .A2(new_n431), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n424), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n661), .A2(KEYINPUT104), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n189), .B1(new_n661), .B2(KEYINPUT104), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n638), .B1(new_n441), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n657), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n260), .ZN(G45));
  NOR3_X1   g483(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n629), .A2(new_n670), .A3(new_n646), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n644), .A2(new_n315), .A3(new_n638), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  AND3_X1   g487(.A1(new_n435), .A2(new_n439), .A3(new_n436), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n439), .B1(new_n435), .B2(new_n436), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n456), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n598), .ZN(new_n677));
  INV_X1    g491(.A(G469), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n603), .B(new_n677), .C1(new_n678), .C2(new_n590), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n676), .A2(new_n680), .A3(new_n371), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n557), .A3(new_n315), .A4(new_n619), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND4_X1  g498(.A1(new_n681), .A2(new_n557), .A3(new_n315), .A4(new_n630), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NAND2_X1  g500(.A1(new_n315), .A2(new_n638), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n559), .A2(new_n676), .A3(new_n680), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT106), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n219), .ZN(G21));
  AOI211_X1 g505(.A(new_n188), .B(new_n679), .C1(new_n313), .C2(new_n314), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n425), .B(new_n434), .C1(new_n446), .C2(new_n422), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n436), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n622), .A2(new_n371), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n622), .A2(new_n371), .A3(KEYINPUT107), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n610), .A2(new_n542), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n692), .A2(new_n699), .A3(new_n557), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  AND3_X1   g516(.A1(new_n622), .A2(new_n638), .A3(new_n694), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n692), .A2(new_n671), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  NAND3_X1  g519(.A1(new_n313), .A2(new_n187), .A3(new_n314), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n629), .A2(new_n670), .A3(new_n646), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n596), .A2(new_n598), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT42), .B1(new_n710), .B2(new_n457), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n457), .A2(KEYINPUT108), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n676), .A2(new_n371), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT42), .A4(new_n710), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n712), .A2(new_n715), .A3(KEYINPUT42), .ZN(new_n719));
  INV_X1    g533(.A(new_n706), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n671), .A3(new_n708), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT109), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n711), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n374), .ZN(G33));
  NOR3_X1   g538(.A1(new_n706), .A2(new_n713), .A3(new_n709), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n648), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n610), .A2(new_n728), .A3(new_n670), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n610), .A2(KEYINPUT110), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n629), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n618), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n729), .B1(new_n733), .B2(new_n728), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n734), .A2(new_n624), .A3(new_n639), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(KEYINPUT44), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n592), .A2(new_n594), .ZN(new_n737));
  XOR2_X1   g551(.A(new_n737), .B(KEYINPUT45), .Z(new_n738));
  OAI21_X1  g552(.A(G469), .B1(new_n738), .B2(G902), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT46), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(G469), .C1(new_n738), .C2(G902), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n603), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n677), .A3(new_n654), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n736), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n706), .B1(new_n735), .B2(KEYINPUT44), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G137), .ZN(G39));
  NAND2_X1  g562(.A1(new_n743), .A2(new_n677), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n743), .A2(KEYINPUT47), .A3(new_n677), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n671), .A3(new_n720), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n441), .A2(new_n456), .A3(new_n372), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n328), .ZN(G42));
  NAND3_X1  g571(.A1(new_n371), .A2(new_n599), .A3(new_n187), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT111), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n759), .A2(new_n441), .A3(new_n664), .ZN(new_n760));
  INV_X1    g574(.A(new_n603), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n590), .A2(new_n678), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT49), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n760), .A2(new_n659), .A3(new_n733), .A4(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n701), .A2(new_n682), .A3(new_n685), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n608), .B(new_n641), .C1(new_n620), .C2(new_n625), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n689), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n631), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n625), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n315), .A2(KEYINPUT112), .A3(new_n557), .A4(new_n630), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n766), .A2(new_n768), .A3(new_n769), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n723), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n725), .A2(new_n648), .B1(new_n710), .B2(new_n703), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n607), .A2(new_n676), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n313), .A2(new_n187), .A3(new_n314), .A4(new_n646), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n549), .A2(new_n639), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT113), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n779), .ZN(new_n783));
  AND4_X1   g597(.A1(KEYINPUT113), .A2(new_n783), .A3(new_n644), .A4(new_n781), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n777), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n704), .A2(new_n649), .A3(new_n672), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n700), .A2(new_n315), .A3(new_n665), .A4(new_n646), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n709), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(KEYINPUT52), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n704), .A2(new_n649), .A3(new_n672), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n791), .B1(new_n792), .B2(new_n788), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n785), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n776), .A2(KEYINPUT53), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT53), .B1(new_n776), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n796), .A2(KEYINPUT114), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n697), .A2(new_n698), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n734), .A2(new_n802), .A3(new_n552), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n188), .A3(new_n659), .A4(new_n680), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(KEYINPUT50), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n804), .B(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n761), .A2(new_n762), .A3(new_n599), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n803), .B(new_n720), .C1(new_n753), .C2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n706), .A2(new_n552), .A3(new_n679), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n441), .A2(new_n371), .A3(new_n664), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n810), .A2(new_n610), .A3(new_n618), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n734), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n703), .A3(new_n810), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n809), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n807), .A2(KEYINPUT51), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT51), .B1(new_n807), .B2(new_n816), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n817), .A2(new_n818), .A3(new_n550), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n803), .A2(new_n692), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n795), .A2(new_n796), .A3(KEYINPUT54), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n801), .A2(new_n819), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n810), .A2(new_n619), .A3(new_n812), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n814), .A2(new_n716), .A3(new_n810), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT48), .Z(new_n826));
  NOR3_X1   g640(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(G952), .A2(G953), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n765), .B1(new_n827), .B2(new_n828), .ZN(G75));
  NOR2_X1   g643(.A1(new_n797), .A2(new_n189), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(G210), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT56), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n303), .A2(new_n305), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n307), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT55), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n833), .A2(new_n837), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n284), .A2(G952), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G51));
  XOR2_X1   g655(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n678), .B2(new_n189), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(G469), .A3(G902), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n776), .A2(new_n794), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n776), .A2(new_n794), .A3(KEYINPUT53), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n844), .B(new_n845), .C1(new_n821), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n602), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n830), .A2(G469), .A3(new_n738), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n840), .B1(new_n855), .B2(new_n856), .ZN(G54));
  NAND3_X1  g671(.A1(new_n830), .A2(KEYINPUT58), .A3(G475), .ZN(new_n858));
  INV_X1    g672(.A(new_n493), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n860), .A2(new_n861), .A3(new_n840), .ZN(G60));
  INV_X1    g676(.A(new_n840), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n612), .A2(new_n614), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n617), .B(KEYINPUT59), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n864), .B(new_n866), .C1(new_n821), .C2(new_n851), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n801), .B2(new_n822), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n863), .B(new_n867), .C1(new_n868), .C2(new_n864), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(G63));
  XNOR2_X1  g684(.A(new_n636), .B(KEYINPUT122), .ZN(new_n871));
  XNOR2_X1  g685(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n363), .A2(new_n189), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(new_n795), .B2(new_n796), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT121), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n874), .C1(new_n795), .C2(new_n796), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n871), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n368), .B(KEYINPUT123), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n878), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n863), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n883), .A2(new_n885), .A3(new_n863), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n883), .B2(new_n863), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n879), .ZN(new_n888));
  XNOR2_X1  g702(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(G66));
  NAND2_X1  g704(.A1(new_n555), .A2(new_n283), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(G953), .ZN(new_n892));
  INV_X1    g706(.A(new_n775), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n892), .B1(new_n893), .B2(G953), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n834), .B1(G898), .B2(new_n284), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n894), .B(new_n895), .ZN(G69));
  NAND2_X1  g710(.A1(new_n405), .A2(new_n411), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n485), .ZN(new_n898));
  NAND2_X1  g712(.A1(G900), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n747), .B1(new_n755), .B2(new_n754), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n716), .A2(new_n315), .A3(new_n700), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n786), .B(new_n726), .C1(new_n901), .C2(new_n744), .ZN(new_n902));
  OR3_X1    g716(.A1(new_n900), .A2(new_n723), .A3(new_n902), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n898), .B(new_n899), .C1(new_n903), .C2(G953), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n786), .B1(new_n667), .B2(new_n657), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n756), .B1(new_n746), .B2(new_n745), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n619), .A2(new_n630), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n655), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n911), .A2(new_n457), .A3(new_n720), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n907), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT127), .A4(new_n913), .ZN(new_n917));
  AOI21_X1  g731(.A(G953), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n898), .B(KEYINPUT125), .Z(new_n919));
  OAI21_X1  g733(.A(new_n904), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n284), .B1(G227), .B2(G900), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G72));
  NAND2_X1  g736(.A1(new_n451), .A2(new_n424), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n916), .A2(new_n917), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n422), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n903), .A2(new_n431), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n893), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(G472), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT63), .Z(new_n929));
  OAI211_X1 g743(.A(new_n929), .B(new_n923), .C1(new_n799), .C2(new_n800), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n923), .A2(new_n929), .ZN(new_n931));
  AND4_X1   g745(.A1(new_n863), .A2(new_n927), .A3(new_n930), .A4(new_n931), .ZN(G57));
endmodule


