//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G902), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  OAI211_X1 g006(.A(G128), .B(new_n189), .C1(new_n190), .C2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(G137), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n196), .A2(new_n198), .A3(new_n199), .A4(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n195), .A2(G137), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n197), .A2(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(G131), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n191), .A2(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n188), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n205), .B(new_n206), .C1(KEYINPUT1), .C2(new_n207), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n193), .A2(new_n201), .A3(new_n204), .A4(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n196), .A2(new_n198), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(G131), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n196), .A2(new_n198), .A3(new_n200), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(G131), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n205), .A2(new_n206), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT0), .B(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n209), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT2), .ZN(new_n221));
  INV_X1    g035(.A(G113), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT64), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(KEYINPUT2), .B2(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT2), .A2(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(G116), .B(G119), .Z(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n223), .A2(new_n225), .B1(KEYINPUT2), .B2(G113), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n220), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n228), .A2(new_n229), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n232), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(KEYINPUT67), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n219), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n237), .ZN(new_n239));
  INV_X1    g053(.A(new_n219), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n241), .B1(new_n239), .B2(new_n240), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n238), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n246));
  NOR2_X1   g060(.A1(G237), .A2(G953), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G210), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n246), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT26), .B(G101), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT29), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n187), .B1(new_n245), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n239), .A2(new_n240), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n209), .A2(KEYINPUT30), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n212), .A2(G131), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n218), .B1(new_n201), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n201), .ZN(new_n261));
  INV_X1    g075(.A(new_n218), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n263), .A2(KEYINPUT65), .A3(KEYINPUT30), .A4(new_n209), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n230), .A2(new_n233), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n219), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n265), .A2(KEYINPUT66), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT66), .B1(new_n265), .B2(new_n268), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n255), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n251), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n219), .B1(new_n233), .B2(new_n230), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n252), .B(new_n273), .C1(new_n243), .C2(new_n244), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n254), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G472), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT71), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n275), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n251), .B2(new_n271), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n280), .B(G472), .C1(new_n282), .C2(new_n254), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n273), .B1(new_n243), .B2(new_n244), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n251), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n252), .A2(new_n255), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n209), .A2(KEYINPUT30), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT65), .B1(new_n289), .B2(new_n263), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n257), .A2(new_n259), .A3(new_n256), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n268), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n265), .A2(KEYINPUT66), .A3(new_n268), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n288), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n287), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n288), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n297), .B(new_n299), .C1(new_n269), .C2(new_n270), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n296), .A2(KEYINPUT69), .A3(new_n297), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n298), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n285), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n299), .B1(new_n269), .B2(new_n270), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n308), .A2(KEYINPUT31), .B1(new_n251), .B2(new_n286), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT69), .B1(new_n296), .B2(new_n297), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n300), .A2(new_n301), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT32), .A3(new_n305), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n284), .A2(new_n307), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G953), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(G221), .A3(G234), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT75), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT22), .B(G137), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT16), .ZN(new_n325));
  OR3_X1    g139(.A1(new_n323), .A2(KEYINPUT16), .A3(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(G146), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n325), .A2(new_n326), .A3(new_n329), .A4(G146), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n191), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n335));
  XNOR2_X1  g149(.A(G119), .B(G128), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(KEYINPUT72), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT24), .B(G110), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(G128), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n343), .B(new_n344), .C1(G119), .C2(new_n207), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G110), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n335), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT72), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n336), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n338), .ZN(new_n350));
  INV_X1    g164(.A(new_n346), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(KEYINPUT73), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n334), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n337), .A2(new_n339), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n325), .A2(new_n326), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n191), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n327), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n345), .A2(G110), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n320), .B1(new_n353), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n328), .A2(new_n330), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n191), .B2(new_n332), .ZN(new_n363));
  INV_X1    g177(.A(new_n352), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT73), .B1(new_n350), .B2(new_n351), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n359), .A3(new_n319), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n368), .B1(new_n187), .B2(G234), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G902), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n361), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n371), .B(KEYINPUT76), .Z(new_n372));
  INV_X1    g186(.A(new_n369), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n361), .A2(new_n367), .A3(new_n187), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n361), .A2(new_n367), .A3(KEYINPUT25), .A4(new_n187), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT3), .B1(new_n380), .B2(G107), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n382));
  INV_X1    g196(.A(G107), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(G104), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(G107), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G101), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT79), .ZN(new_n388));
  INV_X1    g202(.A(G101), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n381), .A2(new_n384), .A3(new_n389), .A4(new_n385), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n390), .A2(KEYINPUT4), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT79), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n392), .A3(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n386), .A2(G101), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n218), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n193), .A2(new_n208), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n380), .A2(G107), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n383), .A2(G104), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n390), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT10), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n193), .A2(new_n390), .A3(new_n402), .A4(new_n208), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT10), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n398), .A2(new_n408), .A3(new_n213), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n315), .A2(G227), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT78), .ZN(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G140), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n213), .B1(new_n398), .B2(new_n408), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n193), .A2(new_n208), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n390), .A2(new_n402), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n213), .B1(new_n421), .B2(new_n406), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n398), .A2(new_n408), .A3(new_n213), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n418), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n406), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n208), .A2(new_n193), .B1(new_n390), .B2(new_n402), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n261), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n423), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n422), .A2(KEYINPUT12), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT80), .A3(new_n409), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n426), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n417), .B1(new_n434), .B2(new_n413), .ZN(new_n435));
  OAI21_X1  g249(.A(G469), .B1(new_n435), .B2(G902), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n415), .A2(new_n424), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n394), .A2(new_n397), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n406), .B(new_n404), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n261), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n414), .B1(new_n441), .B2(new_n409), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n437), .B(new_n187), .C1(new_n438), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT81), .ZN(new_n444));
  INV_X1    g258(.A(new_n187), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n413), .B1(new_n425), .B2(new_n416), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n432), .A2(new_n414), .A3(new_n409), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n437), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n436), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G214), .B1(G237), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G210), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n193), .A2(new_n323), .A3(new_n208), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n215), .B(G125), .C1(new_n216), .C2(new_n217), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G224), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G953), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n459), .B(new_n461), .Z(new_n462));
  INV_X1    g276(.A(KEYINPUT5), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n342), .A3(G116), .ZN(new_n464));
  OAI211_X1 g278(.A(G113), .B(new_n464), .C1(new_n229), .C2(new_n463), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n403), .A2(new_n236), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G110), .B(G122), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n388), .A2(new_n391), .A3(new_n393), .ZN(new_n468));
  OAI22_X1  g282(.A1(new_n230), .A2(new_n233), .B1(KEYINPUT4), .B2(new_n387), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n467), .B(KEYINPUT82), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n470), .A2(KEYINPUT6), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n472), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G902), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n465), .A2(new_n236), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n420), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(KEYINPUT83), .A3(new_n466), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n467), .B(KEYINPUT8), .Z(new_n481));
  AOI22_X1  g295(.A1(new_n465), .A2(new_n236), .B1(new_n390), .B2(new_n402), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n457), .B(new_n458), .C1(new_n486), .C2(new_n461), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n461), .B1(new_n457), .B2(new_n458), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n487), .A2(new_n488), .B1(new_n489), .B2(KEYINPUT7), .ZN(new_n490));
  INV_X1    g304(.A(new_n487), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT84), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n485), .A2(new_n490), .A3(new_n492), .A4(KEYINPUT85), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n470), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n480), .A2(new_n484), .B1(new_n491), .B2(KEYINPUT84), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT85), .B1(new_n495), .B2(new_n490), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n456), .B1(new_n477), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n490), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n470), .A3(new_n493), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n502), .A2(new_n476), .A3(new_n455), .A4(new_n475), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n454), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT9), .B(G234), .ZN(new_n505));
  OAI21_X1  g319(.A(G221), .B1(new_n505), .B2(G902), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT77), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n452), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(G104), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT88), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n188), .A2(KEYINPUT86), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(G214), .A3(new_n247), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n247), .A2(G214), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT86), .B(G143), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n322), .A2(new_n324), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G146), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n333), .ZN(new_n522));
  INV_X1    g336(.A(new_n515), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT86), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G143), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n525), .A2(new_n514), .B1(new_n247), .B2(G214), .ZN(new_n526));
  OAI21_X1  g340(.A(G131), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n519), .B(new_n522), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n199), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n356), .B(new_n327), .C1(new_n527), .C2(new_n530), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n513), .B(new_n529), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n476), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n525), .A2(new_n514), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n247), .A2(G214), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n199), .B1(new_n539), .B2(new_n515), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT17), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n532), .A2(new_n541), .A3(new_n356), .A4(new_n327), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n513), .B1(new_n542), .B2(new_n529), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT89), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n512), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT89), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n476), .A4(new_n535), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n544), .A2(G475), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT87), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT19), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n520), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n332), .A2(KEYINPUT19), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n527), .A2(new_n531), .B1(new_n554), .B2(new_n191), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n540), .A2(KEYINPUT18), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n522), .A2(new_n519), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n331), .A2(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n511), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n550), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n531), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n552), .A2(new_n553), .ZN(new_n562));
  OAI22_X1  g376(.A1(new_n561), .A2(new_n540), .B1(new_n562), .B2(G146), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n529), .B1(new_n563), .B2(new_n362), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(KEYINPUT87), .A3(new_n511), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n542), .A2(new_n559), .A3(new_n529), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(G475), .A2(G902), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT20), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT20), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n567), .A2(new_n571), .A3(new_n568), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n549), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G478), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n505), .A2(new_n368), .A3(G953), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT91), .B1(new_n207), .B2(G143), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT91), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(new_n188), .A3(G128), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n579), .A2(new_n581), .A3(KEYINPUT13), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n207), .A2(G143), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G134), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT90), .ZN(new_n589));
  INV_X1    g403(.A(G116), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n589), .B1(new_n590), .B2(G122), .ZN(new_n591));
  INV_X1    g405(.A(G122), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(KEYINPUT90), .A3(G116), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n590), .A2(G122), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G107), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n591), .A2(new_n593), .B1(new_n590), .B2(G122), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n383), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n582), .A2(new_n195), .A3(new_n586), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n588), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n383), .B1(new_n594), .B2(new_n595), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n594), .A2(KEYINPUT14), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n598), .B1(KEYINPUT14), .B2(new_n383), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n582), .A2(new_n195), .A3(new_n586), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n195), .B1(new_n582), .B2(new_n586), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n606), .B(new_n607), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n602), .A2(new_n603), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n603), .B1(new_n602), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n578), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n582), .A2(new_n583), .B1(new_n207), .B2(G143), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n195), .B1(new_n614), .B2(new_n585), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n594), .A2(new_n383), .A3(new_n595), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n601), .B1(new_n616), .B2(new_n604), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n604), .A2(new_n605), .ZN(new_n619));
  OAI22_X1  g433(.A1(new_n615), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT92), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n602), .A2(new_n603), .A3(new_n610), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n577), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n576), .B1(new_n624), .B2(new_n187), .ZN(new_n625));
  AOI211_X1 g439(.A(new_n445), .B(new_n575), .C1(new_n613), .C2(new_n623), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(G952), .ZN(new_n628));
  AOI211_X1 g442(.A(G953), .B(new_n628), .C1(G234), .C2(G237), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n315), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT21), .B(G898), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n573), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n314), .A2(new_n379), .A3(new_n509), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT93), .B(G101), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G3));
  NAND2_X1  g451(.A1(new_n504), .A2(new_n633), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n611), .A2(new_n612), .A3(new_n578), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n577), .B1(new_n621), .B2(new_n622), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n613), .A2(KEYINPUT33), .A3(new_n623), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n445), .A2(new_n574), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n187), .B1(new_n640), .B2(new_n641), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n574), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n544), .A2(G475), .A3(new_n548), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n567), .A2(new_n571), .A3(new_n568), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n571), .B1(new_n567), .B2(new_n568), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n638), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n507), .B1(new_n436), .B2(new_n451), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n655), .A2(new_n379), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n312), .A2(new_n187), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n657), .A2(G472), .B1(new_n305), .B2(new_n312), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n654), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  OR2_X1    g475(.A1(new_n625), .A2(new_n626), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n573), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n638), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n656), .A3(new_n658), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NAND2_X1  g481(.A1(new_n376), .A2(new_n377), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n369), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n366), .A2(new_n359), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n320), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n370), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n509), .A2(new_n658), .A3(new_n634), .A4(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  AND3_X1   g491(.A1(new_n655), .A2(new_n504), .A3(new_n674), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n630), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n629), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n663), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n678), .A2(new_n314), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(KEYINPUT94), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT94), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n678), .A2(new_n314), .A3(new_n687), .A4(new_n684), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XNOR2_X1  g504(.A(new_n682), .B(KEYINPUT39), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n655), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT40), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n252), .B1(new_n238), .B2(new_n255), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n476), .B1(new_n296), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G472), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n313), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n307), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n498), .A2(new_n503), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT38), .Z(new_n700));
  NOR2_X1   g514(.A1(new_n573), .A2(new_n627), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n453), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n700), .A2(new_n674), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n693), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  NOR2_X1   g519(.A1(new_n653), .A2(new_n683), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n678), .A2(new_n314), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  OR2_X1    g522(.A1(new_n448), .A2(new_n437), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n446), .A2(new_n447), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n449), .A2(new_n710), .A3(new_n437), .A4(new_n187), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n449), .B1(new_n448), .B2(new_n437), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n508), .B(new_n709), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT95), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT95), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n451), .A2(new_n715), .A3(new_n508), .A4(new_n709), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n314), .A3(new_n654), .A4(new_n379), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND4_X1  g534(.A1(new_n717), .A2(new_n314), .A3(new_n664), .A4(new_n379), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  AND2_X1   g536(.A1(new_n634), .A2(new_n674), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n314), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n714), .A2(new_n504), .A3(new_n716), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT96), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n714), .A2(KEYINPUT96), .A3(new_n504), .A4(new_n716), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT97), .B(G119), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G21));
  AOI211_X1 g545(.A(new_n454), .B(new_n632), .C1(new_n498), .C2(new_n503), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n714), .A3(new_n701), .A4(new_n716), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n303), .A2(new_n302), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n308), .A2(KEYINPUT31), .B1(new_n251), .B2(new_n245), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n306), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n304), .A2(new_n445), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT98), .B(G472), .Z(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n737), .B(new_n379), .C1(new_n738), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n733), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n592), .ZN(G24));
  NAND2_X1  g557(.A1(new_n727), .A2(new_n728), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n740), .B1(new_n312), .B2(new_n187), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n736), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n674), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n744), .A2(new_n706), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NOR2_X1   g564(.A1(new_n711), .A2(new_n712), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n432), .A2(KEYINPUT80), .A3(new_n409), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT80), .B1(new_n432), .B2(new_n409), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n413), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n417), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n437), .B1(new_n756), .B2(new_n476), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT99), .B1(new_n751), .B2(new_n757), .ZN(new_n758));
  AND4_X1   g572(.A1(KEYINPUT42), .A2(new_n648), .A3(new_n652), .A4(new_n682), .ZN(new_n759));
  AND4_X1   g573(.A1(new_n508), .A2(new_n498), .A3(new_n453), .A4(new_n503), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT99), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n436), .A2(new_n451), .A3(new_n761), .ZN(new_n762));
  AND4_X1   g576(.A1(new_n758), .A2(new_n759), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT100), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n313), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n312), .A2(KEYINPUT100), .A3(KEYINPUT32), .A4(new_n305), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n307), .A3(new_n284), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n767), .A3(new_n379), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT101), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n763), .A2(new_n767), .A3(KEYINPUT101), .A4(new_n379), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n314), .A2(new_n379), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n758), .A2(new_n760), .A3(new_n762), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n706), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT102), .B(G131), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G33));
  NAND4_X1  g594(.A1(new_n773), .A2(KEYINPUT103), .A3(new_n684), .A4(new_n774), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n774), .A2(new_n314), .A3(new_n379), .A4(new_n684), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT103), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  NAND2_X1  g600(.A1(new_n435), .A2(KEYINPUT45), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT104), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n437), .B1(new_n756), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(G469), .A2(G902), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n451), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n508), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n691), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n699), .A2(new_n454), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n648), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n652), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT43), .ZN(new_n806));
  INV_X1    g620(.A(new_n658), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n807), .A3(new_n674), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n803), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n801), .B(new_n810), .C1(new_n809), .C2(new_n808), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  NAND2_X1  g626(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n799), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n815));
  INV_X1    g629(.A(new_n813), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n798), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n314), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n371), .B(KEYINPUT76), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n669), .A2(new_n819), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n818), .A2(new_n820), .A3(new_n706), .A4(new_n802), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n814), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  NAND4_X1  g637(.A1(new_n805), .A2(new_n379), .A3(new_n508), .A4(new_n453), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n451), .A2(new_n709), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(KEYINPUT49), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n825), .A2(KEYINPUT49), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n698), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n700), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n806), .A2(new_n629), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n745), .A2(new_n820), .A3(new_n736), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n700), .A2(new_n454), .A3(new_n717), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n717), .A2(new_n802), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n837), .A2(new_n838), .B1(new_n748), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n836), .A2(KEYINPUT113), .A3(new_n842), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n379), .A2(new_n839), .A3(new_n629), .A4(new_n829), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n573), .A3(new_n804), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n841), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT114), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n814), .A2(new_n817), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n508), .B2(new_n825), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n834), .A2(new_n803), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT112), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n831), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n653), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n628), .B(G953), .C1(new_n844), .C2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n767), .A2(new_n379), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n840), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g672(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n840), .A2(KEYINPUT115), .A3(KEYINPUT48), .A4(new_n857), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n832), .A2(new_n744), .A3(new_n833), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n856), .A2(new_n860), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n846), .A2(new_n831), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n864), .B2(new_n852), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n854), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n504), .A2(new_n701), .A3(new_n633), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n833), .A2(new_n717), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n718), .A2(new_n869), .A3(new_n665), .A4(new_n675), .ZN(new_n870));
  INV_X1    g684(.A(new_n721), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n870), .A2(new_n729), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT106), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n635), .B2(new_n659), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n635), .A2(new_n659), .A3(new_n873), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n746), .A2(new_n674), .A3(new_n706), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n758), .A2(new_n760), .A3(new_n762), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n683), .B1(new_n669), .B2(new_n673), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n662), .A2(new_n652), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n802), .A2(new_n655), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n878), .A2(new_n879), .B1(new_n818), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n781), .B2(new_n784), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n778), .A2(new_n872), .A3(new_n877), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT107), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n635), .A2(new_n659), .A3(new_n873), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n874), .ZN(new_n888));
  OAI21_X1  g702(.A(G472), .B1(new_n304), .B2(new_n445), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n312), .A2(new_n305), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n655), .A3(new_n379), .A4(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n732), .A2(new_n662), .A3(new_n573), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n890), .A3(new_n674), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n655), .A2(new_n634), .A3(new_n504), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n891), .A2(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n742), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n314), .A2(new_n723), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n744), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(new_n898), .A3(new_n718), .A4(new_n721), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT107), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n778), .A4(new_n884), .ZN(new_n902));
  INV_X1    g716(.A(new_n707), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n686), .B2(new_n688), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n758), .A2(new_n762), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n702), .B1(new_n498), .B2(new_n503), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n507), .B1(new_n682), .B2(KEYINPUT108), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(KEYINPUT108), .B2(new_n682), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n674), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n698), .A2(new_n905), .A3(new_n906), .A4(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n904), .A2(new_n749), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT52), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n904), .A2(KEYINPUT52), .A3(new_n749), .A4(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n886), .A2(new_n902), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT53), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n886), .A2(new_n902), .A3(new_n915), .ZN(new_n919));
  XOR2_X1   g733(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI22_X1  g735(.A1(new_n918), .A2(KEYINPUT109), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n885), .A2(KEYINPUT107), .B1(new_n913), .B2(new_n914), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT53), .B1(new_n923), .B2(new_n902), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT109), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n867), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n916), .A2(new_n920), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n885), .A2(new_n917), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n915), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n867), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT111), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  OAI22_X1  g747(.A1(new_n924), .A2(new_n925), .B1(new_n916), .B2(new_n920), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n918), .A2(KEYINPUT109), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT54), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT111), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n937), .A3(new_n931), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n866), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(G952), .A2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n830), .B1(new_n939), .B2(new_n940), .ZN(G75));
  AOI21_X1  g755(.A(new_n921), .B1(new_n923), .B2(new_n902), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n929), .A2(new_n915), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n187), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n456), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n473), .A2(new_n474), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n462), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT55), .ZN(new_n949));
  NOR2_X1   g763(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n950));
  AND2_X1   g764(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n946), .B(new_n949), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n315), .A2(G952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT56), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n949), .B1(new_n946), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT116), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(G51));
  OAI21_X1  g775(.A(KEYINPUT54), .B1(new_n942), .B2(new_n943), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT118), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n931), .A3(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(KEYINPUT118), .B(KEYINPUT54), .C1(new_n942), .C2(new_n943), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n792), .B(KEYINPUT57), .Z(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT119), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n964), .A2(KEYINPUT119), .A3(new_n965), .A4(new_n966), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n710), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n945), .A2(new_n788), .A3(new_n790), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n953), .B1(new_n971), .B2(new_n972), .ZN(G54));
  NAND3_X1  g787(.A1(new_n945), .A2(KEYINPUT58), .A3(G475), .ZN(new_n974));
  INV_X1    g788(.A(new_n567), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n953), .ZN(G60));
  NAND2_X1  g792(.A1(new_n642), .A2(new_n643), .ZN(new_n979));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT59), .Z(new_n981));
  NOR2_X1   g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n964), .A2(new_n965), .A3(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n983), .A2(KEYINPUT120), .A3(new_n954), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT120), .B1(new_n983), .B2(new_n954), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n981), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n933), .A2(new_n938), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n979), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n986), .A2(new_n989), .ZN(G63));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT60), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n944), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n361), .A2(new_n367), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n954), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n672), .B2(new_n993), .ZN(new_n996));
  XNOR2_X1  g810(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G66));
  INV_X1    g812(.A(KEYINPUT122), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n631), .A2(new_n460), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n900), .A2(G953), .ZN(new_n1002));
  MUX2_X1   g816(.A(new_n1001), .B(new_n999), .S(new_n1002), .Z(new_n1003));
  OAI21_X1  g817(.A(new_n947), .B1(G898), .B2(new_n315), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1003), .B(new_n1004), .Z(G69));
  OAI21_X1  g819(.A(new_n265), .B1(KEYINPUT30), .B2(new_n240), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(new_n562), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G900), .A2(G953), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n857), .A2(new_n906), .ZN(new_n1009));
  OR3_X1    g823(.A1(new_n800), .A2(KEYINPUT124), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(KEYINPUT124), .B1(new_n800), .B2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n904), .A2(new_n749), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1013), .A2(new_n778), .A3(new_n785), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1012), .A2(new_n811), .A3(new_n822), .A4(new_n1014), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1007), .B(new_n1008), .C1(new_n1015), .C2(G953), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT123), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n803), .B1(new_n653), .B2(new_n663), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n773), .A2(new_n692), .A3(new_n1018), .ZN(new_n1019));
  AND3_X1   g833(.A1(new_n811), .A2(new_n822), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1013), .A2(new_n704), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(KEYINPUT62), .ZN(new_n1022));
  OR2_X1    g836(.A1(new_n1021), .A2(KEYINPUT62), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1024), .A2(new_n315), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n1016), .B(new_n1017), .C1(new_n1025), .C2(new_n1007), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1016), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1007), .B1(new_n1024), .B2(new_n315), .ZN(new_n1028));
  OAI21_X1  g842(.A(KEYINPUT123), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n315), .B1(G227), .B2(G900), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1030), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1031), .A2(new_n1032), .ZN(G72));
  NAND2_X1  g847(.A1(G472), .A2(G902), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT63), .Z(new_n1035));
  INV_X1    g849(.A(new_n900), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1035), .B1(new_n1015), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n271), .B(KEYINPUT125), .Z(new_n1038));
  NOR2_X1   g852(.A1(new_n1038), .A2(new_n252), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n953), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1038), .A2(new_n252), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n1020), .A2(new_n900), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1041), .B1(new_n1042), .B2(new_n1035), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT126), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g859(.A(KEYINPUT126), .B(new_n1041), .C1(new_n1042), .C2(new_n1035), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1040), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n922), .A2(new_n926), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1035), .ZN(new_n1049));
  OR2_X1    g863(.A1(new_n272), .A2(KEYINPUT127), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n296), .B1(new_n272), .B2(KEYINPUT127), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1047), .B1(new_n1048), .B2(new_n1052), .ZN(G57));
endmodule


