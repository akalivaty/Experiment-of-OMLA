//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  NOR3_X1   g0009(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n210), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT64), .B(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G50), .A2(G226), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n212), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n215), .B1(new_n211), .B2(new_n214), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G226), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(G232), .Z(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND2_X1  g0041(.A1(G33), .A2(G41), .ZN(new_n242));
  NAND3_X1  g0042(.A1(new_n242), .A2(G1), .A3(G13), .ZN(new_n243));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  OAI21_X1  g0044(.A(new_n244), .B1(G41), .B2(G45), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n243), .A2(G238), .A3(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G41), .ZN(new_n247));
  INV_X1    g0047(.A(G45), .ZN(new_n248));
  AOI21_X1  g0048(.A(G1), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G274), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(G226), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  OAI211_X1 g0055(.A(G232), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n243), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n251), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT13), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT72), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n258), .A2(new_n259), .ZN(new_n264));
  INV_X1    g0064(.A(new_n251), .ZN(new_n265));
  AND4_X1   g0065(.A1(new_n263), .A2(new_n264), .A3(new_n261), .A4(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n260), .B2(new_n261), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G200), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n270), .A2(KEYINPUT65), .A3(new_n209), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT65), .B1(new_n270), .B2(new_n209), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G68), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n275), .A2(G50), .B1(G20), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G77), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n208), .A2(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT11), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n270), .A2(new_n209), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n244), .A2(G13), .A3(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n287), .A2(new_n244), .A3(G13), .A4(G20), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n284), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n244), .A2(G20), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G68), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n286), .A2(new_n276), .A3(new_n288), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT12), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n274), .A2(KEYINPUT11), .A3(new_n280), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n283), .A2(new_n292), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n260), .A2(new_n261), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n264), .A2(new_n261), .A3(new_n265), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n269), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n262), .A2(G179), .A3(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT73), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT73), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n262), .A2(new_n306), .A3(G179), .A4(new_n300), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n260), .A2(new_n263), .A3(new_n261), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n297), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT14), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT14), .B1(new_n268), .B2(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n308), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT74), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n296), .B(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n303), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT75), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n312), .B1(new_n311), .B2(new_n313), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n268), .A2(KEYINPUT14), .A3(G169), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n322), .A2(new_n323), .B1(new_n307), .B2(new_n305), .ZN(new_n324));
  INV_X1    g0124(.A(new_n318), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT75), .B1(new_n326), .B2(new_n303), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n259), .A2(new_n249), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G226), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n250), .ZN(new_n330));
  OR2_X1    g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G223), .A3(G1698), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(G222), .A3(new_n252), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n334), .B(new_n335), .C1(new_n216), .C2(new_n333), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n330), .B1(new_n336), .B2(new_n259), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G179), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n313), .B2(new_n337), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n275), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT66), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G58), .ZN(new_n344));
  OR3_X1    g0144(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT8), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n340), .B1(new_n346), .B2(new_n279), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n274), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n286), .A2(new_n288), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n273), .A2(G50), .A3(new_n290), .A4(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT68), .ZN(new_n351));
  INV_X1    g0151(.A(new_n349), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n202), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n350), .B2(new_n353), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n348), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n339), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n336), .A2(new_n259), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n358), .A2(G190), .A3(new_n250), .A4(new_n329), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n337), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT9), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(new_n356), .ZN(new_n363));
  OAI211_X1 g0163(.A(KEYINPUT9), .B(new_n348), .C1(new_n354), .C2(new_n355), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT71), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n364), .A2(new_n365), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT10), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT10), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(new_n363), .C1(new_n366), .C2(new_n367), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n357), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n373));
  OAI211_X1 g0173(.A(G223), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n374));
  OAI211_X1 g0174(.A(G226), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n259), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n243), .A2(G232), .A3(new_n245), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n250), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(G190), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT76), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n380), .B1(new_n377), .B2(new_n259), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT76), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n383), .B1(new_n388), .B2(new_n360), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n343), .A2(new_n345), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n290), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n273), .A2(new_n349), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n391), .A2(new_n392), .B1(new_n349), .B2(new_n390), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n333), .B2(G20), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n253), .A2(new_n254), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n276), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n344), .A2(new_n276), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n201), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n275), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n395), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n398), .B2(new_n208), .ZN(new_n406));
  NOR4_X1   g0206(.A1(new_n253), .A2(new_n254), .A3(new_n396), .A4(G20), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n404), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(KEYINPUT16), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n284), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n394), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n373), .B1(new_n389), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g0213(.A(new_n384), .B(new_n380), .C1(new_n259), .C2(new_n377), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT76), .B1(new_n378), .B2(new_n381), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n313), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n382), .A2(G179), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n284), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n408), .A2(new_n409), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n395), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n393), .B1(new_n422), .B2(new_n410), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT18), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n360), .B1(new_n414), .B2(new_n415), .ZN(new_n425));
  INV_X1    g0225(.A(new_n383), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(KEYINPUT77), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n423), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n412), .A2(new_n431), .A3(new_n416), .A4(new_n418), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n413), .A2(new_n424), .A3(new_n430), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n333), .A2(G238), .A3(G1698), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n333), .A2(G232), .A3(new_n252), .ZN(new_n435));
  INV_X1    g0235(.A(G107), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n434), .B(new_n435), .C1(new_n436), .C2(new_n333), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n259), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n328), .A2(G244), .B1(G274), .B2(new_n249), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n298), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(G200), .B2(new_n440), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n291), .A2(G77), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT15), .B(G87), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n208), .A2(new_n216), .B1(new_n444), .B2(new_n279), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n341), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n284), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n216), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n443), .B(new_n449), .C1(new_n450), .C2(new_n349), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT70), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n451), .A2(KEYINPUT70), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n442), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n440), .A2(G169), .ZN(new_n456));
  INV_X1    g0256(.A(G179), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(new_n440), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n451), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n433), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  AND4_X1   g0261(.A1(new_n321), .A2(new_n327), .A3(new_n372), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n248), .A2(G1), .ZN(new_n464));
  AND2_X1   g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n243), .ZN(new_n468));
  INV_X1    g0268(.A(G270), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT82), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G274), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT82), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n467), .A2(new_n473), .A3(G270), .A4(new_n243), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G264), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n476));
  OAI211_X1 g0276(.A(G257), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n331), .A2(G303), .A3(new_n332), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT83), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n479), .A2(new_n480), .A3(new_n259), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n479), .B2(new_n259), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n470), .B(new_n475), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n286), .A2(new_n484), .A3(new_n288), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT84), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT84), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n286), .A2(new_n487), .A3(new_n484), .A4(new_n288), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n484), .B1(new_n244), .B2(G33), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n486), .A2(new_n488), .B1(new_n289), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G33), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G97), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  AOI21_X1  g0293(.A(G20), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n208), .A2(new_n484), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n284), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT20), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(KEYINPUT20), .B(new_n284), .C1(new_n494), .C2(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n313), .B1(new_n490), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n483), .A2(new_n501), .A3(KEYINPUT21), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT85), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n483), .A2(new_n501), .A3(KEYINPUT85), .A4(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n490), .A2(new_n500), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n483), .A2(new_n457), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n483), .A2(new_n501), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT21), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n483), .A2(G190), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n479), .A2(new_n259), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT83), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n479), .A2(new_n480), .A3(new_n259), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n470), .A2(new_n474), .A3(new_n472), .ZN(new_n517));
  AOI21_X1  g0317(.A(G200), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n500), .B(new_n490), .C1(new_n512), .C2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n506), .A2(new_n511), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G257), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n472), .B1(new_n521), .B2(new_n468), .ZN(new_n522));
  OAI21_X1  g0322(.A(G244), .B1(new_n253), .B2(new_n254), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n523), .A2(new_n524), .B1(G33), .B2(G283), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(G1698), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(G244), .C1(new_n254), .C2(new_n253), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n333), .B2(G250), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n525), .B(new_n527), .C1(new_n252), .C2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n522), .B1(new_n529), .B2(new_n259), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G179), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n217), .B1(new_n331), .B2(new_n332), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n527), .B(new_n493), .C1(new_n532), .C2(KEYINPUT4), .ZN(new_n533));
  OAI21_X1  g0333(.A(G250), .B1(new_n253), .B2(new_n254), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n252), .B1(new_n534), .B2(KEYINPUT4), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n259), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n467), .A2(new_n243), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(G257), .B1(G274), .B2(new_n471), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n313), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  XNOR2_X1  g0340(.A(G97), .B(G107), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT78), .ZN(new_n542));
  OR3_X1    g0342(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT6), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(KEYINPUT6), .ZN(new_n544));
  INV_X1    g0344(.A(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT6), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n543), .A2(G20), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n397), .A2(new_n399), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G107), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n275), .A2(G77), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n284), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n352), .A2(new_n545), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n244), .A2(G33), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n273), .A2(new_n349), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n555), .B2(new_n545), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n531), .A2(new_n540), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT79), .B1(new_n530), .B2(new_n360), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n536), .A2(new_n538), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT79), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(G200), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n536), .A2(G190), .A3(new_n538), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n552), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n558), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(G250), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n568));
  OAI211_X1 g0368(.A(G257), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G294), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n259), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n467), .A2(G264), .A3(new_n243), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT87), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT87), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n467), .A2(new_n575), .A3(G264), .A4(new_n243), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n572), .A2(new_n574), .A3(new_n472), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n360), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n572), .A2(new_n298), .A3(new_n472), .A4(new_n573), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n208), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT22), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT22), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n333), .A2(new_n583), .A3(new_n208), .A4(G87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT86), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(KEYINPUT86), .B(KEYINPUT23), .C1(new_n208), .C2(G107), .ZN(new_n589));
  OR3_X1    g0389(.A1(new_n208), .A2(KEYINPUT23), .A3(G107), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n588), .A2(new_n589), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n585), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n585), .A2(new_n593), .A3(KEYINPUT24), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n284), .A3(new_n597), .ZN(new_n598));
  OR3_X1    g0398(.A1(new_n349), .A2(KEYINPUT25), .A3(G107), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n273), .A2(G107), .A3(new_n349), .A4(new_n554), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT25), .B1(new_n349), .B2(G107), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n580), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n597), .A2(new_n284), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n592), .B1(new_n582), .B2(new_n584), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(KEYINPUT24), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n602), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n572), .A2(new_n472), .A3(new_n573), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n608), .A2(new_n313), .B1(new_n577), .B2(new_n457), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n333), .A2(new_n208), .A3(G68), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT19), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n257), .B2(G20), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n208), .B1(new_n257), .B2(new_n614), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT81), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(KEYINPUT81), .B(new_n208), .C1(new_n257), .C2(new_n614), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n284), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n352), .A2(new_n444), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n273), .A2(G87), .A3(new_n349), .A4(new_n554), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(G244), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n627));
  OAI211_X1 g0427(.A(G238), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n628));
  NAND2_X1  g0428(.A1(G33), .A2(G116), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT80), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT80), .A4(new_n629), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n259), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n464), .A2(G274), .ZN(new_n635));
  INV_X1    g0435(.A(G250), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n464), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n243), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n634), .A2(G190), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n633), .A2(new_n259), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n640), .A2(new_n632), .B1(new_n243), .B2(new_n637), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n626), .B(new_n639), .C1(new_n360), .C2(new_n641), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n623), .B(new_n624), .C1(new_n444), .C2(new_n555), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n634), .A2(new_n457), .A3(new_n638), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n643), .B(new_n644), .C1(new_n641), .C2(G169), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n567), .A2(new_n612), .A3(new_n647), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n463), .A2(new_n520), .A3(new_n648), .ZN(G372));
  NAND2_X1  g0449(.A1(new_n424), .A2(new_n432), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n326), .B1(new_n302), .B2(new_n460), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n413), .A2(new_n430), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n369), .A2(new_n371), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n357), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n560), .A2(new_n457), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n548), .A2(G107), .B1(G77), .B2(new_n275), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n420), .B1(new_n658), .B2(new_n547), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n657), .A2(new_n539), .B1(new_n659), .B2(new_n556), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT26), .B1(new_n646), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n558), .A2(new_n645), .A3(new_n642), .A4(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n661), .A2(new_n645), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n506), .A2(new_n511), .A3(new_n610), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n665), .A2(new_n647), .A3(new_n567), .A4(new_n603), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n656), .B1(new_n463), .B2(new_n668), .ZN(G369));
  AND2_X1   g0469(.A1(new_n506), .A2(new_n511), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n244), .A2(new_n208), .A3(G13), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT88), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n670), .A2(new_n507), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n507), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n520), .A2(new_n679), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n678), .A2(G330), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n607), .A2(new_n609), .A3(new_n677), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT89), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT89), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n607), .A2(new_n677), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n683), .B(new_n684), .C1(new_n611), .C2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n670), .A2(new_n677), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n688), .A2(new_n686), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n610), .A2(new_n677), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n687), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n213), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR4_X1   g0495(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n207), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n677), .B1(new_n664), .B2(new_n666), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI211_X1 g0502(.A(KEYINPUT29), .B(new_n677), .C1(new_n664), .C2(new_n666), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g0504(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n634), .A2(new_n638), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n572), .A2(new_n574), .A3(new_n576), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n707), .A2(new_n560), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT91), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(KEYINPUT30), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(new_n508), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n708), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n641), .A2(new_n530), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n516), .A2(new_n517), .A3(G179), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n483), .A2(new_n707), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n560), .A2(new_n457), .A3(new_n577), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n677), .B(new_n706), .C1(new_n718), .C2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n677), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n713), .A2(new_n717), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT92), .B1(new_n719), .B2(new_n720), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n560), .A2(new_n457), .A3(new_n577), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n516), .A2(new_n517), .B1(new_n634), .B2(new_n638), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT92), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n723), .B1(new_n724), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n722), .B1(new_n731), .B2(KEYINPUT31), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n648), .A2(new_n520), .A3(new_n677), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n704), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n699), .B1(new_n737), .B2(G1), .ZN(G364));
  AND2_X1   g0538(.A1(new_n208), .A2(G13), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G45), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n695), .A2(G1), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n681), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n678), .A2(new_n680), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n743), .B1(G330), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n741), .B(KEYINPUT93), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n693), .A2(new_n398), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n748), .A2(G355), .B1(new_n484), .B2(new_n693), .ZN(new_n749));
  INV_X1    g0549(.A(new_n207), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G45), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n237), .B2(G45), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n693), .A2(new_n333), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n749), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n209), .B1(G20), .B2(new_n313), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n747), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n759), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n208), .A2(G190), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n457), .A3(G200), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT95), .Z(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n436), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n208), .A2(new_n298), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n457), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n457), .A2(new_n360), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n763), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G58), .A2(new_n772), .B1(new_n775), .B2(G68), .ZN(new_n776));
  INV_X1    g0576(.A(new_n769), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n777), .A2(new_n360), .A3(G179), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n763), .A2(new_n770), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n778), .A2(G87), .B1(new_n450), .B2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n298), .A2(G179), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n208), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n545), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n773), .A2(new_n769), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n398), .B(new_n784), .C1(G50), .C2(new_n786), .ZN(new_n787));
  AND4_X1   g0587(.A1(new_n768), .A2(new_n776), .A3(new_n781), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n763), .A2(new_n457), .A3(new_n360), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT94), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  INV_X1    g0596(.A(new_n778), .ZN(new_n797));
  INV_X1    g0597(.A(G303), .ZN(new_n798));
  INV_X1    g0598(.A(G322), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n797), .A2(new_n798), .B1(new_n771), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G326), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n785), .A2(new_n801), .B1(new_n779), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT33), .B(G317), .Z(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n398), .B1(new_n804), .B2(new_n774), .C1(new_n805), .C2(new_n783), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n800), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n793), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n808), .A2(G329), .B1(new_n765), .B2(G283), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n788), .A2(new_n796), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n758), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n761), .B1(new_n762), .B2(new_n810), .C1(new_n744), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n745), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT96), .Z(G396));
  NOR2_X1   g0614(.A1(new_n759), .A2(new_n756), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT97), .Z(new_n816));
  OAI21_X1  g0616(.A(new_n746), .B1(G77), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n771), .A2(new_n805), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n785), .A2(new_n798), .B1(new_n779), .B2(new_n484), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(G107), .C2(new_n778), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n333), .B(new_n784), .C1(G283), .C2(new_n775), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n808), .A2(G311), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n765), .A2(G87), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n786), .A2(G137), .B1(new_n780), .B2(G159), .ZN(new_n825));
  INV_X1    g0625(.A(G143), .ZN(new_n826));
  INV_X1    g0626(.A(G150), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n771), .C1(new_n827), .C2(new_n774), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT34), .Z(new_n829));
  OAI21_X1  g0629(.A(new_n333), .B1(new_n797), .B2(new_n202), .ZN(new_n830));
  INV_X1    g0630(.A(new_n783), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(G58), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n765), .A2(G68), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n793), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n824), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n817), .B1(new_n836), .B2(new_n759), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n460), .A2(new_n723), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n677), .A2(new_n451), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n454), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n839), .B1(new_n459), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n837), .B1(new_n842), .B2(new_n757), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n700), .A2(new_n842), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n700), .A2(new_n842), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n735), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n742), .B1(new_n846), .B2(new_n847), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(KEYINPUT98), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n849), .A2(KEYINPUT98), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n843), .B1(new_n851), .B2(new_n852), .ZN(G384));
  NAND3_X1  g0653(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(KEYINPUT35), .ZN(new_n856));
  NOR4_X1   g0656(.A1(new_n856), .A2(new_n208), .A3(new_n484), .A4(new_n209), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT99), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n857), .A2(new_n858), .B1(KEYINPUT35), .B2(new_n855), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT36), .Z(new_n861));
  OR3_X1    g0661(.A1(new_n207), .A2(new_n216), .A3(new_n401), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n276), .A2(G50), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT100), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n244), .B(G13), .C1(new_n862), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n405), .A2(new_n274), .A3(new_n410), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n675), .B1(new_n394), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n433), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n427), .A2(new_n423), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  INV_X1    g0671(.A(new_n675), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n416), .B2(new_n418), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n870), .B(new_n871), .C1(new_n423), .C2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(G169), .B1(new_n385), .B2(new_n387), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n675), .B1(new_n875), .B2(new_n417), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n394), .A2(new_n867), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n876), .A2(new_n877), .B1(new_n423), .B2(new_n427), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n874), .B1(new_n878), .B2(new_n871), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n869), .B2(new_n879), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT102), .B(KEYINPUT39), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n869), .A2(new_n879), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT39), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n870), .B1(new_n423), .B2(new_n873), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n423), .A2(new_n675), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n874), .A2(new_n891), .B1(new_n433), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n887), .B1(new_n893), .B2(KEYINPUT38), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT102), .B1(new_n894), .B2(KEYINPUT39), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n883), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n326), .A2(new_n723), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n839), .B1(new_n700), .B2(new_n842), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n318), .A2(new_n677), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n302), .B(new_n901), .C1(new_n324), .C2(new_n325), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT101), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n316), .A2(new_n318), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT101), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n302), .A4(new_n901), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n318), .B(new_n677), .C1(new_n316), .C2(new_n303), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n900), .A2(new_n888), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n651), .B2(new_n872), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n898), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n462), .B1(new_n702), .B2(new_n703), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n656), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n911), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n907), .B1(new_n902), .B2(KEYINPUT101), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n905), .B1(new_n319), .B2(new_n901), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n842), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n731), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n733), .B2(new_n705), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n725), .A2(new_n729), .ZN(new_n921));
  OAI211_X1 g0721(.A(KEYINPUT31), .B(new_n677), .C1(new_n921), .C2(new_n718), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT103), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n724), .A2(new_n730), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n925), .A2(KEYINPUT103), .A3(KEYINPUT31), .A4(new_n677), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n920), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT40), .B1(new_n886), .B2(new_n887), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(KEYINPUT104), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n918), .B(new_n928), .C1(new_n929), .C2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n894), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n561), .B1(new_n560), .B2(G200), .ZN(new_n934));
  AOI211_X1 g0734(.A(KEYINPUT79), .B(new_n360), .C1(new_n536), .C2(new_n538), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n660), .B1(new_n936), .B2(new_n565), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n937), .A2(new_n646), .A3(new_n611), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n506), .A2(new_n511), .A3(new_n519), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(new_n939), .A3(new_n723), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n731), .B1(new_n940), .B2(new_n706), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n924), .A2(new_n926), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n908), .B(new_n842), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n933), .B1(new_n943), .B2(KEYINPUT104), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n932), .B1(new_n944), .B2(new_n930), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n941), .A2(new_n942), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n463), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n945), .B(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(G330), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n914), .A2(new_n950), .B1(new_n244), .B2(new_n739), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n914), .A2(new_n950), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n866), .B1(new_n951), .B2(new_n952), .ZN(G367));
  NAND2_X1  g0753(.A1(new_n740), .A2(G1), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n677), .B1(new_n659), .B2(new_n556), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n567), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n660), .B2(new_n723), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT44), .B1(new_n691), .B2(new_n957), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n691), .A2(KEYINPUT45), .A3(new_n957), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT45), .B1(new_n691), .B2(new_n957), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n958), .B(new_n959), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT106), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n687), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n681), .A2(new_n686), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n688), .B1(new_n966), .B2(new_n687), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(new_n689), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n736), .ZN(new_n969));
  INV_X1    g0769(.A(new_n687), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n962), .A2(new_n963), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n965), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n737), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n694), .B(KEYINPUT41), .Z(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n954), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n689), .A2(new_n957), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT42), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n723), .A2(new_n626), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n645), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n647), .B2(new_n979), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT43), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n977), .A2(KEYINPUT42), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n660), .B1(new_n956), .B2(new_n610), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n723), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n978), .A2(new_n983), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT105), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n978), .A2(new_n984), .A3(new_n986), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n981), .B(new_n982), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n970), .A2(new_n957), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n981), .A2(new_n758), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n233), .A2(new_n754), .ZN(new_n995));
  INV_X1    g0795(.A(new_n760), .ZN(new_n996));
  INV_X1    g0796(.A(new_n444), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n996), .B1(new_n693), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n797), .A2(new_n344), .B1(new_n774), .B2(new_n794), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G143), .B2(new_n786), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n831), .A2(G68), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n771), .A2(new_n827), .B1(new_n779), .B2(new_n202), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n764), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n398), .B(new_n1003), .C1(new_n450), .C2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(KEYINPUT108), .B(G137), .Z(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n808), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1001), .A2(new_n1002), .A3(new_n1005), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT46), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n797), .B2(new_n484), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n778), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(new_n805), .C2(new_n774), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT107), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n808), .A2(G317), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n764), .A2(new_n545), .B1(new_n771), .B2(new_n798), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n398), .B1(new_n785), .B2(new_n802), .C1(new_n783), .C2(new_n436), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(G283), .C2(new_n780), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1015), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1009), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT47), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n759), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n746), .B1(new_n995), .B2(new_n999), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n976), .A2(new_n993), .B1(new_n994), .B2(new_n1026), .ZN(G387));
  AOI21_X1  g0827(.A(new_n968), .B1(G1), .B2(new_n740), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n686), .A2(new_n811), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n748), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1030), .A2(new_n696), .B1(G107), .B2(new_n213), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n230), .A2(G45), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n696), .B(new_n248), .C1(new_n276), .C2(new_n278), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT109), .Z(new_n1034));
  NOR2_X1   g0834(.A1(new_n341), .A2(G50), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n754), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1031), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n746), .B1(new_n1038), .B2(new_n996), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n808), .A2(G150), .B1(new_n390), .B2(new_n775), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n545), .B2(new_n766), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n778), .A2(new_n450), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n202), .B2(new_n771), .C1(new_n276), .C2(new_n779), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n831), .A2(new_n997), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n333), .C1(new_n794), .C2(new_n785), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT110), .Z(new_n1047));
  OAI22_X1  g0847(.A1(new_n785), .A2(new_n799), .B1(new_n774), .B2(new_n802), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT111), .Z(new_n1049));
  AOI22_X1  g0849(.A1(G317), .A2(new_n772), .B1(new_n780), .B2(G303), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT48), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G294), .A2(new_n778), .B1(new_n831), .B2(G283), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1052), .B2(KEYINPUT48), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1053), .A2(KEYINPUT49), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n333), .B1(new_n1004), .B2(G116), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n801), .C2(new_n793), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT49), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1047), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1039), .B1(new_n1061), .B2(new_n759), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1028), .B1(new_n1029), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n969), .A2(new_n695), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n968), .A2(new_n736), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1063), .A2(new_n1066), .ZN(G393));
  NAND2_X1  g0867(.A1(new_n965), .A2(new_n971), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1068), .A2(new_n694), .A3(new_n969), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n962), .B(new_n687), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1064), .B2(new_n954), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n760), .B1(new_n545), .B2(new_n213), .C1(new_n240), .C2(new_n754), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n746), .A2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G317), .A2(new_n786), .B1(new_n772), .B2(G311), .ZN(new_n1074));
  XOR2_X1   g0874(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1075));
  XNOR2_X1  g0875(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n768), .B(new_n1076), .C1(new_n799), .C2(new_n793), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n778), .A2(G283), .B1(G294), .B2(new_n780), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n333), .B1(new_n775), .B2(G303), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n484), .C2(new_n783), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n797), .A2(new_n276), .B1(new_n774), .B2(new_n202), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n783), .A2(new_n278), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n333), .B1(new_n779), .B2(new_n341), .ZN(new_n1083));
  OR3_X1    g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n785), .A2(new_n827), .B1(new_n771), .B2(new_n794), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1086), .B(new_n823), .C1(new_n826), .C2(new_n793), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1077), .A2(new_n1080), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1073), .B1(new_n1088), .B2(new_n759), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n957), .B2(new_n811), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1069), .A2(new_n1071), .A3(new_n1090), .ZN(G390));
  NAND2_X1  g0891(.A1(new_n895), .A2(new_n889), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n915), .A2(new_n916), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n897), .B1(new_n899), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1092), .A2(new_n1094), .A3(new_n882), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n897), .B(new_n894), .C1(new_n899), .C2(new_n1093), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n734), .A2(G330), .A3(new_n842), .A4(new_n908), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n842), .A2(G330), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n908), .C1(new_n941), .C2(new_n942), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n954), .B(new_n1098), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n896), .A2(new_n756), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n779), .A2(new_n545), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n436), .A2(new_n774), .B1(new_n771), .B2(new_n484), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G283), .C2(new_n786), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n333), .B(new_n1082), .C1(G87), .C2(new_n778), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n808), .A2(G294), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n833), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n778), .A2(G150), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT53), .Z(new_n1111));
  INV_X1    g0911(.A(KEYINPUT113), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1006), .A2(new_n774), .B1(new_n779), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n808), .A2(G125), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1111), .B(new_n1115), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G128), .A2(new_n786), .B1(new_n772), .B2(G132), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n398), .B1(new_n1004), .B2(G50), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n794), .C2(new_n783), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1109), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n759), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n816), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n747), .B1(new_n346), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1103), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1102), .A2(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1125), .A2(KEYINPUT114), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1098), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n928), .A2(G330), .A3(new_n462), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1128), .A2(new_n912), .A3(new_n656), .ZN(new_n1129));
  OAI211_X1 g0929(.A(G330), .B(new_n842), .C1(new_n732), .C2(new_n733), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1093), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1101), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n900), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n842), .A2(G330), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1093), .B1(new_n946), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(new_n899), .A3(new_n1097), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1129), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1127), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1137), .B(new_n1098), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n694), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1125), .A2(KEYINPUT114), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1126), .A2(new_n1141), .A3(new_n1142), .ZN(G378));
  XOR2_X1   g0943(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1144));
  NOR2_X1   g0944(.A1(new_n372), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n356), .A2(new_n872), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT55), .Z(new_n1148));
  NAND2_X1  g0948(.A1(new_n372), .A2(new_n1144), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1148), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n945), .A2(G330), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n945), .B2(G330), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n909), .B1(new_n651), .B2(new_n872), .C1(new_n896), .C2(new_n897), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n931), .B1(new_n888), .B2(new_n930), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(new_n943), .ZN(new_n1159));
  OAI21_X1  g0959(.A(KEYINPUT104), .B1(new_n946), .B2(new_n917), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n894), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1159), .B1(new_n1161), .B2(KEYINPUT40), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1152), .B1(new_n1162), .B2(new_n949), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n945), .A2(G330), .A3(new_n1153), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n911), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(KEYINPUT118), .B1(new_n1157), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1156), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1163), .A2(new_n911), .A3(new_n1164), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT118), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1129), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1140), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT57), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(new_n1167), .A3(new_n1168), .A4(KEYINPUT57), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT119), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n1140), .B2(new_n1172), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1179), .A2(KEYINPUT119), .A3(new_n1168), .A4(new_n1167), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1177), .A2(new_n694), .A3(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1174), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(G125), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n785), .A2(new_n1183), .B1(new_n774), .B2(new_n834), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n780), .A2(G137), .ZN(new_n1185));
  INV_X1    g0985(.A(G128), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1185), .B1(new_n1186), .B2(new_n771), .C1(new_n797), .C2(new_n1113), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1184), .B(new_n1187), .C1(G150), .C2(new_n831), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n808), .A2(G124), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n1004), .C2(G159), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n333), .A2(G41), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n545), .B2(new_n774), .C1(new_n436), .C2(new_n771), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n786), .A2(G116), .B1(new_n780), .B2(new_n997), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1004), .A2(G58), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1197), .A2(new_n1042), .A3(new_n1002), .A4(new_n1198), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1196), .B(new_n1199), .C1(G283), .C2(new_n808), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G50), .B(new_n1195), .C1(new_n491), .C2(new_n247), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT115), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1194), .A2(new_n1201), .A3(new_n1202), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n759), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT116), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n741), .B(new_n1207), .C1(new_n202), .C2(new_n815), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1153), .A2(new_n756), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1171), .B2(new_n954), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1182), .A2(new_n1212), .ZN(G375));
  NAND3_X1  g1013(.A1(new_n1133), .A2(new_n1129), .A3(new_n1136), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1138), .A2(new_n975), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1093), .A2(new_n756), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n746), .B1(G68), .B2(new_n816), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n766), .A2(new_n278), .B1(new_n793), .B2(new_n798), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n333), .B1(new_n778), .B2(G97), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G116), .A2(new_n775), .B1(new_n772), .B2(G283), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n786), .A2(G294), .B1(new_n780), .B2(G107), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1044), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n774), .A2(new_n1113), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n778), .B2(G159), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n827), .B2(new_n779), .C1(new_n793), .C2(new_n1186), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n772), .A2(new_n1007), .B1(new_n786), .B2(G132), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n831), .A2(G50), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1227), .A2(new_n333), .A3(new_n1198), .A4(new_n1228), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1219), .A2(new_n1223), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1218), .B1(new_n1230), .B2(new_n759), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1216), .A2(new_n954), .B1(new_n1217), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1215), .A2(new_n1232), .ZN(G381));
  INV_X1    g1033(.A(G378), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1182), .A2(new_n1234), .A3(new_n1212), .ZN(new_n1235));
  OR4_X1    g1035(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1236));
  OR4_X1    g1036(.A1(G387), .A2(new_n1235), .A3(G381), .A4(new_n1236), .ZN(G407));
  NAND2_X1  g1037(.A1(new_n676), .A2(G213), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT120), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G407), .B(G213), .C1(new_n1235), .C2(new_n1240), .ZN(G409));
  INV_X1    g1041(.A(KEYINPUT124), .ZN(new_n1242));
  INV_X1    g1042(.A(G396), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(G393), .B(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G387), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1244), .B1(G387), .B2(KEYINPUT123), .ZN(new_n1247));
  INV_X1    g1047(.A(G390), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G387), .A2(KEYINPUT123), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1244), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G390), .B1(new_n1252), .B2(new_n1245), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1249), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1242), .B1(new_n1254), .B2(KEYINPUT61), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  OAI211_X1 g1056(.A(KEYINPUT124), .B(new_n1256), .C1(new_n1249), .C2(new_n1253), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G378), .B(new_n1212), .C1(new_n1174), .C2(new_n1181), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1169), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n975), .B(new_n1173), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1167), .A2(new_n1168), .A3(new_n954), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1210), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT121), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1262), .A2(KEYINPUT121), .A3(new_n1210), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1261), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1234), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1239), .B1(new_n1258), .B2(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1214), .B(KEYINPUT60), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(new_n694), .A3(new_n1138), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1271), .A2(G384), .A3(new_n1232), .ZN(new_n1272));
  AOI21_X1  g1072(.A(G384), .B1(new_n1271), .B2(new_n1232), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1255), .A2(new_n1257), .B1(new_n1269), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1258), .A2(new_n1268), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n1238), .A3(new_n1274), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1274), .A2(G213), .A3(new_n676), .A4(G2897), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1239), .A2(G2897), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1282), .A2(KEYINPUT122), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT122), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1279), .A2(new_n1238), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1276), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1278), .B1(new_n1281), .B2(new_n1289), .ZN(new_n1290));
  XOR2_X1   g1090(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1291));
  INV_X1    g1091(.A(new_n1269), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1287), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1280), .A2(KEYINPUT126), .A3(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1269), .A2(KEYINPUT62), .A3(new_n1274), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT126), .B1(new_n1280), .B2(new_n1294), .ZN(new_n1298));
  OAI211_X1 g1098(.A(KEYINPUT127), .B(new_n1293), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1254), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1280), .A2(new_n1294), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT127), .B1(new_n1304), .B2(new_n1293), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1290), .B1(new_n1300), .B2(new_n1305), .ZN(G405));
  XNOR2_X1  g1106(.A(new_n1254), .B(new_n1275), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G375), .A2(G378), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1235), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1307), .B(new_n1309), .ZN(G402));
endmodule


