//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(KEYINPUT1), .ZN(new_n202));
  OAI21_X1  g001(.A(new_n202), .B1(G113gat), .B2(G120gat), .ZN(new_n203));
  AND2_X1   g002(.A1(G113gat), .A2(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT68), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n206), .B(KEYINPUT68), .C1(new_n204), .C2(new_n203), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT69), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT25), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n214));
  AND2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  AND4_X1   g017(.A1(new_n212), .A2(new_n214), .A3(new_n216), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n214), .A2(new_n216), .A3(new_n218), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n225), .A2(new_n226), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n231), .B1(new_n220), .B2(new_n221), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n231), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n229), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n228), .B1(new_n236), .B2(new_n212), .ZN(new_n237));
  INV_X1    g036(.A(new_n220), .ZN(new_n238));
  OAI211_X1 g037(.A(KEYINPUT65), .B(new_n224), .C1(new_n223), .C2(KEYINPUT27), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT28), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT27), .ZN(new_n242));
  AOI21_X1  g041(.A(G190gat), .B1(new_n242), .B2(G183gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n238), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(KEYINPUT26), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT67), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n213), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G169gat), .ZN(new_n252));
  INV_X1    g051(.A(G176gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n254), .B(KEYINPUT66), .C1(new_n215), .C2(KEYINPUT26), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(new_n213), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n251), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n239), .A2(new_n243), .A3(new_n240), .A4(new_n244), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n246), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n211), .B1(new_n237), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n215), .B1(new_n254), .B2(new_n217), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n225), .B(new_n226), .C1(new_n234), .C2(new_n231), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n214), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n266), .A2(KEYINPUT25), .B1(new_n227), .B2(new_n219), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n246), .A2(new_n259), .A3(new_n260), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(KEYINPUT69), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n210), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT69), .B1(new_n267), .B2(new_n268), .ZN(new_n271));
  INV_X1    g070(.A(new_n210), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275));
  AND4_X1   g074(.A1(KEYINPUT73), .A2(new_n274), .A3(KEYINPUT34), .A4(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n277), .B1(new_n274), .B2(new_n275), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n266), .A2(KEYINPUT25), .ZN(new_n281));
  AND4_X1   g080(.A1(KEYINPUT69), .A2(new_n268), .A3(new_n281), .A4(new_n228), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n272), .B1(new_n282), .B2(new_n271), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n210), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n275), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT71), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G15gat), .B(G43gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(G71gat), .B(G99gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n275), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n270), .B2(new_n273), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n293), .B2(KEYINPUT32), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n295), .A3(new_n286), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n288), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n288), .A2(new_n294), .A3(KEYINPUT72), .A4(new_n296), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n291), .A2(new_n286), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n285), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n280), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g105(.A(new_n304), .B(new_n279), .C1(new_n299), .C2(new_n300), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n267), .A2(new_n268), .ZN(new_n309));
  AND2_X1   g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n312));
  NAND2_X1  g111(.A1(G211gat), .A2(G218gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT22), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(KEYINPUT74), .A3(new_n314), .ZN(new_n318));
  XNOR2_X1  g117(.A(G197gat), .B(G204gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n321));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n320), .B2(new_n321), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n312), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n322), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(KEYINPUT75), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT76), .A3(new_n323), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT29), .B1(new_n267), .B2(new_n268), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n311), .B(new_n331), .C1(new_n310), .C2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n310), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n311), .A2(KEYINPUT77), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n309), .A2(new_n336), .A3(new_n310), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n333), .B1(new_n338), .B2(new_n331), .ZN(new_n339));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT78), .ZN(new_n341));
  XNOR2_X1  g140(.A(G64gat), .B(G92gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT80), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n349), .A3(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n333), .ZN(new_n352));
  INV_X1    g151(.A(new_n334), .ZN(new_n353));
  INV_X1    g152(.A(new_n337), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n336), .B1(new_n309), .B2(new_n310), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n331), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n352), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n343), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n339), .A2(KEYINPUT30), .A3(new_n344), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n351), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G141gat), .ZN(new_n364));
  INV_X1    g163(.A(G148gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(KEYINPUT81), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G155gat), .B(G162gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G155gat), .ZN(new_n371));
  INV_X1    g170(.A(G162gat), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT2), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n366), .A2(new_n367), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n366), .A3(new_n367), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(new_n369), .A3(new_n368), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n377), .A3(KEYINPUT3), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n272), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n210), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n378), .A2(new_n210), .A3(KEYINPUT4), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(KEYINPUT83), .A2(KEYINPUT5), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n378), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT4), .B1(new_n378), .B2(new_n210), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n394), .A2(new_n386), .A3(new_n382), .A4(new_n389), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT0), .ZN(new_n398));
  XNOR2_X1  g197(.A(G57gat), .B(G85gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n378), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n272), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n383), .ZN(new_n404));
  INV_X1    g203(.A(new_n386), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(KEYINPUT5), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n396), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT6), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n401), .B1(new_n396), .B2(new_n406), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n363), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n380), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n331), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n379), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n328), .A2(new_n327), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n320), .B2(new_n322), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n419), .B1(new_n423), .B2(new_n378), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n329), .A2(new_n416), .A3(new_n323), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT3), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n378), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n426), .B1(new_n418), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n430), .A3(G22gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(G22gat), .B1(new_n425), .B2(new_n430), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n434));
  XNOR2_X1  g233(.A(G78gat), .B(G106gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT31), .B(G50gat), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n435), .B(new_n436), .Z(new_n437));
  OAI22_X1  g236(.A1(new_n432), .A2(new_n433), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n433), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n431), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n437), .B(KEYINPUT84), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n308), .A2(new_n415), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT35), .ZN(new_n444));
  INV_X1    g243(.A(new_n441), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n439), .A2(new_n445), .A3(new_n431), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n306), .A2(new_n307), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n361), .B1(new_n348), .B2(new_n350), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT86), .B1(new_n412), .B2(new_n410), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n396), .A2(new_n406), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n400), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n411), .A4(new_n407), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n450), .A2(new_n409), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT87), .B(KEYINPUT35), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n448), .A2(new_n449), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n301), .A2(new_n305), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n279), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n301), .A2(new_n305), .A3(new_n280), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT36), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n306), .B2(new_n307), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n442), .B1(new_n449), .B2(new_n413), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n353), .B(new_n331), .C1(new_n354), .C2(new_n355), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n311), .B1(new_n332), .B2(new_n310), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(new_n357), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT38), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(new_n343), .C1(new_n358), .C2(KEYINPUT37), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n345), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT38), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n344), .B1(new_n339), .B2(new_n468), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n358), .A2(KEYINPUT37), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n447), .B1(new_n455), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n382), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n385), .A2(new_n387), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n405), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n482), .A2(KEYINPUT39), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n482), .B(KEYINPUT39), .C1(new_n405), .C2(new_n404), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n400), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n486), .A2(KEYINPUT85), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n407), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n487), .B2(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n363), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n466), .B1(new_n479), .B2(new_n490), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n444), .A2(new_n458), .B1(new_n465), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT18), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  OR2_X1    g293(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OR3_X1    g296(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n497), .A2(G29gat), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G43gat), .B(G50gat), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n501), .A2(KEYINPUT90), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT15), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n501), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n498), .A2(new_n499), .ZN(new_n506));
  INV_X1    g305(.A(G29gat), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n495), .B2(new_n496), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n505), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n500), .A2(new_n502), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n494), .B(new_n504), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G8gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(G1gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G1gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT16), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(KEYINPUT93), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT93), .ZN(new_n522));
  INV_X1    g321(.A(new_n520), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(new_n516), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(KEYINPUT91), .ZN(new_n526));
  XOR2_X1   g325(.A(G15gat), .B(G22gat), .Z(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT92), .A3(new_n518), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT91), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n515), .A2(new_n529), .A3(new_n519), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(new_n515), .B2(G1gat), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n526), .A2(new_n528), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G8gat), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n512), .B1(new_n509), .B2(new_n510), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT17), .B1(new_n536), .B2(new_n503), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n536), .A2(new_n503), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n534), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n513), .A2(new_n535), .A3(new_n537), .A4(new_n539), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n493), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(new_n543), .B2(new_n544), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT18), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n546), .B(KEYINPUT13), .Z(new_n551));
  AND2_X1   g350(.A1(new_n540), .A2(new_n541), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n540), .A2(new_n541), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G113gat), .B(G141gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G169gat), .B(G197gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT12), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n548), .A2(new_n550), .A3(new_n554), .A4(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n554), .B1(new_n549), .B2(KEYINPUT18), .ZN(new_n563));
  AOI211_X1 g362(.A(new_n493), .B(new_n547), .C1(new_n543), .C2(new_n544), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n492), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT21), .ZN(new_n569));
  INV_X1    g368(.A(G64gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT95), .B1(new_n570), .B2(G57gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n572));
  INV_X1    g371(.A(G57gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(G64gat), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n571), .B(new_n574), .C1(new_n573), .C2(G64gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  OR2_X1    g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n570), .A2(G57gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n573), .A2(G64gat), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT9), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n577), .A2(new_n576), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n535), .B1(new_n569), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT96), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G155gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n588), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n569), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G127gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n591), .A2(new_n598), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT7), .ZN(new_n603));
  OR2_X1    g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(G85gat), .A2(G92gat), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(KEYINPUT8), .B2(new_n605), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n606), .B1(new_n603), .B2(new_n608), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n513), .A2(new_n537), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n540), .A2(new_n612), .ZN(new_n615));
  NAND2_X1  g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G190gat), .B(G218gat), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT97), .ZN(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n620), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n614), .A2(new_n626), .A3(new_n615), .A4(new_n618), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n621), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n625), .B1(new_n621), .B2(new_n627), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n601), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT98), .B1(new_n603), .B2(new_n608), .ZN(new_n633));
  OAI22_X1  g432(.A1(new_n586), .A2(new_n633), .B1(new_n610), .B2(new_n611), .ZN(new_n634));
  INV_X1    g433(.A(new_n611), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n579), .A2(new_n575), .B1(new_n583), .B2(new_n584), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n603), .A2(new_n608), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n635), .A2(new_n636), .A3(new_n639), .A4(new_n609), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n634), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n636), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n634), .A2(new_n640), .ZN(new_n647));
  INV_X1    g446(.A(new_n645), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT99), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n646), .A2(new_n649), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n632), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n568), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n413), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n518), .ZN(G1324gat));
  NAND3_X1  g463(.A1(new_n568), .A2(new_n363), .A3(new_n661), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n665), .A2(G8gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT16), .B(G8gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT42), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(KEYINPUT42), .B2(new_n668), .ZN(G1325gat));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT36), .B1(new_n460), .B2(new_n461), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n306), .A2(new_n307), .A3(new_n463), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT101), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G15gat), .B1(new_n662), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n308), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(G15gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n662), .B2(new_n680), .ZN(G1326gat));
  NOR2_X1   g480(.A1(new_n662), .A2(new_n442), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT43), .B(G22gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  INV_X1    g483(.A(new_n601), .ZN(new_n685));
  INV_X1    g484(.A(new_n631), .ZN(new_n686));
  INV_X1    g485(.A(new_n660), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n568), .A2(new_n685), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n688), .A2(G29gat), .A3(new_n413), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(KEYINPUT45), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n491), .A3(new_n675), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n444), .A2(new_n458), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n629), .B2(new_n630), .ZN(new_n695));
  INV_X1    g494(.A(new_n630), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(new_n628), .A3(KEYINPUT103), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(KEYINPUT44), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n492), .B2(new_n631), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n660), .B(KEYINPUT102), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(new_n567), .A3(new_n601), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n413), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n689), .A2(KEYINPUT45), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n690), .A2(new_n708), .A3(new_n709), .ZN(G1328gat));
  NOR3_X1   g509(.A1(new_n688), .A2(new_n449), .A3(new_n497), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT46), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n497), .B1(new_n707), .B2(new_n449), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1329gat));
  OAI21_X1  g513(.A(G43gat), .B1(new_n707), .B2(new_n677), .ZN(new_n715));
  OR3_X1    g514(.A1(new_n688), .A2(G43gat), .A3(new_n679), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n715), .A2(KEYINPUT47), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n707), .B2(new_n442), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n688), .A2(G50gat), .A3(new_n442), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(KEYINPUT48), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1331gat));
  NOR3_X1   g527(.A1(new_n632), .A2(new_n704), .A3(new_n566), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n693), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n413), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(new_n573), .ZN(G1332gat));
  INV_X1    g531(.A(new_n730), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n449), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT104), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n736), .B(new_n737), .Z(G1333gat));
  NOR3_X1   g537(.A1(new_n730), .A2(G71gat), .A3(new_n679), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n733), .A2(new_n676), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(G71gat), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n733), .A2(new_n447), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g543(.A1(new_n601), .A2(new_n566), .A3(new_n687), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n703), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746), .B2(new_n413), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n601), .A2(new_n566), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n686), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT51), .B1(new_n693), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  AOI211_X1 g551(.A(new_n752), .B(new_n749), .C1(new_n691), .C2(new_n692), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n687), .A2(G85gat), .A3(new_n413), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT105), .Z(new_n756));
  OAI21_X1  g555(.A(new_n747), .B1(new_n754), .B2(new_n756), .ZN(G1336gat));
  OAI21_X1  g556(.A(G92gat), .B1(new_n746), .B2(new_n449), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n449), .A2(G92gat), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n705), .B(new_n759), .C1(new_n751), .C2(new_n753), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT52), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n758), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1337gat));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n766));
  INV_X1    g565(.A(G99gat), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n703), .A2(new_n745), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(new_n676), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n308), .A2(new_n767), .A3(new_n660), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT106), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n754), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n766), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G99gat), .B1(new_n746), .B2(new_n677), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n774), .B(KEYINPUT107), .C1(new_n754), .C2(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1338gat));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n442), .A2(G106gat), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n705), .B(new_n778), .C1(new_n751), .C2(new_n753), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n465), .A2(new_n491), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT35), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n448), .B2(new_n415), .ZN(new_n783));
  AND4_X1   g582(.A1(new_n308), .A2(new_n449), .A3(new_n442), .A4(new_n457), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n780), .B1(new_n785), .B2(new_n686), .ZN(new_n786));
  INV_X1    g585(.A(new_n700), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n691), .B2(new_n692), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n447), .B(new_n745), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT109), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G106gat), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n789), .A2(KEYINPUT109), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n777), .B(new_n779), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n789), .A2(KEYINPUT108), .A3(G106gat), .ZN(new_n794));
  INV_X1    g593(.A(new_n779), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT108), .B1(new_n789), .B2(G106gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n793), .B1(new_n797), .B2(new_n777), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n563), .A2(new_n564), .A3(new_n562), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n543), .A2(new_n547), .A3(new_n544), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n552), .A2(new_n553), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n551), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n559), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT112), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n561), .A2(new_n807), .A3(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n642), .A2(new_n648), .A3(new_n643), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n646), .A2(KEYINPUT54), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT110), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n646), .A2(new_n812), .A3(KEYINPUT54), .A4(new_n809), .ZN(new_n813));
  XNOR2_X1  g612(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n644), .A2(new_n645), .A3(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n654), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n657), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n654), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(KEYINPUT110), .B2(new_n810), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT55), .B1(new_n820), .B2(new_n813), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n806), .A2(new_n698), .A3(new_n808), .A4(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n566), .A2(new_n822), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n660), .A2(new_n561), .A3(new_n804), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n698), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n799), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n800), .A2(new_n805), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n660), .A2(new_n829), .B1(new_n566), .B2(new_n822), .ZN(new_n830));
  OAI211_X1 g629(.A(KEYINPUT113), .B(new_n823), .C1(new_n830), .C2(new_n698), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n685), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n661), .A2(new_n567), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n413), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n449), .A3(new_n448), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT115), .ZN(new_n836));
  INV_X1    g635(.A(G113gat), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(new_n837), .A3(new_n566), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n447), .B1(new_n832), .B2(new_n833), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n363), .A2(new_n413), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n679), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(new_n566), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n839), .B1(new_n844), .B2(G113gat), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n844), .A2(new_n839), .A3(G113gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n838), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  NOR2_X1   g646(.A1(new_n687), .A2(G120gat), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT116), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n836), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n840), .A2(new_n843), .ZN(new_n851));
  OAI21_X1  g650(.A(G120gat), .B1(new_n851), .B2(new_n704), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1341gat));
  OAI21_X1  g652(.A(G127gat), .B1(new_n851), .B2(new_n685), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n601), .A2(new_n595), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n835), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT117), .Z(G1342gat));
  OR3_X1    g656(.A1(new_n835), .A2(G134gat), .A3(new_n631), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n851), .B2(new_n631), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(G1343gat));
  NOR2_X1   g661(.A1(new_n676), .A2(new_n442), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n834), .A2(new_n863), .A3(new_n449), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n566), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n825), .A2(new_n826), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n631), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n601), .B1(new_n868), .B2(new_n823), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n632), .A2(new_n566), .A3(new_n660), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n447), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT57), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n676), .A2(new_n842), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n442), .B1(new_n832), .B2(new_n833), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n567), .A2(new_n364), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n866), .A2(new_n364), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT58), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n877), .A2(new_n878), .ZN(new_n883));
  AOI21_X1  g682(.A(G141gat), .B1(new_n865), .B2(new_n566), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT118), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n881), .A2(new_n885), .ZN(G1344gat));
  NAND3_X1  g685(.A1(new_n865), .A2(new_n365), .A3(new_n660), .ZN(new_n887));
  AOI211_X1 g686(.A(KEYINPUT59), .B(new_n365), .C1(new_n877), .C2(new_n660), .ZN(new_n888));
  XOR2_X1   g687(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n889));
  NOR2_X1   g688(.A1(new_n442), .A2(KEYINPUT57), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n806), .A2(new_n686), .A3(new_n808), .A4(new_n822), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n868), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n685), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n891), .B1(new_n894), .B2(new_n833), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n832), .A2(new_n833), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n447), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(KEYINPUT57), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n873), .A3(new_n660), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n889), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n887), .B1(new_n888), .B2(new_n900), .ZN(G1345gat));
  AOI21_X1  g700(.A(G155gat), .B1(new_n865), .B2(new_n601), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n601), .A2(G155gat), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT120), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n877), .B2(new_n904), .ZN(G1346gat));
  AOI21_X1  g704(.A(G162gat), .B1(new_n865), .B2(new_n686), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n699), .A2(new_n372), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n877), .B2(new_n907), .ZN(G1347gat));
  NAND4_X1  g707(.A1(new_n840), .A2(new_n413), .A3(new_n308), .A4(new_n363), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n252), .A3(new_n567), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n414), .B1(new_n832), .B2(new_n833), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n448), .A2(new_n363), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT121), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n566), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n910), .B1(new_n919), .B2(new_n252), .ZN(G1348gat));
  OAI21_X1  g719(.A(G176gat), .B1(new_n909), .B2(new_n704), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n687), .A2(G176gat), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n917), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(G1349gat));
  OAI21_X1  g725(.A(G183gat), .B1(new_n909), .B2(new_n685), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n242), .A2(G183gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n601), .A2(new_n928), .A3(new_n244), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n927), .B1(new_n913), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n909), .B2(new_n631), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT61), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n699), .A2(G190gat), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n918), .A2(KEYINPUT123), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT123), .B1(new_n918), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1351gat));
  NAND3_X1  g736(.A1(new_n911), .A2(new_n863), .A3(new_n363), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(G197gat), .B1(new_n939), .B2(new_n566), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n894), .A2(new_n833), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n890), .ZN(new_n942));
  AND4_X1   g741(.A1(new_n413), .A2(new_n674), .A3(new_n363), .A4(new_n675), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n942), .B(new_n943), .C1(new_n876), .C2(new_n875), .ZN(new_n944));
  INV_X1    g743(.A(G197gat), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n944), .A2(new_n945), .A3(new_n567), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n940), .A2(new_n946), .ZN(G1352gat));
  OAI21_X1  g746(.A(G204gat), .B1(new_n944), .B2(new_n704), .ZN(new_n948));
  OR3_X1    g747(.A1(new_n938), .A2(G204gat), .A3(new_n687), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n949), .A2(new_n951), .A3(KEYINPUT62), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n949), .B2(KEYINPUT62), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n948), .B(new_n950), .C1(new_n952), .C2(new_n953), .ZN(G1353gat));
  INV_X1    g753(.A(G211gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n955), .A3(new_n601), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n957), .A2(KEYINPUT126), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n898), .A2(new_n959), .A3(new_n601), .A4(new_n943), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT125), .B1(new_n944), .B2(new_n685), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n955), .B1(KEYINPUT126), .B2(new_n957), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n958), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n958), .ZN(new_n965));
  INV_X1    g764(.A(new_n963), .ZN(new_n966));
  AOI211_X1 g765(.A(new_n965), .B(new_n966), .C1(new_n960), .C2(new_n961), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n956), .B1(new_n964), .B2(new_n967), .ZN(G1354gat));
  AND2_X1   g767(.A1(new_n944), .A2(KEYINPUT127), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n686), .B1(new_n944), .B2(KEYINPUT127), .ZN(new_n970));
  OAI21_X1  g769(.A(G218gat), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n699), .A2(G218gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n938), .B2(new_n972), .ZN(G1355gat));
endmodule


