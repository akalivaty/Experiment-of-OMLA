//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n580, new_n581, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n594, new_n595,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n644,
    new_n647, new_n649, new_n650, new_n651, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n450), .B(new_n451), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT69), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n467), .A2(new_n468), .A3(G137), .A4(new_n461), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n462), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n471), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  AOI211_X1 g050(.A(KEYINPUT68), .B(new_n461), .C1(new_n472), .C2(new_n473), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT70), .ZN(G160));
  NOR2_X1   g053(.A1(new_n463), .A2(new_n464), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(new_n461), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G138), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n467), .A2(KEYINPUT4), .A3(G138), .A4(new_n461), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n467), .A2(G126), .A3(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  OAI21_X1  g074(.A(G62), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(KEYINPUT71), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G62), .C1(new_n498), .C2(new_n499), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n497), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(G50), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n498), .A2(new_n499), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n504), .A2(new_n511), .ZN(G166));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n513), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(new_n497), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(KEYINPUT72), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT73), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n514), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n523), .A2(new_n519), .A3(KEYINPUT73), .A4(G543), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(G51), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n529), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n509), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n530), .B(new_n532), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT74), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G51), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n523), .A2(new_n519), .A3(G543), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n538), .B1(new_n541), .B2(new_n524), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n543));
  NOR3_X1   g118(.A1(new_n542), .A2(new_n543), .A3(new_n535), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n537), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n506), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n527), .A2(new_n528), .B1(new_n517), .B2(new_n518), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G90), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n541), .A2(new_n524), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n553), .B1(new_n554), .B2(G52), .ZN(G171));
  NAND2_X1  g130(.A1(new_n551), .A2(G81), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n557));
  OAI21_X1  g132(.A(G56), .B1(new_n498), .B2(new_n499), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n557), .B1(new_n560), .B2(G651), .ZN(new_n561));
  AOI211_X1 g136(.A(KEYINPUT75), .B(new_n497), .C1(new_n558), .C2(new_n559), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n556), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n541), .B2(new_n524), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT76), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n556), .ZN(new_n567));
  INV_X1    g142(.A(new_n559), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n529), .B2(G56), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT75), .B1(new_n569), .B2(new_n497), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n560), .A2(new_n557), .A3(G651), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(G43), .B1(new_n520), .B2(new_n525), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G860), .ZN(G153));
  NAND4_X1  g153(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g154(.A1(G1), .A2(G3), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT8), .ZN(new_n581));
  NAND4_X1  g156(.A1(G319), .A2(G483), .A3(G661), .A4(new_n581), .ZN(G188));
  INV_X1    g157(.A(G53), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT9), .B1(new_n539), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT9), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n515), .A2(new_n585), .A3(G53), .A4(new_n519), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n529), .A2(new_n509), .A3(G91), .ZN(new_n588));
  XNOR2_X1  g163(.A(KEYINPUT77), .B(G65), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n529), .A2(new_n589), .B1(G78), .B2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n590), .B2(new_n497), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n587), .A2(new_n592), .ZN(G299));
  NOR2_X1   g168(.A1(new_n520), .A2(new_n525), .ZN(new_n594));
  INV_X1    g169(.A(G52), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n550), .B(new_n552), .C1(new_n594), .C2(new_n595), .ZN(G301));
  OAI21_X1  g171(.A(KEYINPUT78), .B1(new_n504), .B2(new_n511), .ZN(new_n597));
  NAND2_X1  g172(.A1(G75), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G62), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n527), .B2(new_n528), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n600), .B2(new_n502), .ZN(new_n601));
  INV_X1    g176(.A(new_n503), .ZN(new_n602));
  OAI21_X1  g177(.A(G651), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n603), .A2(new_n604), .A3(new_n510), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n597), .A2(new_n605), .ZN(G303));
  NAND3_X1  g181(.A1(new_n515), .A2(G49), .A3(new_n519), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n551), .A2(G87), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(G288));
  INV_X1    g185(.A(G61), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n527), .B2(new_n528), .ZN(new_n612));
  AND2_X1   g187(.A1(G73), .A2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(G651), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G86), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n527), .B2(new_n528), .ZN(new_n616));
  AND2_X1   g191(.A1(G48), .A2(G543), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n509), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(G305));
  NAND2_X1  g194(.A1(G72), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G60), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n506), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n622), .A2(G651), .B1(new_n551), .B2(G85), .ZN(new_n623));
  INV_X1    g198(.A(G47), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n594), .B2(new_n624), .ZN(G290));
  NAND2_X1  g200(.A1(G301), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(G54), .B1(new_n520), .B2(new_n525), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n551), .B2(G92), .ZN(new_n630));
  AND4_X1   g205(.A1(new_n629), .A2(new_n529), .A3(new_n509), .A4(G92), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g207(.A1(new_n529), .A2(G66), .ZN(new_n633));
  NAND2_X1  g208(.A1(G79), .A2(G543), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT80), .Z(new_n635));
  OAI21_X1  g210(.A(G651), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G92), .ZN(new_n637));
  OAI21_X1  g212(.A(KEYINPUT79), .B1(new_n533), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n551), .A2(new_n629), .A3(G92), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT10), .A3(new_n639), .ZN(new_n640));
  AND4_X1   g215(.A1(new_n627), .A2(new_n632), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n626), .B1(new_n641), .B2(G868), .ZN(G284));
  OAI21_X1  g217(.A(new_n626), .B1(new_n641), .B2(G868), .ZN(G321));
  NOR2_X1   g218(.A1(G299), .A2(G868), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(G168), .B2(G868), .ZN(G297));
  XOR2_X1   g220(.A(G297), .B(KEYINPUT81), .Z(G280));
  INV_X1    g221(.A(G559), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n641), .B1(new_n647), .B2(G860), .ZN(G148));
  NAND2_X1  g223(.A1(new_n641), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G868), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n577), .B2(G868), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT82), .Z(G323));
  XNOR2_X1  g227(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g228(.A1(G123), .A2(new_n482), .B1(new_n480), .B2(G135), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n656));
  INV_X1    g231(.A(G111), .ZN(new_n657));
  AOI22_X1  g232(.A1(new_n655), .A2(new_n656), .B1(new_n657), .B2(G2105), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n656), .B2(new_n655), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(G2096), .Z(new_n661));
  XOR2_X1   g236(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT13), .ZN(new_n665));
  INV_X1    g240(.A(G2100), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n661), .A2(new_n667), .A3(new_n668), .ZN(G156));
  INV_X1    g244(.A(KEYINPUT14), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2427), .B(G2438), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2430), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT15), .B(G2435), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n673), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2451), .B(G2454), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT16), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1341), .B(G1348), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2443), .B(G2446), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G14), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(G401));
  XOR2_X1   g260(.A(G2072), .B(G2078), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  XOR2_X1   g263(.A(G2084), .B(G2090), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT18), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n686), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n688), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI211_X1 g270(.A(new_n689), .B(new_n695), .C1(new_n694), .C2(new_n686), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n694), .A2(new_n689), .ZN(new_n697));
  AOI211_X1 g272(.A(new_n691), .B(new_n696), .C1(new_n693), .C2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G2096), .B(G2100), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G227));
  XOR2_X1   g276(.A(G1971), .B(G1976), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT19), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1956), .B(G2474), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1961), .B(G1966), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n703), .A2(new_n706), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT20), .Z(new_n710));
  AOI211_X1 g285(.A(new_n708), .B(new_n710), .C1(new_n703), .C2(new_n707), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1991), .B(G1996), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1981), .B(G1986), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(G229));
  NOR2_X1   g292(.A1(G6), .A2(G16), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n614), .A2(new_n618), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT32), .ZN(new_n721));
  INV_X1    g296(.A(G1981), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G22), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G166), .B2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(G1971), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(G23), .ZN(new_n729));
  INV_X1    g304(.A(G288), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n724), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT33), .B(G1976), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n723), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(KEYINPUT34), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT88), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n724), .A2(G24), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n624), .B1(new_n541), .B2(new_n524), .ZN(new_n738));
  INV_X1    g313(.A(new_n623), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n737), .B1(new_n740), .B2(new_n724), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT87), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1986), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n734), .A2(KEYINPUT34), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n480), .A2(G131), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n482), .A2(G119), .ZN(new_n746));
  OR2_X1    g321(.A1(G95), .A2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n747), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  MUX2_X1   g324(.A(G25), .B(new_n749), .S(G29), .Z(new_n750));
  XOR2_X1   g325(.A(KEYINPUT35), .B(G1991), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT86), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n750), .B(new_n752), .Z(new_n753));
  NAND4_X1  g328(.A1(new_n736), .A2(new_n743), .A3(new_n744), .A4(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G32), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n482), .A2(G129), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT93), .Z(new_n760));
  AND3_X1   g335(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT26), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n761), .B(new_n763), .C1(G141), .C2(new_n480), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n758), .B1(new_n766), .B2(new_n757), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(G160), .A2(G29), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT24), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n757), .B1(new_n772), .B2(G34), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(KEYINPUT91), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n772), .B2(G34), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(KEYINPUT91), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT97), .Z(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n724), .A2(G5), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G171), .B2(new_n724), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT96), .Z(new_n785));
  AOI211_X1 g360(.A(new_n770), .B(new_n781), .C1(new_n782), .C2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT98), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n577), .A2(new_n724), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n724), .B2(G19), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G1341), .ZN(new_n792));
  NOR2_X1   g367(.A1(G29), .A2(G33), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT89), .Z(new_n794));
  AND2_X1   g369(.A1(new_n467), .A2(G127), .ZN(new_n795));
  AND2_X1   g370(.A1(G115), .A2(G2104), .ZN(new_n796));
  OAI21_X1  g371(.A(G2105), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT25), .ZN(new_n798));
  NAND2_X1  g373(.A1(G103), .A2(G2104), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(G2105), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n480), .A2(G139), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n794), .B1(new_n803), .B2(new_n757), .ZN(new_n804));
  INV_X1    g379(.A(G2072), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT92), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n757), .A2(G35), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G162), .B2(new_n757), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT29), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n807), .B1(G2090), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n757), .A2(G26), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT28), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n480), .A2(G140), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n482), .A2(G128), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n461), .A2(G116), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n814), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n813), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G2067), .ZN(new_n820));
  INV_X1    g395(.A(G2078), .ZN(new_n821));
  NAND2_X1  g396(.A1(G164), .A2(G29), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G27), .B2(G29), .ZN(new_n823));
  OAI221_X1 g398(.A(new_n820), .B1(new_n821), .B2(new_n823), .C1(new_n767), .C2(new_n769), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n804), .A2(new_n805), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT90), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G11), .ZN(new_n828));
  INV_X1    g403(.A(G28), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(KEYINPUT30), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT95), .ZN(new_n831));
  AOI21_X1  g406(.A(G29), .B1(new_n829), .B2(KEYINPUT30), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n757), .B2(new_n660), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n821), .B2(new_n823), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n826), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n811), .A2(new_n824), .A3(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n785), .A2(new_n782), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n791), .A2(G1341), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n792), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(G16), .A2(G21), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G168), .B2(G16), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G1966), .ZN(new_n843));
  NOR2_X1   g418(.A1(G4), .A2(G16), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n641), .B2(G16), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(G1348), .Z(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n779), .B2(new_n778), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n810), .A2(G2090), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n724), .A2(G20), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT23), .Z(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G299), .B2(G16), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G1956), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT99), .ZN(new_n854));
  NOR4_X1   g429(.A1(new_n840), .A2(new_n843), .A3(new_n847), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n788), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n756), .A2(new_n856), .ZN(G311));
  XNOR2_X1  g432(.A(new_n754), .B(KEYINPUT36), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(new_n855), .A3(new_n788), .ZN(G150));
  NAND2_X1  g434(.A1(G80), .A2(G543), .ZN(new_n860));
  INV_X1    g435(.A(G67), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n506), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G651), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n551), .A2(G93), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n554), .B2(G55), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT76), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n574), .B1(new_n572), .B2(new_n573), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(new_n573), .A3(new_n572), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT38), .Z(new_n873));
  NAND4_X1  g448(.A1(new_n627), .A2(new_n632), .A3(new_n636), .A4(new_n640), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n874), .A2(new_n647), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n873), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n877));
  AOI21_X1  g452(.A(G860), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n877), .B2(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n867), .A2(G860), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT37), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(G145));
  XNOR2_X1  g457(.A(new_n818), .B(new_n495), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n765), .ZN(new_n884));
  INV_X1    g459(.A(new_n803), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n749), .B(new_n664), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n480), .A2(G142), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n482), .A2(G130), .ZN(new_n891));
  OR2_X1    g466(.A1(G106), .A2(G2105), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n892), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n889), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT100), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n888), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n888), .A2(new_n896), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(KEYINPUT101), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(KEYINPUT101), .B2(new_n898), .ZN(new_n900));
  XNOR2_X1  g475(.A(G160), .B(new_n486), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(new_n660), .Z(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n888), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n897), .B1(new_n904), .B2(new_n895), .ZN(new_n905));
  INV_X1    g480(.A(new_n902), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g484(.A(new_n872), .B(new_n649), .ZN(new_n910));
  NOR2_X1   g485(.A1(G299), .A2(KEYINPUT102), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(new_n587), .B2(new_n592), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n911), .A2(new_n874), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n874), .A2(KEYINPUT102), .A3(G299), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT103), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(G299), .A2(KEYINPUT102), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n591), .B1(new_n584), .B2(new_n586), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n912), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n641), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n874), .A2(KEYINPUT102), .A3(G299), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n917), .B1(new_n910), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n910), .A2(KEYINPUT103), .A3(new_n916), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G166), .B(G305), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(G290), .A2(G288), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n740), .A2(new_n730), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n931), .A2(KEYINPUT104), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n740), .A2(new_n730), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n738), .A2(G288), .A3(new_n739), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n932), .A2(KEYINPUT104), .A3(new_n933), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n930), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n941), .B(KEYINPUT42), .Z(new_n942));
  OR2_X1    g517(.A1(new_n929), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n929), .A2(new_n942), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(G868), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G868), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT105), .B1(new_n867), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n947), .B1(new_n945), .B2(new_n949), .ZN(G295));
  AOI21_X1  g525(.A(new_n947), .B1(new_n945), .B2(new_n949), .ZN(G331));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n537), .A2(new_n544), .A3(G171), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n526), .A2(KEYINPUT74), .A3(new_n536), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n543), .B1(new_n542), .B2(new_n535), .ZN(new_n955));
  AOI21_X1  g530(.A(G301), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n866), .B1(new_n566), .B2(new_n575), .ZN(new_n957));
  INV_X1    g532(.A(new_n871), .ZN(new_n958));
  OAI22_X1  g533(.A1(new_n953), .A2(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(G171), .B1(new_n537), .B2(new_n544), .ZN(new_n960));
  NAND3_X1  g535(.A1(G301), .A2(new_n954), .A3(new_n955), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n870), .A2(new_n960), .A3(new_n871), .A4(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n916), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n962), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n925), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n924), .A2(new_n925), .A3(new_n965), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n941), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G37), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n959), .A2(new_n962), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n941), .B(new_n963), .C1(new_n973), .C2(new_n926), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n971), .A2(KEYINPUT107), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n972), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT41), .B1(new_n914), .B2(new_n915), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(KEYINPUT106), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(new_n964), .A3(new_n966), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n941), .B1(new_n981), .B2(new_n963), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n976), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n975), .A2(new_n983), .A3(KEYINPUT43), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n964), .B1(new_n924), .B2(new_n925), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n941), .B1(new_n985), .B2(new_n963), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n977), .A2(new_n986), .A3(KEYINPUT43), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n952), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n971), .A2(new_n990), .A3(new_n972), .A4(new_n974), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT43), .B1(new_n977), .B2(new_n986), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n992), .A3(new_n952), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT108), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n959), .A2(new_n962), .B1(new_n925), .B2(new_n965), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n980), .A2(new_n997), .B1(new_n973), .B2(new_n916), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n972), .B(new_n974), .C1(new_n998), .C2(new_n941), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n990), .B1(new_n999), .B2(new_n976), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n987), .B1(new_n1000), .B2(new_n975), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n996), .B(new_n993), .C1(new_n1001), .C2(new_n952), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n995), .A2(new_n1002), .ZN(G397));
  OAI211_X1 g578(.A(new_n470), .B(G40), .C1(new_n475), .C2(new_n476), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT109), .B(G1384), .Z(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT45), .B1(new_n495), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1996), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n766), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT110), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1008), .ZN(new_n1012));
  INV_X1    g587(.A(G2067), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n818), .B(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT111), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(G1996), .B2(new_n765), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1011), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n749), .B(new_n752), .Z(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1008), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(G290), .B(G1986), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1012), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n730), .A2(G1976), .ZN(new_n1022));
  INV_X1    g597(.A(G1384), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n495), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n474), .A2(G2105), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT68), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n474), .A2(new_n471), .A3(G2105), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1024), .A2(G40), .A3(new_n470), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT113), .B1(new_n1029), .B2(G8), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n495), .A2(new_n1023), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT113), .B(G8), .C1(new_n1004), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1022), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n597), .A2(new_n605), .A3(G8), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n597), .A2(new_n605), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT112), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n495), .A2(new_n1043), .A3(KEYINPUT45), .A4(new_n1006), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT45), .B1(new_n495), .B2(new_n1023), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1004), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1971), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n495), .A2(new_n1049), .A3(new_n1023), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1049), .B1(new_n495), .B2(new_n1023), .ZN(new_n1052));
  NOR4_X1   g627(.A1(new_n1051), .A2(new_n1004), .A3(new_n1052), .A4(G2090), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1040), .B(G8), .C1(new_n1048), .C2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1022), .B(new_n1056), .C1(new_n1030), .C2(new_n1033), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT49), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT114), .B1(G305), .B2(G1981), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n614), .A2(new_n618), .A3(new_n1060), .A4(new_n722), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n722), .B1(new_n614), .B2(new_n618), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1058), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1064), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(KEYINPUT49), .A3(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1065), .B(new_n1067), .C1(new_n1030), .C2(new_n1033), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1035), .A2(new_n1054), .A3(new_n1057), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n954), .A2(new_n955), .A3(G8), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT126), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT51), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n1023), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT45), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1031), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n495), .A2(KEYINPUT118), .A3(KEYINPUT45), .A4(new_n1023), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1005), .A2(new_n1077), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1966), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1051), .A2(new_n1004), .A3(new_n1052), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1081), .A2(new_n1082), .B1(new_n1083), .B2(new_n779), .ZN(new_n1084));
  INV_X1    g659(.A(G8), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1074), .B(new_n1071), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1084), .A2(new_n1071), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1083), .A2(new_n779), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(G8), .B(new_n1073), .C1(new_n1091), .C2(G286), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1086), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n727), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1053), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT117), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(G8), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1040), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1045), .A2(new_n821), .A3(new_n1047), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1052), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1005), .A2(new_n1105), .A3(new_n1050), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1103), .A2(new_n1104), .B1(new_n782), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1104), .A2(G2078), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1047), .A2(new_n1080), .A3(new_n1077), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1111));
  NAND2_X1  g686(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n470), .A2(G40), .A3(new_n1025), .A4(new_n1108), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1007), .A2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1111), .A2(new_n1112), .B1(new_n1045), .B2(new_n1115), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1110), .A2(new_n1113), .B1(new_n1107), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1070), .A2(new_n1093), .A3(new_n1102), .A4(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1045), .A2(new_n1009), .A3(new_n1047), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT58), .B(G1341), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1029), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT59), .B1(new_n1122), .B2(new_n577), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1124), .B(new_n576), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT57), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1127), .A2(KEYINPUT57), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n919), .B2(new_n1129), .ZN(new_n1130));
  AND4_X1   g705(.A1(new_n587), .A2(new_n592), .A3(new_n1129), .A4(new_n1128), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT124), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(G299), .A2(new_n1127), .A3(KEYINPUT57), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n919), .A2(new_n1129), .A3(new_n1128), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G1956), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1106), .A2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1045), .A2(new_n1047), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(KEYINPUT61), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1139), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1144), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1126), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1004), .A2(new_n1031), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1013), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1153), .B(KEYINPUT60), .C1(new_n1083), .C2(G1348), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1154), .A2(KEYINPUT125), .A3(new_n874), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n874), .B1(new_n1154), .B2(KEYINPUT125), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1155), .A2(new_n1156), .B1(KEYINPUT125), .B2(new_n1154), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1153), .B1(new_n1083), .B2(G1348), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1151), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1143), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1158), .A2(new_n641), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1145), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1118), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(G2090), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1094), .A2(new_n727), .B1(new_n1083), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1085), .B1(new_n1168), .B2(new_n1097), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1040), .B1(new_n1169), .B2(new_n1099), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1110), .A2(G171), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1170), .A2(new_n1069), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1071), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1091), .B2(G8), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1087), .B1(new_n1174), .B2(new_n1074), .ZN(new_n1175));
  AOI21_X1  g750(.A(KEYINPUT62), .B1(new_n1175), .B2(new_n1092), .ZN(new_n1176));
  AND4_X1   g751(.A1(KEYINPUT62), .A2(new_n1086), .A3(new_n1092), .A4(new_n1088), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1172), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT127), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1172), .B(new_n1180), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1166), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1068), .A2(new_n1057), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT113), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1184), .B1(new_n1152), .B2(new_n1085), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1185), .A2(new_n1032), .B1(G1976), .B2(new_n730), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT52), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1183), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(G288), .A2(G1976), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT116), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1063), .B1(new_n1068), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT115), .ZN(new_n1195));
  OAI22_X1  g770(.A1(new_n1190), .A2(new_n1054), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1084), .A2(new_n1085), .A3(G286), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1102), .A2(new_n1189), .A3(new_n1054), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(KEYINPUT119), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT119), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1070), .A2(new_n1200), .A3(new_n1102), .A4(new_n1197), .ZN(new_n1201));
  XNOR2_X1  g776(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1199), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1101), .B1(new_n1168), .B2(new_n1085), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1197), .A2(new_n1204), .A3(KEYINPUT63), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1205), .A2(new_n1069), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1206), .A2(KEYINPUT121), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT121), .ZN(new_n1208));
  NOR3_X1   g783(.A1(new_n1205), .A2(new_n1069), .A3(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1196), .B1(new_n1203), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1182), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI211_X1 g788(.A(KEYINPUT122), .B(new_n1196), .C1(new_n1203), .C2(new_n1210), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1021), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1008), .B1(new_n1015), .B2(new_n766), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT46), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1012), .A2(new_n1009), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1219), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1220), .B(KEYINPUT47), .Z(new_n1221));
  NOR2_X1   g796(.A1(new_n749), .A2(new_n752), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1017), .A2(new_n1222), .ZN(new_n1223));
  OR2_X1    g798(.A1(new_n818), .A2(G2067), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1008), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NOR3_X1   g800(.A1(new_n1008), .A2(G1986), .A3(G290), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n1226), .B(KEYINPUT48), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1019), .A2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g803(.A1(new_n1221), .A2(new_n1225), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1215), .A2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g805(.A(new_n700), .B(G319), .C1(new_n684), .C2(new_n683), .ZN(new_n1232));
  NOR2_X1   g806(.A1(G229), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n992), .ZN(new_n1234));
  NAND3_X1  g808(.A1(new_n1233), .A2(new_n908), .A3(new_n1234), .ZN(G225));
  INV_X1    g809(.A(G225), .ZN(G308));
endmodule


