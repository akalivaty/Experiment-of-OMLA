

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U554 ( .A1(n633), .A2(n984), .ZN(n522) );
  XOR2_X1 U555 ( .A(KEYINPUT101), .B(n634), .Z(n523) );
  INV_X1 U556 ( .A(KEYINPUT103), .ZN(n641) );
  XNOR2_X1 U557 ( .A(n642), .B(n641), .ZN(n645) );
  INV_X1 U558 ( .A(KEYINPUT29), .ZN(n652) );
  XNOR2_X1 U559 ( .A(n653), .B(n652), .ZN(n654) );
  INV_X1 U560 ( .A(KEYINPUT107), .ZN(n671) );
  INV_X1 U561 ( .A(KEYINPUT12), .ZN(n622) );
  XNOR2_X1 U562 ( .A(n622), .B(KEYINPUT73), .ZN(n623) );
  XNOR2_X1 U563 ( .A(n624), .B(n623), .ZN(n626) );
  NOR2_X1 U564 ( .A1(G543), .A2(G651), .ZN(n791) );
  INV_X1 U565 ( .A(G2105), .ZN(n529) );
  XNOR2_X1 U566 ( .A(n525), .B(KEYINPUT65), .ZN(n907) );
  NOR2_X1 U567 ( .A1(n632), .A2(n631), .ZN(n984) );
  AND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n903) );
  NAND2_X1 U569 ( .A1(n903), .A2(G114), .ZN(n524) );
  XNOR2_X1 U570 ( .A(n524), .B(KEYINPUT92), .ZN(n527) );
  NAND2_X1 U571 ( .A1(n529), .A2(G2104), .ZN(n525) );
  NAND2_X1 U572 ( .A1(G102), .A2(n907), .ZN(n526) );
  NAND2_X1 U573 ( .A1(n527), .A2(n526), .ZN(n533) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XOR2_X1 U575 ( .A(KEYINPUT17), .B(n528), .Z(n908) );
  NAND2_X1 U576 ( .A1(G138), .A2(n908), .ZN(n531) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n529), .ZN(n904) );
  NAND2_X1 U578 ( .A1(G126), .A2(n904), .ZN(n530) );
  NAND2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U580 ( .A1(n533), .A2(n532), .ZN(G164) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n576) );
  NOR2_X1 U582 ( .A1(G651), .A2(n576), .ZN(n795) );
  NAND2_X1 U583 ( .A1(G48), .A2(n795), .ZN(n534) );
  XNOR2_X1 U584 ( .A(n534), .B(KEYINPUT84), .ZN(n543) );
  NAND2_X1 U585 ( .A1(G86), .A2(n791), .ZN(n537) );
  INV_X1 U586 ( .A(G651), .ZN(n538) );
  NOR2_X1 U587 ( .A1(G543), .A2(n538), .ZN(n535) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n535), .Z(n799) );
  NAND2_X1 U589 ( .A1(G61), .A2(n799), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n541) );
  NOR2_X1 U591 ( .A1(n576), .A2(n538), .ZN(n792) );
  NAND2_X1 U592 ( .A1(n792), .A2(G73), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT2), .B(n539), .Z(n540) );
  NOR2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(G305) );
  NAND2_X1 U596 ( .A1(G52), .A2(n795), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G64), .A2(n799), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n550) );
  NAND2_X1 U599 ( .A1(G90), .A2(n791), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G77), .A2(n792), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U602 ( .A(KEYINPUT9), .B(n548), .Z(n549) );
  NOR2_X1 U603 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U604 ( .A(KEYINPUT69), .B(n551), .Z(G171) );
  NAND2_X1 U605 ( .A1(n792), .A2(G76), .ZN(n552) );
  XNOR2_X1 U606 ( .A(KEYINPUT77), .B(n552), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n791), .A2(G89), .ZN(n553) );
  XOR2_X1 U608 ( .A(n553), .B(KEYINPUT4), .Z(n554) );
  NOR2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U610 ( .A(KEYINPUT5), .B(n556), .Z(n557) );
  XNOR2_X1 U611 ( .A(KEYINPUT78), .B(n557), .ZN(n563) );
  XNOR2_X1 U612 ( .A(KEYINPUT79), .B(KEYINPUT6), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G51), .A2(n795), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G63), .A2(n799), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U616 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U618 ( .A(n564), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U619 ( .A1(G88), .A2(n791), .ZN(n565) );
  XNOR2_X1 U620 ( .A(n565), .B(KEYINPUT86), .ZN(n568) );
  NAND2_X1 U621 ( .A1(G50), .A2(n795), .ZN(n566) );
  XOR2_X1 U622 ( .A(KEYINPUT85), .B(n566), .Z(n567) );
  NAND2_X1 U623 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U624 ( .A1(G75), .A2(n792), .ZN(n570) );
  NAND2_X1 U625 ( .A1(G62), .A2(n799), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U627 ( .A1(n572), .A2(n571), .ZN(G166) );
  XNOR2_X1 U628 ( .A(KEYINPUT93), .B(G166), .ZN(G303) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G49), .A2(n795), .ZN(n574) );
  NAND2_X1 U631 ( .A1(G74), .A2(G651), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U633 ( .A1(n799), .A2(n575), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n576), .A2(G87), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n578), .A2(n577), .ZN(G288) );
  NAND2_X1 U636 ( .A1(G47), .A2(n795), .ZN(n580) );
  NAND2_X1 U637 ( .A1(G60), .A2(n799), .ZN(n579) );
  NAND2_X1 U638 ( .A1(n580), .A2(n579), .ZN(n586) );
  NAND2_X1 U639 ( .A1(n791), .A2(G85), .ZN(n581) );
  XNOR2_X1 U640 ( .A(n581), .B(KEYINPUT66), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G72), .A2(n792), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U643 ( .A(KEYINPUT67), .B(n584), .Z(n585) );
  NOR2_X1 U644 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U645 ( .A(KEYINPUT68), .B(n587), .Z(G290) );
  NAND2_X1 U646 ( .A1(n908), .A2(G137), .ZN(n761) );
  INV_X1 U647 ( .A(n761), .ZN(n592) );
  INV_X1 U648 ( .A(G40), .ZN(n590) );
  NAND2_X1 U649 ( .A1(G113), .A2(n903), .ZN(n589) );
  NAND2_X1 U650 ( .A1(G125), .A2(n904), .ZN(n588) );
  NAND2_X1 U651 ( .A1(n589), .A2(n588), .ZN(n764) );
  OR2_X1 U652 ( .A1(n590), .A2(n764), .ZN(n591) );
  NOR2_X1 U653 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U654 ( .A1(G101), .A2(n907), .ZN(n593) );
  XOR2_X1 U655 ( .A(n593), .B(KEYINPUT23), .Z(n762) );
  NAND2_X1 U656 ( .A1(n594), .A2(n762), .ZN(n709) );
  XNOR2_X1 U657 ( .A(n709), .B(KEYINPUT99), .ZN(n595) );
  NOR2_X1 U658 ( .A1(G164), .A2(G1384), .ZN(n710) );
  NAND2_X1 U659 ( .A1(n595), .A2(n710), .ZN(n656) );
  NAND2_X1 U660 ( .A1(G8), .A2(n656), .ZN(n703) );
  NOR2_X1 U661 ( .A1(G1981), .A2(G305), .ZN(n596) );
  XOR2_X1 U662 ( .A(n596), .B(KEYINPUT24), .Z(n597) );
  NOR2_X1 U663 ( .A1(n703), .A2(n597), .ZN(n708) );
  NOR2_X1 U664 ( .A1(G1966), .A2(n703), .ZN(n670) );
  INV_X1 U665 ( .A(n656), .ZN(n620) );
  BUF_X1 U666 ( .A(n620), .Z(n607) );
  INV_X1 U667 ( .A(G1961), .ZN(n992) );
  NAND2_X1 U668 ( .A1(n656), .A2(n992), .ZN(n600) );
  XNOR2_X1 U669 ( .A(G2078), .B(KEYINPUT100), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n598), .B(KEYINPUT25), .ZN(n954) );
  NAND2_X1 U671 ( .A1(n607), .A2(n954), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n662) );
  NAND2_X1 U673 ( .A1(n662), .A2(G171), .ZN(n655) );
  NAND2_X1 U674 ( .A1(G53), .A2(n795), .ZN(n602) );
  NAND2_X1 U675 ( .A1(G65), .A2(n799), .ZN(n601) );
  NAND2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G91), .A2(n791), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G78), .A2(n792), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n771) );
  NAND2_X1 U681 ( .A1(n607), .A2(G2072), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n608), .B(KEYINPUT27), .ZN(n610) );
  AND2_X1 U683 ( .A1(G1956), .A2(n656), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n648) );
  NAND2_X1 U685 ( .A1(n771), .A2(n648), .ZN(n647) );
  NAND2_X1 U686 ( .A1(G66), .A2(n799), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G92), .A2(n791), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G79), .A2(n792), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G54), .A2(n795), .ZN(n613) );
  XNOR2_X1 U691 ( .A(KEYINPUT75), .B(n613), .ZN(n614) );
  NOR2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n618), .B(KEYINPUT15), .ZN(n619) );
  XOR2_X1 U695 ( .A(KEYINPUT76), .B(n619), .Z(n979) );
  NAND2_X1 U696 ( .A1(n620), .A2(G1996), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n621), .B(KEYINPUT26), .ZN(n633) );
  NAND2_X1 U698 ( .A1(G81), .A2(n791), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G68), .A2(n792), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT13), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G43), .A2(n795), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n799), .A2(G56), .ZN(n630) );
  XOR2_X1 U705 ( .A(KEYINPUT14), .B(n630), .Z(n631) );
  NAND2_X1 U706 ( .A1(G1341), .A2(n656), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n522), .A2(n523), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n635), .B(KEYINPUT64), .ZN(n643) );
  OR2_X1 U709 ( .A1(n979), .A2(n643), .ZN(n640) );
  INV_X1 U710 ( .A(G2067), .ZN(n865) );
  NOR2_X1 U711 ( .A1(n656), .A2(n865), .ZN(n636) );
  XOR2_X1 U712 ( .A(n636), .B(KEYINPUT102), .Z(n638) );
  NAND2_X1 U713 ( .A1(n656), .A2(G1348), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n979), .A2(n643), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n651) );
  NOR2_X1 U719 ( .A1(n771), .A2(n648), .ZN(n649) );
  XOR2_X1 U720 ( .A(n649), .B(KEYINPUT28), .Z(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n668) );
  NOR2_X1 U723 ( .A1(G2084), .A2(n656), .ZN(n673) );
  NOR2_X1 U724 ( .A1(n673), .A2(n670), .ZN(n657) );
  NAND2_X1 U725 ( .A1(G8), .A2(n657), .ZN(n658) );
  XNOR2_X1 U726 ( .A(KEYINPUT105), .B(n658), .ZN(n660) );
  XOR2_X1 U727 ( .A(KEYINPUT30), .B(KEYINPUT104), .Z(n659) );
  XNOR2_X1 U728 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U729 ( .A1(G168), .A2(n661), .ZN(n664) );
  NOR2_X1 U730 ( .A1(G171), .A2(n662), .ZN(n663) );
  NOR2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n666) );
  XOR2_X1 U732 ( .A(KEYINPUT31), .B(KEYINPUT106), .Z(n665) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n680) );
  INV_X1 U735 ( .A(n680), .ZN(n669) );
  NOR2_X2 U736 ( .A1(n670), .A2(n669), .ZN(n672) );
  XNOR2_X1 U737 ( .A(n672), .B(n671), .ZN(n675) );
  NAND2_X1 U738 ( .A1(G8), .A2(n673), .ZN(n674) );
  NAND2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n686) );
  NOR2_X1 U740 ( .A1(G1971), .A2(n703), .ZN(n676) );
  XNOR2_X1 U741 ( .A(n676), .B(KEYINPUT108), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n656), .A2(G2090), .ZN(n677) );
  NOR2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n679), .A2(G303), .ZN(n682) );
  NAND2_X1 U745 ( .A1(G286), .A2(n680), .ZN(n681) );
  NAND2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U747 ( .A1(G8), .A2(n683), .ZN(n684) );
  XNOR2_X1 U748 ( .A(KEYINPUT32), .B(n684), .ZN(n685) );
  NAND2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n702) );
  NOR2_X1 U750 ( .A1(G1976), .A2(G288), .ZN(n692) );
  NOR2_X1 U751 ( .A1(G1971), .A2(G303), .ZN(n687) );
  NOR2_X1 U752 ( .A1(n692), .A2(n687), .ZN(n982) );
  INV_X1 U753 ( .A(KEYINPUT33), .ZN(n688) );
  AND2_X1 U754 ( .A1(n982), .A2(n688), .ZN(n689) );
  NAND2_X1 U755 ( .A1(n702), .A2(n689), .ZN(n699) );
  INV_X1 U756 ( .A(n703), .ZN(n690) );
  NAND2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n988) );
  AND2_X1 U758 ( .A1(n690), .A2(n988), .ZN(n691) );
  OR2_X1 U759 ( .A1(KEYINPUT33), .A2(n691), .ZN(n695) );
  NAND2_X1 U760 ( .A1(n692), .A2(KEYINPUT33), .ZN(n693) );
  OR2_X1 U761 ( .A1(n693), .A2(n703), .ZN(n694) );
  NAND2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n697) );
  XOR2_X1 U763 ( .A(G1981), .B(G305), .Z(n976) );
  INV_X1 U764 ( .A(n976), .ZN(n696) );
  NOR2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n706) );
  NOR2_X1 U767 ( .A1(G2090), .A2(G303), .ZN(n700) );
  NAND2_X1 U768 ( .A1(G8), .A2(n700), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n742) );
  NOR2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n756) );
  XOR2_X1 U774 ( .A(n865), .B(KEYINPUT37), .Z(n711) );
  XNOR2_X1 U775 ( .A(n711), .B(KEYINPUT94), .ZN(n754) );
  NAND2_X1 U776 ( .A1(G104), .A2(n907), .ZN(n713) );
  NAND2_X1 U777 ( .A1(G140), .A2(n908), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U779 ( .A(KEYINPUT34), .B(n714), .ZN(n720) );
  NAND2_X1 U780 ( .A1(n903), .A2(G116), .ZN(n715) );
  XOR2_X1 U781 ( .A(KEYINPUT95), .B(n715), .Z(n717) );
  NAND2_X1 U782 ( .A1(n904), .A2(G128), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U784 ( .A(KEYINPUT35), .B(n718), .Z(n719) );
  NOR2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U786 ( .A(KEYINPUT36), .B(n721), .ZN(n900) );
  NOR2_X1 U787 ( .A1(n754), .A2(n900), .ZN(n932) );
  NAND2_X1 U788 ( .A1(n756), .A2(n932), .ZN(n752) );
  NAND2_X1 U789 ( .A1(G107), .A2(n903), .ZN(n723) );
  NAND2_X1 U790 ( .A1(G119), .A2(n904), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U792 ( .A(KEYINPUT96), .B(n724), .ZN(n728) );
  NAND2_X1 U793 ( .A1(G95), .A2(n907), .ZN(n726) );
  NAND2_X1 U794 ( .A1(G131), .A2(n908), .ZN(n725) );
  NAND2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n914) );
  INV_X1 U797 ( .A(G1991), .ZN(n850) );
  NOR2_X1 U798 ( .A1(n914), .A2(n850), .ZN(n739) );
  XOR2_X1 U799 ( .A(KEYINPUT38), .B(KEYINPUT98), .Z(n730) );
  NAND2_X1 U800 ( .A1(G105), .A2(n907), .ZN(n729) );
  XNOR2_X1 U801 ( .A(n730), .B(n729), .ZN(n735) );
  NAND2_X1 U802 ( .A1(G117), .A2(n903), .ZN(n732) );
  NAND2_X1 U803 ( .A1(G129), .A2(n904), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U805 ( .A(KEYINPUT97), .B(n733), .Z(n734) );
  NOR2_X1 U806 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U807 ( .A1(n908), .A2(G141), .ZN(n736) );
  NAND2_X1 U808 ( .A1(n737), .A2(n736), .ZN(n899) );
  AND2_X1 U809 ( .A1(n899), .A2(G1996), .ZN(n738) );
  NOR2_X1 U810 ( .A1(n739), .A2(n738), .ZN(n929) );
  INV_X1 U811 ( .A(n929), .ZN(n740) );
  NAND2_X1 U812 ( .A1(n740), .A2(n756), .ZN(n745) );
  NAND2_X1 U813 ( .A1(n752), .A2(n745), .ZN(n741) );
  NOR2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n744) );
  XNOR2_X1 U815 ( .A(G1986), .B(G290), .ZN(n994) );
  NAND2_X1 U816 ( .A1(n994), .A2(n756), .ZN(n743) );
  NAND2_X1 U817 ( .A1(n744), .A2(n743), .ZN(n759) );
  NOR2_X1 U818 ( .A1(G1996), .A2(n899), .ZN(n945) );
  INV_X1 U819 ( .A(n745), .ZN(n748) );
  NOR2_X1 U820 ( .A1(G1986), .A2(G290), .ZN(n746) );
  AND2_X1 U821 ( .A1(n850), .A2(n914), .ZN(n928) );
  NOR2_X1 U822 ( .A1(n746), .A2(n928), .ZN(n747) );
  NOR2_X1 U823 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U824 ( .A(KEYINPUT109), .B(n749), .Z(n750) );
  NOR2_X1 U825 ( .A1(n945), .A2(n750), .ZN(n751) );
  XNOR2_X1 U826 ( .A(n751), .B(KEYINPUT39), .ZN(n753) );
  NAND2_X1 U827 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U828 ( .A1(n754), .A2(n900), .ZN(n942) );
  NAND2_X1 U829 ( .A1(n755), .A2(n942), .ZN(n757) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U831 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U832 ( .A(n760), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U833 ( .A(G171), .ZN(G301) );
  AND2_X1 U834 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U835 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U836 ( .A1(n764), .A2(n763), .ZN(G160) );
  INV_X1 U837 ( .A(G132), .ZN(G219) );
  INV_X1 U838 ( .A(G82), .ZN(G220) );
  XOR2_X1 U839 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n766) );
  NAND2_X1 U840 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U841 ( .A(n766), .B(n765), .ZN(G223) );
  XOR2_X1 U842 ( .A(G223), .B(KEYINPUT72), .Z(n832) );
  NAND2_X1 U843 ( .A1(n832), .A2(G567), .ZN(n767) );
  XOR2_X1 U844 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  NAND2_X1 U845 ( .A1(n984), .A2(G860), .ZN(G153) );
  NAND2_X1 U846 ( .A1(G301), .A2(G868), .ZN(n768) );
  XNOR2_X1 U847 ( .A(n768), .B(KEYINPUT74), .ZN(n770) );
  INV_X1 U848 ( .A(G868), .ZN(n804) );
  NAND2_X1 U849 ( .A1(n804), .A2(n979), .ZN(n769) );
  NAND2_X1 U850 ( .A1(n770), .A2(n769), .ZN(G284) );
  INV_X1 U851 ( .A(n771), .ZN(G299) );
  XOR2_X1 U852 ( .A(KEYINPUT80), .B(G868), .Z(n772) );
  NOR2_X1 U853 ( .A1(G286), .A2(n772), .ZN(n775) );
  NOR2_X1 U854 ( .A1(G868), .A2(G299), .ZN(n773) );
  XOR2_X1 U855 ( .A(KEYINPUT81), .B(n773), .Z(n774) );
  NOR2_X1 U856 ( .A1(n775), .A2(n774), .ZN(G297) );
  INV_X1 U857 ( .A(G860), .ZN(n776) );
  NAND2_X1 U858 ( .A1(n776), .A2(G559), .ZN(n777) );
  INV_X1 U859 ( .A(n979), .ZN(n873) );
  NAND2_X1 U860 ( .A1(n777), .A2(n873), .ZN(n778) );
  XNOR2_X1 U861 ( .A(n778), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U862 ( .A1(G868), .A2(n873), .ZN(n779) );
  NOR2_X1 U863 ( .A1(G559), .A2(n779), .ZN(n781) );
  AND2_X1 U864 ( .A1(n804), .A2(n984), .ZN(n780) );
  NOR2_X1 U865 ( .A1(n781), .A2(n780), .ZN(G282) );
  NAND2_X1 U866 ( .A1(G123), .A2(n904), .ZN(n782) );
  XNOR2_X1 U867 ( .A(n782), .B(KEYINPUT18), .ZN(n785) );
  NAND2_X1 U868 ( .A1(G111), .A2(n903), .ZN(n783) );
  XNOR2_X1 U869 ( .A(n783), .B(KEYINPUT82), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U871 ( .A1(G99), .A2(n907), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G135), .A2(n908), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n927) );
  XNOR2_X1 U875 ( .A(n927), .B(G2096), .ZN(n790) );
  INV_X1 U876 ( .A(G2100), .ZN(n863) );
  NAND2_X1 U877 ( .A1(n790), .A2(n863), .ZN(G156) );
  NAND2_X1 U878 ( .A1(G93), .A2(n791), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G80), .A2(n792), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U881 ( .A1(G55), .A2(n795), .ZN(n796) );
  XNOR2_X1 U882 ( .A(KEYINPUT83), .B(n796), .ZN(n797) );
  NOR2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U884 ( .A1(n799), .A2(G67), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n801), .A2(n800), .ZN(n806) );
  NAND2_X1 U886 ( .A1(n873), .A2(G559), .ZN(n802) );
  XOR2_X1 U887 ( .A(n984), .B(n802), .Z(n813) );
  NOR2_X1 U888 ( .A1(G860), .A2(n813), .ZN(n803) );
  XOR2_X1 U889 ( .A(n806), .B(n803), .Z(G145) );
  NAND2_X1 U890 ( .A1(n804), .A2(n806), .ZN(n805) );
  XNOR2_X1 U891 ( .A(n805), .B(KEYINPUT88), .ZN(n816) );
  XOR2_X1 U892 ( .A(G299), .B(G166), .Z(n812) );
  XNOR2_X1 U893 ( .A(G290), .B(G305), .ZN(n807) );
  XNOR2_X1 U894 ( .A(n807), .B(n806), .ZN(n808) );
  XNOR2_X1 U895 ( .A(KEYINPUT87), .B(n808), .ZN(n810) );
  XNOR2_X1 U896 ( .A(G288), .B(KEYINPUT19), .ZN(n809) );
  XNOR2_X1 U897 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U898 ( .A(n812), .B(n811), .ZN(n872) );
  XNOR2_X1 U899 ( .A(n872), .B(n813), .ZN(n814) );
  NAND2_X1 U900 ( .A1(G868), .A2(n814), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n816), .A2(n815), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2078), .A2(G2084), .ZN(n817) );
  XNOR2_X1 U903 ( .A(n817), .B(KEYINPUT89), .ZN(n818) );
  XNOR2_X1 U904 ( .A(KEYINPUT20), .B(n818), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n819), .A2(G2090), .ZN(n820) );
  XNOR2_X1 U906 ( .A(KEYINPUT21), .B(n820), .ZN(n821) );
  NAND2_X1 U907 ( .A1(n821), .A2(G2072), .ZN(G158) );
  XOR2_X1 U908 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U909 ( .A(KEYINPUT90), .B(G44), .ZN(n822) );
  XNOR2_X1 U910 ( .A(n822), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U911 ( .A1(G108), .A2(G120), .ZN(n823) );
  NOR2_X1 U912 ( .A1(G237), .A2(n823), .ZN(n824) );
  NAND2_X1 U913 ( .A1(G69), .A2(n824), .ZN(n837) );
  NAND2_X1 U914 ( .A1(n837), .A2(G567), .ZN(n829) );
  NOR2_X1 U915 ( .A1(G220), .A2(G219), .ZN(n825) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n825), .Z(n826) );
  NOR2_X1 U917 ( .A1(G218), .A2(n826), .ZN(n827) );
  NAND2_X1 U918 ( .A1(G96), .A2(n827), .ZN(n836) );
  NAND2_X1 U919 ( .A1(n836), .A2(G2106), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(n926) );
  NAND2_X1 U921 ( .A1(G661), .A2(G483), .ZN(n830) );
  XOR2_X1 U922 ( .A(KEYINPUT91), .B(n830), .Z(n831) );
  NOR2_X1 U923 ( .A1(n926), .A2(n831), .ZN(n835) );
  NAND2_X1 U924 ( .A1(n835), .A2(G36), .ZN(G176) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U927 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G108), .ZN(G238) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n837), .A2(n836), .ZN(n838) );
  XOR2_X1 U936 ( .A(n838), .B(KEYINPUT112), .Z(G261) );
  INV_X1 U937 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U938 ( .A(KEYINPUT110), .B(G2454), .ZN(n847) );
  XNOR2_X1 U939 ( .A(G2430), .B(G2435), .ZN(n845) );
  XOR2_X1 U940 ( .A(G2451), .B(G2427), .Z(n840) );
  XNOR2_X1 U941 ( .A(G2438), .B(G2446), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U943 ( .A(n841), .B(G2443), .Z(n843) );
  XNOR2_X1 U944 ( .A(G1341), .B(G1348), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  NAND2_X1 U948 ( .A1(n848), .A2(G14), .ZN(n849) );
  XNOR2_X1 U949 ( .A(KEYINPUT111), .B(n849), .ZN(G401) );
  XNOR2_X1 U950 ( .A(G1996), .B(KEYINPUT114), .ZN(n860) );
  XOR2_X1 U951 ( .A(G1976), .B(G1956), .Z(n852) );
  XOR2_X1 U952 ( .A(n850), .B(G1961), .Z(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U954 ( .A(G1981), .B(G1971), .Z(n854) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1966), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U957 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U958 ( .A(G2474), .B(KEYINPUT41), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(G229) );
  XOR2_X1 U961 ( .A(KEYINPUT113), .B(G2090), .Z(n862) );
  XNOR2_X1 U962 ( .A(G2084), .B(G2078), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n867) );
  XOR2_X1 U965 ( .A(n865), .B(G2072), .Z(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U967 ( .A(G2096), .B(KEYINPUT43), .Z(n869) );
  XNOR2_X1 U968 ( .A(G2678), .B(KEYINPUT42), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U970 ( .A(n871), .B(n870), .Z(G227) );
  XOR2_X1 U971 ( .A(n872), .B(G286), .Z(n875) );
  XOR2_X1 U972 ( .A(n873), .B(n984), .Z(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U974 ( .A(n876), .B(G301), .Z(n877) );
  NOR2_X1 U975 ( .A1(G37), .A2(n877), .ZN(G397) );
  NAND2_X1 U976 ( .A1(G124), .A2(n904), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n878), .B(KEYINPUT44), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G112), .A2(n903), .ZN(n879) );
  XOR2_X1 U979 ( .A(KEYINPUT115), .B(n879), .Z(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G100), .A2(n907), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G136), .A2(n908), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  NOR2_X1 U984 ( .A1(n885), .A2(n884), .ZN(G162) );
  XOR2_X1 U985 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n887) );
  XNOR2_X1 U986 ( .A(n927), .B(KEYINPUT48), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n898) );
  NAND2_X1 U988 ( .A1(G103), .A2(n907), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G139), .A2(n908), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G115), .A2(n903), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G127), .A2(n904), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U996 ( .A(KEYINPUT117), .B(n895), .Z(n935) );
  XNOR2_X1 U997 ( .A(G164), .B(n935), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n896), .B(G162), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U1000 ( .A(n900), .B(n899), .Z(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n918) );
  NAND2_X1 U1002 ( .A1(G118), .A2(n903), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(G130), .A2(n904), .ZN(n905) );
  NAND2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(G106), .A2(n907), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n908), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1008 ( .A(n911), .B(KEYINPUT45), .Z(n912) );
  NOR2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n915) );
  XOR2_X1 U1010 ( .A(n915), .B(n914), .Z(n916) );
  XNOR2_X1 U1011 ( .A(G160), .B(n916), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n919), .ZN(n920) );
  XNOR2_X1 U1014 ( .A(KEYINPUT118), .B(n920), .ZN(G395) );
  OR2_X1 U1015 ( .A1(n926), .A2(G401), .ZN(n923) );
  NOR2_X1 U1016 ( .A1(G229), .A2(G227), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(G397), .A2(G395), .ZN(n924) );
  NAND2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(n926), .ZN(G319) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n934) );
  XNOR2_X1 U1024 ( .A(G160), .B(G2084), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1027 ( .A1(n934), .A2(n933), .ZN(n941) );
  XNOR2_X1 U1028 ( .A(G2072), .B(n935), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(G164), .B(G2078), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n938), .Z(n939) );
  XNOR2_X1 U1032 ( .A(KEYINPUT119), .B(n939), .ZN(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n943), .A2(n942), .ZN(n948) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(n946), .B(KEYINPUT51), .ZN(n947) );
  NOR2_X1 U1038 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1039 ( .A(KEYINPUT52), .B(n949), .ZN(n950) );
  INV_X1 U1040 ( .A(KEYINPUT55), .ZN(n972) );
  NAND2_X1 U1041 ( .A1(n950), .A2(n972), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n951), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1043 ( .A(G29), .B(KEYINPUT123), .ZN(n974) );
  XOR2_X1 U1044 ( .A(G1996), .B(G32), .Z(n953) );
  XOR2_X1 U1045 ( .A(G2067), .B(G26), .Z(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1047 ( .A(n954), .B(G27), .Z(n955) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n963) );
  XOR2_X1 U1049 ( .A(G1991), .B(G25), .Z(n957) );
  NAND2_X1 U1050 ( .A1(n957), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(n958), .B(KEYINPUT120), .ZN(n961) );
  XOR2_X1 U1052 ( .A(G2072), .B(KEYINPUT121), .Z(n959) );
  XNOR2_X1 U1053 ( .A(G33), .B(n959), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n964), .ZN(n968) );
  XOR2_X1 U1057 ( .A(KEYINPUT122), .B(G34), .Z(n966) );
  XNOR2_X1 U1058 ( .A(G2084), .B(KEYINPUT54), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n966), .B(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(G35), .B(G2090), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1063 ( .A(n972), .B(n971), .Z(n973) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n975), .ZN(n1029) );
  INV_X1 U1066 ( .A(G16), .ZN(n1025) );
  XOR2_X1 U1067 ( .A(n1025), .B(KEYINPUT56), .Z(n1001) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(KEYINPUT57), .B(n978), .ZN(n999) );
  XOR2_X1 U1071 ( .A(n979), .B(G1348), .Z(n981) );
  NAND2_X1 U1072 ( .A1(G1971), .A2(G303), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n991) );
  XOR2_X1 U1074 ( .A(G299), .B(G1956), .Z(n983) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n987) );
  XOR2_X1 U1076 ( .A(G1341), .B(n984), .Z(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT124), .B(n985), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n996) );
  XOR2_X1 U1081 ( .A(n992), .B(G301), .Z(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(KEYINPUT125), .B(n997), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1027) );
  XOR2_X1 U1087 ( .A(G5), .B(G1961), .Z(n1015) );
  XOR2_X1 U1088 ( .A(G1966), .B(G21), .Z(n1012) );
  XNOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(n1002), .B(G4), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G1956), .B(G20), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(KEYINPUT126), .B(G1981), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G6), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(n1010), .B(KEYINPUT60), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(KEYINPUT127), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1022) );
  XNOR2_X1 U1102 ( .A(G1971), .B(G22), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G23), .B(G1976), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(G1986), .B(G24), .Z(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT58), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1032), .ZN(G150) );
  INV_X1 U1115 ( .A(G150), .ZN(G311) );
endmodule

