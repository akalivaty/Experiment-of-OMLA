//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  AND2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OR3_X1    g0007(.A1(new_n207), .A2(KEYINPUT65), .A3(G13), .ZN(new_n208));
  OAI21_X1  g0008(.A(KEYINPUT65), .B1(new_n207), .B2(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(G58), .A2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n211), .A2(new_n212), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(new_n212), .B2(new_n211), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT67), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n207), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n221), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT69), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  INV_X1    g0044(.A(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT68), .B(G50), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G77), .ZN(new_n255));
  OR2_X1    g0055(.A1(KEYINPUT72), .A2(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT72), .A2(G1698), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n256), .A2(new_n251), .A3(new_n253), .A4(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G222), .ZN(new_n259));
  INV_X1    g0059(.A(G223), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G1698), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n255), .B1(new_n258), .B2(new_n259), .C1(new_n260), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT73), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n264), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n274), .A2(new_n275), .A3(new_n268), .ZN(new_n276));
  XOR2_X1   g0076(.A(KEYINPUT70), .B(G226), .Z(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G169), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n213), .ZN(new_n283));
  INV_X1    g0083(.A(G20), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n203), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G150), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(G33), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n283), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G13), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n292), .A2(new_n284), .A3(G1), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n283), .ZN(new_n294));
  INV_X1    g0094(.A(G50), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(new_n271), .B2(G20), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n294), .A2(new_n296), .B1(new_n295), .B2(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n278), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n267), .B2(new_n268), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n281), .A2(new_n298), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT76), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n300), .B2(G190), .ZN(new_n305));
  INV_X1    g0105(.A(G41), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n214), .B1(new_n250), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n265), .B2(new_n266), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  NOR4_X1   g0109(.A1(new_n308), .A2(KEYINPUT76), .A3(new_n309), .A4(new_n299), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT9), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT75), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n291), .B2(new_n297), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n291), .A2(new_n313), .A3(new_n297), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n316), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n318), .A2(KEYINPUT9), .A3(new_n314), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n317), .A2(new_n319), .B1(new_n320), .B2(new_n300), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n311), .A2(new_n321), .A3(KEYINPUT10), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT10), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n269), .A2(G190), .A3(new_n278), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT76), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n300), .A2(new_n304), .A3(G190), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT9), .B1(new_n318), .B2(new_n314), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n315), .A2(new_n312), .A3(new_n316), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n328), .A2(new_n329), .B1(new_n279), .B2(G200), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n323), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n303), .B1(new_n322), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT77), .ZN(new_n334));
  INV_X1    g0134(.A(G226), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n258), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n256), .A2(new_n257), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n337), .A2(KEYINPUT77), .A3(G226), .A4(new_n261), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G97), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n262), .B2(new_n232), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n268), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n273), .B1(new_n276), .B2(G238), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n342), .A2(new_n343), .B1(KEYINPUT78), .B2(KEYINPUT13), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n342), .A2(KEYINPUT78), .A3(KEYINPUT13), .A4(new_n343), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n309), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n341), .B1(new_n338), .B2(new_n336), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n343), .B1(new_n348), .B2(new_n307), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n343), .B(KEYINPUT13), .C1(new_n348), .C2(new_n307), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G200), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n294), .A2(KEYINPUT74), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT74), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n293), .B2(new_n283), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n271), .A2(G20), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n354), .A2(new_n356), .A3(G68), .A4(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G68), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n286), .A2(G50), .B1(G20), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n204), .B2(new_n289), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n283), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT11), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n293), .A2(new_n359), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT12), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(KEYINPUT11), .A3(new_n283), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n358), .A2(new_n364), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT79), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n353), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n347), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n369), .ZN(new_n372));
  INV_X1    g0172(.A(new_n346), .ZN(new_n373));
  OAI21_X1  g0173(.A(G179), .B1(new_n373), .B2(new_n344), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n351), .A2(G169), .A3(new_n352), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT14), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n351), .A2(new_n377), .A3(G169), .A4(new_n352), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n371), .B1(new_n372), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n288), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n286), .B1(G20), .B2(G77), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n289), .B2(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(new_n283), .B1(new_n204), .B2(new_n293), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n354), .A2(new_n356), .A3(G77), .A4(new_n357), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n254), .A2(G107), .ZN(new_n388));
  INV_X1    g0188(.A(G238), .ZN(new_n389));
  OAI221_X1 g0189(.A(new_n388), .B1(new_n258), .B2(new_n232), .C1(new_n389), .C2(new_n262), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n268), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n273), .B1(new_n276), .B2(G244), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n387), .B1(G190), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n320), .B2(new_n393), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n393), .A2(new_n301), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n387), .B1(new_n393), .B2(G169), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n333), .A2(new_n380), .A3(new_n395), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n294), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n381), .A2(new_n357), .ZN(new_n402));
  INV_X1    g0202(.A(new_n293), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n401), .A2(new_n402), .B1(new_n403), .B2(new_n381), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n283), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT81), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT81), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT7), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n284), .B2(new_n254), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n407), .B(G20), .C1(new_n251), .C2(new_n253), .ZN(new_n413));
  OAI21_X1  g0213(.A(G68), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n245), .A2(new_n359), .ZN(new_n415));
  OAI21_X1  g0215(.A(G20), .B1(new_n415), .B2(new_n216), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n286), .A2(G159), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n406), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT81), .B(KEYINPUT7), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n261), .A2(new_n423), .A3(G20), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n252), .A2(G33), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT80), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT80), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n251), .A2(new_n253), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n284), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n424), .B1(new_n430), .B2(new_n407), .ZN(new_n431));
  OAI211_X1 g0231(.A(KEYINPUT16), .B(new_n419), .C1(new_n431), .C2(new_n359), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n422), .A2(KEYINPUT82), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT82), .B1(new_n422), .B2(new_n432), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n405), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n273), .B1(new_n276), .B2(G232), .ZN(new_n436));
  INV_X1    g0236(.A(G87), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n258), .A2(new_n260), .B1(new_n250), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT83), .B1(new_n262), .B2(new_n335), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT83), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n261), .A2(new_n440), .A3(G226), .A4(G1698), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n438), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n436), .B1(new_n442), .B2(new_n307), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G169), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n436), .B(G179), .C1(new_n442), .C2(new_n307), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n435), .A2(KEYINPUT18), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT84), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n435), .A2(KEYINPUT84), .A3(KEYINPUT18), .A4(new_n446), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT18), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT82), .ZN(new_n452));
  INV_X1    g0252(.A(new_n432), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n423), .B1(new_n261), .B2(G20), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n284), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n418), .B1(new_n456), .B2(G68), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n283), .B1(new_n457), .B2(KEYINPUT16), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n452), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n422), .A2(KEYINPUT82), .A3(new_n432), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n404), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n446), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n451), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n449), .A2(new_n450), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n443), .A2(new_n320), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n436), .B(new_n309), .C1(new_n442), .C2(new_n307), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n405), .B(new_n467), .C1(new_n433), .C2(new_n434), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT85), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(KEYINPUT17), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n459), .A2(new_n460), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n472), .A2(new_n405), .A3(new_n467), .A4(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n464), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n400), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT21), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n271), .B2(G33), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n354), .A2(new_n356), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n293), .A2(new_n479), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n282), .A2(new_n213), .B1(G20), .B2(new_n479), .ZN(new_n483));
  AOI21_X1  g0283(.A(G20), .B1(G33), .B2(G283), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n250), .A2(G97), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT90), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n484), .B2(new_n485), .ZN(new_n489));
  OAI211_X1 g0289(.A(KEYINPUT20), .B(new_n483), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n484), .A2(new_n485), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT90), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n487), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT20), .B1(new_n494), .B2(new_n483), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n481), .B(new_n482), .C1(new_n491), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G169), .ZN(new_n497));
  INV_X1    g0297(.A(G45), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(G1), .ZN(new_n499));
  XNOR2_X1  g0299(.A(KEYINPUT5), .B(G41), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n268), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G270), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n307), .A2(G274), .A3(new_n499), .A4(new_n500), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n251), .A2(new_n253), .A3(G257), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n256), .A2(new_n257), .ZN(new_n506));
  INV_X1    g0306(.A(G303), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n505), .A2(new_n506), .B1(new_n261), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n251), .A2(new_n253), .A3(G264), .A4(G1698), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n268), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT89), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n254), .A2(G303), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n514), .B(new_n509), .C1(new_n506), .C2(new_n505), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(KEYINPUT89), .A3(new_n268), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n504), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n478), .B1(new_n497), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n496), .ZN(new_n519));
  INV_X1    g0319(.A(new_n504), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n515), .A2(KEYINPUT89), .A3(new_n268), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT89), .B1(new_n515), .B2(new_n268), .ZN(new_n522));
  OAI211_X1 g0322(.A(G190), .B(new_n520), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n519), .B(new_n523), .C1(new_n320), .C2(new_n517), .ZN(new_n524));
  AOI211_X1 g0324(.A(new_n301), .B(new_n504), .C1(new_n513), .C2(new_n516), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n496), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n527), .A2(new_n496), .A3(KEYINPUT21), .A4(G169), .ZN(new_n528));
  AND4_X1   g0328(.A1(new_n518), .A2(new_n524), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n251), .A2(new_n253), .A3(G257), .A4(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G294), .ZN(new_n531));
  INV_X1    g0331(.A(G250), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n531), .C1(new_n258), .C2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n268), .B1(G264), .B2(new_n501), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n534), .A2(KEYINPUT91), .A3(new_n309), .A4(new_n503), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT91), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n268), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n501), .A2(G264), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n503), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n536), .B1(new_n539), .B2(new_n320), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(G190), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n251), .A2(new_n253), .A3(new_n284), .A4(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT22), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n261), .A2(new_n545), .A3(new_n284), .A4(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(G20), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT23), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n284), .B2(G107), .ZN(new_n551));
  INV_X1    g0351(.A(G107), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(KEYINPUT23), .A3(G20), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n549), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT24), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n547), .A2(new_n557), .A3(new_n554), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n406), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n403), .A2(G107), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n560), .B(KEYINPUT25), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n294), .B1(G1), .B2(new_n250), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n552), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n542), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(G97), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n293), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n562), .B2(new_n566), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n456), .A2(G107), .ZN(new_n569));
  NAND2_X1  g0369(.A1(KEYINPUT6), .A2(G97), .ZN(new_n570));
  OR3_X1    g0370(.A1(new_n570), .A2(KEYINPUT87), .A3(G107), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT87), .B1(new_n570), .B2(G107), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n566), .A2(new_n552), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n571), .B(new_n572), .C1(new_n575), .C2(KEYINPUT6), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G20), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n286), .A2(G77), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT86), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n569), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n568), .B1(new_n580), .B2(new_n283), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  INV_X1    g0383(.A(G244), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n258), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n337), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G283), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n268), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n500), .A2(new_n499), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(G257), .A3(new_n307), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n503), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n280), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n593), .B1(new_n589), .B2(new_n268), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n301), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n582), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n597), .A2(new_n309), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n597), .A2(G200), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n581), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n565), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n251), .A2(new_n253), .A3(G244), .A4(G1698), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n548), .B(new_n604), .C1(new_n258), .C2(new_n389), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT88), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n337), .A2(G238), .A3(new_n261), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n608), .A2(KEYINPUT88), .A3(new_n548), .A4(new_n604), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n268), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n307), .A2(G274), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n499), .A2(new_n532), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n613), .A2(new_n499), .B1(new_n307), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n611), .A2(G190), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n261), .A2(new_n284), .A3(G68), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT19), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n284), .B1(new_n340), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n574), .A2(new_n437), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n618), .B1(new_n289), .B2(new_n566), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n283), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n383), .A2(new_n293), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n294), .B(G87), .C1(G1), .C2(new_n250), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n307), .B1(new_n607), .B2(new_n609), .ZN(new_n629));
  INV_X1    g0429(.A(new_n615), .ZN(new_n630));
  OAI21_X1  g0430(.A(G200), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n616), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n611), .A2(new_n301), .A3(new_n615), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n280), .B1(new_n629), .B2(new_n630), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n624), .B(new_n625), .C1(new_n383), .C2(new_n562), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n539), .A2(new_n280), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n534), .A2(new_n301), .A3(new_n503), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n637), .B(new_n638), .C1(new_n559), .C2(new_n563), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n632), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n477), .A2(new_n529), .A3(new_n603), .A4(new_n640), .ZN(G372));
  NOR3_X1   g0441(.A1(new_n461), .A2(new_n451), .A3(new_n462), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT18), .B1(new_n435), .B2(new_n446), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n379), .A2(new_n372), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n371), .B2(new_n399), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n644), .B1(new_n646), .B2(new_n475), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT10), .B1(new_n311), .B2(new_n321), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n327), .A2(new_n323), .A3(new_n330), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n303), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n477), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n627), .A2(KEYINPUT92), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT92), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n624), .A2(new_n656), .A3(new_n625), .A4(new_n626), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n616), .A2(new_n658), .A3(new_n631), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n636), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n597), .A2(G169), .ZN(new_n662));
  AOI211_X1 g0462(.A(G179), .B(new_n593), .C1(new_n589), .C2(new_n268), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n662), .A2(new_n581), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n660), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n632), .A3(new_n636), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT26), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n565), .A2(new_n599), .A3(new_n602), .A4(new_n659), .ZN(new_n669));
  AND4_X1   g0469(.A1(new_n518), .A2(new_n639), .A3(new_n526), .A4(new_n528), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n636), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n653), .B1(new_n654), .B2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n518), .A2(new_n526), .A3(new_n528), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n271), .A2(new_n284), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n519), .A2(new_n681), .ZN(new_n682));
  MUX2_X1   g0482(.A(new_n529), .B(new_n674), .S(new_n682), .Z(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n680), .B1(new_n559), .B2(new_n563), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n565), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n639), .ZN(new_n689));
  INV_X1    g0489(.A(new_n639), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n681), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n674), .A2(new_n681), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n691), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n210), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n574), .A2(new_n437), .A3(new_n479), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n701), .A2(new_n271), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n218), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(new_n701), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT28), .Z(new_n706));
  INV_X1    g0506(.A(KEYINPUT96), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n666), .A2(new_n661), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n664), .A2(new_n659), .A3(new_n636), .A4(KEYINPUT26), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n602), .A2(new_n599), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n518), .A2(new_n639), .A3(new_n526), .A4(new_n528), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(new_n565), .A4(new_n659), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n713), .A3(new_n636), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT95), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n714), .A2(new_n715), .A3(new_n681), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n714), .B2(new_n681), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n707), .B(KEYINPUT29), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n708), .A2(new_n709), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n681), .B1(new_n720), .B2(new_n671), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT95), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n714), .A2(new_n715), .A3(new_n681), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n719), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n672), .A2(new_n680), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT96), .B1(new_n725), .B2(KEYINPUT29), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n718), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT94), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n527), .B1(new_n629), .B2(new_n630), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n595), .A2(new_n301), .A3(new_n539), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n611), .A2(new_n597), .A3(new_n534), .A4(new_n615), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n517), .A2(G179), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n539), .A2(new_n301), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n597), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n611), .A2(new_n615), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(KEYINPUT94), .A3(new_n527), .A4(new_n739), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n590), .A2(new_n594), .A3(new_n534), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n629), .A2(new_n630), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n525), .A2(new_n741), .A3(KEYINPUT30), .A4(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n732), .A2(new_n736), .A3(new_n740), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n680), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n603), .A2(new_n529), .A3(new_n640), .A4(new_n681), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n738), .A2(new_n527), .A3(new_n739), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n736), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n681), .A2(new_n746), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(KEYINPUT93), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n747), .A2(new_n748), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n728), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n706), .B1(new_n760), .B2(G1), .ZN(G364));
  NOR2_X1   g0561(.A1(new_n292), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n271), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n701), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n686), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G330), .B2(new_n683), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n765), .A2(KEYINPUT97), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(KEYINPUT97), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n213), .B1(G20), .B2(new_n280), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n284), .A2(new_n301), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n309), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n773), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n777), .A2(new_n309), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n261), .B1(new_n776), .B2(new_n295), .C1(new_n245), .C2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n782), .A2(KEYINPUT98), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(KEYINPUT98), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n780), .B1(new_n786), .B2(G77), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n774), .A2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n359), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n284), .A2(G179), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n437), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n791), .A2(new_n309), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n552), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n301), .A2(new_n320), .A3(G190), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n566), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n790), .A2(new_n793), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n791), .A2(new_n309), .A3(new_n320), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT99), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G159), .ZN(new_n806));
  OAI21_X1  g0606(.A(KEYINPUT32), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OR3_X1    g0607(.A1(new_n805), .A2(KEYINPUT32), .A3(new_n806), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n787), .A2(new_n800), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n794), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G317), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n812), .A2(KEYINPUT33), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(KEYINPUT33), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n789), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n811), .B(new_n815), .C1(G326), .C2(new_n775), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n781), .A2(G311), .ZN(new_n817));
  INV_X1    g0617(.A(G322), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n779), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G294), .B2(new_n797), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n254), .B1(new_n792), .B2(new_n507), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT100), .ZN(new_n822));
  INV_X1    g0622(.A(new_n805), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G329), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n816), .A2(new_n820), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n772), .B1(new_n809), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(G13), .A2(G33), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(G20), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n771), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n700), .A2(new_n254), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n831), .A2(G355), .B1(new_n479), .B2(new_n700), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n248), .A2(new_n498), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n427), .A2(new_n429), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n700), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(G45), .B2(new_n218), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n832), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n770), .B(new_n826), .C1(new_n830), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n829), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n683), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n767), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  NAND2_X1  g0642(.A1(new_n387), .A2(new_n680), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n395), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n399), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n398), .A2(new_n681), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n848), .B(new_n681), .C1(new_n671), .C2(new_n668), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n847), .B1(new_n672), .B2(new_n680), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n765), .B1(new_n758), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n758), .B2(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(new_n770), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n771), .A2(new_n827), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT101), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n794), .A2(new_n437), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n789), .A2(new_n810), .B1(new_n776), .B2(new_n507), .ZN(new_n858));
  INV_X1    g0658(.A(new_n792), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n857), .B(new_n858), .C1(G107), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(G294), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n254), .B1(new_n566), .B2(new_n798), .C1(new_n779), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n785), .A2(new_n479), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n862), .B(new_n863), .C1(G311), .C2(new_n823), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n778), .A2(G143), .B1(new_n775), .B2(G137), .ZN(new_n865));
  INV_X1    g0665(.A(G150), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n865), .B1(new_n866), .B2(new_n789), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n786), .B2(G159), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n868), .A2(KEYINPUT34), .ZN(new_n869));
  INV_X1    g0669(.A(new_n834), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(G50), .B2(new_n859), .ZN(new_n871));
  INV_X1    g0671(.A(new_n794), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n872), .A2(G68), .B1(new_n797), .B2(G58), .ZN(new_n873));
  INV_X1    g0673(.A(G132), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n871), .B(new_n873), .C1(new_n874), .C2(new_n805), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n868), .B2(KEYINPUT34), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n860), .A2(new_n864), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n854), .B1(G77), .B2(new_n856), .C1(new_n877), .C2(new_n772), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT102), .Z(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n828), .B2(new_n848), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n853), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(G384));
  AOI211_X1 g0682(.A(new_n479), .B(new_n215), .C1(new_n576), .C2(KEYINPUT35), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(KEYINPUT35), .B2(new_n576), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT36), .ZN(new_n885));
  OAI21_X1  g0685(.A(G77), .B1(new_n245), .B2(new_n359), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n218), .A2(new_n886), .B1(G50), .B2(new_n359), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(G1), .A3(new_n292), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT103), .Z(new_n890));
  AND3_X1   g0690(.A1(new_n744), .A2(KEYINPUT106), .A3(new_n680), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT106), .B1(new_n744), .B2(new_n680), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT31), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n744), .A2(new_n751), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n748), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n654), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT107), .Z(new_n898));
  OAI21_X1  g0698(.A(new_n419), .B1(new_n431), .B2(new_n359), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n421), .A2(KEYINPUT104), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n283), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n405), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n678), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n476), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n903), .B1(new_n446), .B2(new_n904), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n468), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n435), .A2(new_n446), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n435), .A2(new_n904), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n468), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n905), .B1(new_n464), .B2(new_n475), .ZN(new_n918));
  INV_X1    g0718(.A(new_n915), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n371), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n372), .A2(new_n680), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n645), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n372), .B(new_n680), .C1(new_n371), .C2(new_n379), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n847), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT40), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(new_n893), .C2(new_n895), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n921), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n926), .B1(new_n893), .B2(new_n895), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n911), .A2(new_n912), .A3(new_n468), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT37), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n914), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n463), .A2(new_n447), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n912), .B1(new_n475), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT105), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI211_X1 g0738(.A(KEYINPUT105), .B(new_n912), .C1(new_n475), .C2(new_n935), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n917), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n931), .B1(new_n940), .B2(new_n916), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n930), .B1(new_n941), .B2(new_n927), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n898), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n685), .B1(new_n898), .B2(new_n942), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n924), .A2(new_n925), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n849), .B2(new_n846), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n921), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n644), .A2(new_n678), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT39), .ZN(new_n951));
  INV_X1    g0751(.A(new_n912), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n471), .A2(new_n474), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n644), .B2(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n954), .A2(KEYINPUT105), .B1(new_n914), .B2(new_n933), .ZN(new_n955));
  INV_X1    g0755(.A(new_n939), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT38), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n918), .A2(new_n919), .A3(new_n917), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n951), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n916), .A2(new_n920), .A3(KEYINPUT39), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n645), .A2(new_n680), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n949), .B(new_n950), .C1(new_n961), .C2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n652), .B1(new_n727), .B2(new_n477), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n945), .A2(new_n966), .B1(new_n271), .B2(new_n762), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n945), .A2(new_n966), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n890), .B1(new_n967), .B2(new_n968), .ZN(G367));
  INV_X1    g0769(.A(new_n835), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n238), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n830), .B1(new_n210), .B2(new_n383), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n854), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n794), .A2(new_n204), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n254), .B(new_n974), .C1(G150), .C2(new_n778), .ZN(new_n975));
  INV_X1    g0775(.A(G137), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n975), .B1(new_n976), .B2(new_n805), .C1(new_n785), .C2(new_n295), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n798), .A2(new_n359), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G143), .B2(new_n775), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n245), .B2(new_n792), .C1(new_n806), .C2(new_n789), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n834), .B1(G303), .B2(new_n778), .ZN(new_n981));
  XOR2_X1   g0781(.A(KEYINPUT110), .B(G317), .Z(new_n982));
  OAI221_X1 g0782(.A(new_n981), .B1(new_n805), .B2(new_n982), .C1(new_n785), .C2(new_n810), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT109), .B1(new_n792), .B2(new_n479), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n788), .A2(G294), .B1(new_n775), .B2(G311), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n872), .A2(G97), .B1(new_n797), .B2(G107), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n985), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n977), .A2(new_n980), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT47), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n973), .B1(new_n991), .B2(new_n771), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n658), .A2(new_n681), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n660), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n636), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n992), .B1(new_n996), .B2(new_n839), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n711), .B1(new_n581), .B2(new_n681), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n664), .A2(new_n680), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n696), .A2(new_n691), .A3(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT45), .Z(new_n1002));
  INV_X1    g0802(.A(new_n1000), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT44), .B1(new_n697), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n697), .A2(KEYINPUT44), .A3(new_n1003), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n694), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n692), .B(new_n695), .Z(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(new_n686), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n760), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n701), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n764), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT108), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n693), .A2(new_n1000), .A3(new_n674), .A4(new_n681), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT42), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n599), .B1(new_n998), .B2(new_n639), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1016), .A2(KEYINPUT42), .B1(new_n681), .B2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1017), .A2(new_n1019), .B1(KEYINPUT43), .B2(new_n996), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1020), .B(new_n1021), .Z(new_n1022));
  NOR2_X1   g0822(.A1(new_n694), .A2(new_n1003), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1014), .A2(new_n1015), .A3(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1006), .B(new_n694), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n759), .A2(new_n1010), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n759), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n763), .B1(new_n1029), .B2(new_n1012), .ZN(new_n1030));
  AOI21_X1  g0830(.A(KEYINPUT108), .B1(new_n1030), .B2(new_n1024), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n997), .B1(new_n1026), .B2(new_n1031), .ZN(G387));
  INV_X1    g0832(.A(new_n1028), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n759), .A2(new_n1010), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n701), .A3(new_n1034), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n235), .A2(new_n498), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1036), .A2(new_n835), .B1(new_n702), .B2(new_n831), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n381), .B2(new_n295), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n288), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n498), .B1(new_n359), .B2(new_n204), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n702), .A4(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1037), .A2(new_n1042), .B1(G107), .B2(new_n210), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n770), .B1(new_n1043), .B2(new_n830), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n823), .A2(G326), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n870), .B1(new_n479), .B2(new_n794), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n982), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n778), .A2(new_n1047), .B1(new_n788), .B2(G311), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n818), .B2(new_n776), .C1(new_n785), .C2(new_n507), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n859), .A2(G294), .B1(new_n797), .B2(G283), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1045), .B(new_n1046), .C1(new_n1055), .C2(KEYINPUT49), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(KEYINPUT49), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n798), .A2(new_n383), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G50), .B2(new_n778), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT111), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n805), .A2(new_n866), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n806), .A2(new_n776), .B1(new_n789), .B2(new_n288), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n834), .B1(new_n782), .B2(new_n359), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n204), .A2(new_n792), .B1(new_n794), .B2(new_n566), .ZN(new_n1064));
  NOR4_X1   g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1056), .A2(new_n1057), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1044), .B1(new_n693), .B2(new_n839), .C1(new_n1066), .C2(new_n772), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1035), .B(new_n1067), .C1(new_n763), .C2(new_n1010), .ZN(G393));
  NAND2_X1  g0868(.A1(new_n1008), .A2(new_n1033), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n701), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT112), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1069), .A2(new_n1070), .A3(KEYINPUT112), .A4(new_n701), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n970), .A2(new_n242), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n830), .B1(new_n210), .B2(new_n566), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n854), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n870), .B(new_n857), .C1(new_n786), .C2(new_n381), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n789), .A2(new_n295), .B1(new_n792), .B2(new_n359), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G77), .B2(new_n797), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n823), .A2(G143), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n778), .A2(G159), .B1(new_n775), .B2(G150), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT51), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n778), .A2(G311), .B1(new_n775), .B2(G317), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n789), .A2(new_n507), .B1(new_n792), .B2(new_n810), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G116), .B2(new_n797), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n261), .B(new_n795), .C1(G294), .C2(new_n781), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(new_n818), .C2(new_n805), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1083), .A2(new_n1085), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1078), .B1(new_n1092), .B2(new_n771), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n1000), .B2(new_n839), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1008), .B2(new_n763), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1075), .A2(new_n1096), .ZN(G390));
  OAI211_X1 g0897(.A(new_n926), .B(G330), .C1(new_n893), .C2(new_n895), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT113), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n948), .A2(new_n962), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n959), .B2(new_n960), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n940), .A2(new_n916), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n722), .A2(new_n723), .A3(new_n846), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n845), .A3(new_n946), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n963), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1101), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n948), .A2(new_n962), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT39), .B1(new_n940), .B2(new_n916), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n916), .A2(new_n920), .A3(KEYINPUT39), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n757), .A2(new_n848), .A3(new_n946), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(KEYINPUT113), .B2(new_n1098), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1116), .A3(new_n1107), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1109), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1118), .A2(new_n763), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n961), .A2(new_n827), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n854), .B1(new_n381), .B2(new_n856), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n261), .B1(new_n779), .B2(new_n874), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G159), .B2(new_n797), .ZN(new_n1123));
  INV_X1    g0923(.A(G125), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1123), .B1(new_n1124), .B2(new_n805), .C1(new_n785), .C2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n792), .A2(new_n866), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT53), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n788), .A2(G137), .B1(new_n872), .B2(G50), .ZN(new_n1129));
  INV_X1    g0929(.A(G128), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1128), .B(new_n1129), .C1(new_n1130), .C2(new_n776), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n261), .B(new_n793), .C1(G116), .C2(new_n778), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n861), .B2(new_n805), .C1(new_n785), .C2(new_n566), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n872), .A2(G68), .B1(new_n797), .B2(G77), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n789), .B2(new_n552), .C1(new_n810), .C2(new_n776), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1126), .A2(new_n1131), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1121), .B1(new_n1136), .B2(new_n771), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1119), .B1(new_n1120), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n701), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1105), .A2(new_n845), .ZN(new_n1140));
  OAI211_X1 g0940(.A(G330), .B(new_n848), .C1(new_n893), .C2(new_n895), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n947), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1114), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n756), .A2(G330), .A3(new_n848), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n947), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1098), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n849), .A2(new_n846), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n477), .B(G330), .C1(new_n893), .C2(new_n895), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n965), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1139), .B1(new_n1118), .B2(new_n1151), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n965), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1109), .A2(new_n1153), .A3(new_n1117), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(KEYINPUT114), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT114), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1138), .B1(new_n1156), .B2(new_n1158), .ZN(G378));
  AOI21_X1  g0959(.A(new_n678), .B1(new_n315), .B2(new_n316), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n650), .B2(new_n303), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n303), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1163), .B(new_n1160), .C1(new_n648), .C2(new_n649), .ZN(new_n1164));
  OAI21_X1  g0964(.A(KEYINPUT119), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n332), .A2(new_n1160), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT119), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n650), .A2(new_n303), .A3(new_n1161), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  XOR2_X1   g0969(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1170));
  AND3_X1   g0970(.A1(new_n1165), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n942), .A2(G330), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n942), .B2(G330), .ZN(new_n1175));
  OAI21_X1  g0975(.A(KEYINPUT120), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n949), .A2(new_n950), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1177), .B1(new_n1178), .B2(new_n962), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(KEYINPUT120), .B(new_n964), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n764), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n552), .A2(new_n779), .B1(new_n782), .B2(new_n383), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n978), .B(new_n1184), .C1(G283), .C2(new_n823), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n775), .A2(G116), .B1(new_n859), .B2(G77), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n788), .A2(G97), .B1(new_n872), .B2(G58), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n834), .A2(G41), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT58), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n295), .B1(G33), .B2(G41), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n779), .A2(new_n1130), .B1(new_n792), .B2(new_n1125), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT115), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n781), .A2(G137), .B1(new_n775), .B2(G125), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n788), .A2(G132), .B1(G150), .B2(new_n797), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT59), .Z(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT116), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n823), .A2(G124), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G33), .B(G41), .C1(new_n872), .C2(G159), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1197), .A2(KEYINPUT116), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1190), .B1(new_n1188), .B2(new_n1191), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT117), .Z(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n771), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT118), .Z(new_n1206));
  AOI211_X1 g1006(.A(new_n764), .B(new_n701), .C1(new_n295), .C2(new_n855), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n1173), .C2(new_n828), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1183), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1179), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n928), .B1(new_n916), .B2(new_n920), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n931), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n957), .B2(new_n958), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1213), .B1(new_n1215), .B2(KEYINPUT40), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1212), .B1(new_n1216), .B2(new_n685), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n942), .A2(new_n1173), .A3(G330), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n964), .A3(new_n1218), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1211), .A2(KEYINPUT57), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT121), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n965), .A2(new_n1150), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1154), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1221), .B1(new_n1154), .B2(new_n1223), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT122), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1220), .B(KEYINPUT122), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1113), .A2(new_n1116), .A3(new_n1107), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1100), .B1(new_n1113), .B2(new_n1107), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1151), .ZN(new_n1233));
  OAI21_X1  g1033(.A(KEYINPUT121), .B1(new_n1233), .B2(new_n1222), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1154), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1234), .A2(new_n1235), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n701), .B1(new_n1236), .B2(KEYINPUT57), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1210), .B1(new_n1230), .B2(new_n1237), .ZN(G375));
  NOR2_X1   g1038(.A1(new_n1223), .A2(new_n1149), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1239), .A2(new_n1012), .A3(new_n1153), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT123), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n947), .A2(new_n827), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n854), .B1(G68), .B2(new_n856), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n789), .A2(new_n479), .B1(new_n776), .B2(new_n861), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1058), .B(new_n1244), .C1(G97), .C2(new_n859), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n786), .A2(G107), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n823), .A2(G303), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n261), .B(new_n974), .C1(G283), .C2(new_n778), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n778), .A2(G137), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n789), .B2(new_n1125), .C1(new_n874), .C2(new_n776), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT124), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n823), .A2(G128), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n859), .A2(G159), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n872), .A2(G58), .B1(new_n797), .B2(G50), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n870), .B1(G150), .B2(new_n781), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1249), .B1(new_n1252), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1243), .B1(new_n1258), .B2(new_n771), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1149), .A2(new_n764), .B1(new_n1242), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1241), .A2(new_n1260), .ZN(G381));
  INV_X1    g1061(.A(G390), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1260), .A4(new_n1241), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1138), .A2(new_n1155), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OR4_X1    g1066(.A1(G387), .A2(new_n1264), .A3(G375), .A4(new_n1266), .ZN(G407));
  INV_X1    g1067(.A(G375), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n679), .A2(G213), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1265), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G407), .A2(G213), .A3(new_n1271), .ZN(G409));
  OAI211_X1 g1072(.A(G378), .B(new_n1210), .C1(new_n1230), .C2(new_n1237), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1236), .A2(new_n1013), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1211), .A2(new_n1219), .A3(new_n764), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1208), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1265), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(KEYINPUT125), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1151), .A2(KEYINPUT60), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1139), .B1(new_n1239), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1239), .B2(new_n1281), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(G384), .A3(new_n1260), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G384), .B1(new_n1283), .B2(new_n1260), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1280), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1286), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(KEYINPUT126), .A3(new_n1284), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1273), .A2(new_n1291), .A3(new_n1277), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1279), .A2(new_n1269), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1279), .A2(new_n1269), .A3(new_n1292), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1270), .A2(G2897), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1287), .A2(new_n1289), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1288), .A2(new_n1284), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(G2897), .A3(new_n1270), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1296), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G393), .B(new_n841), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1015), .B1(new_n1014), .B2(new_n1025), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1030), .A2(new_n1024), .A3(KEYINPUT108), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(G390), .A3(new_n997), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G390), .B1(new_n1308), .B2(new_n997), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1305), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT61), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G387), .A2(new_n1262), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(new_n1304), .A3(new_n1309), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1278), .A2(new_n1290), .A3(KEYINPUT63), .A4(new_n1269), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1317), .B2(KEYINPUT127), .ZN(new_n1318));
  OR2_X1    g1118(.A1(new_n1317), .A2(KEYINPUT127), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1295), .A2(new_n1303), .A3(new_n1318), .A4(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1270), .B1(new_n1273), .B2(new_n1277), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1313), .B1(new_n1321), .B2(new_n1301), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1293), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1321), .A2(KEYINPUT62), .A3(new_n1290), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1322), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1312), .A2(new_n1315), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1320), .B1(new_n1326), .B2(new_n1328), .ZN(G405));
  OAI21_X1  g1129(.A(new_n1273), .B1(new_n1268), .B2(new_n1266), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1290), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1331), .B1(new_n1332), .B2(new_n1330), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(new_n1327), .ZN(G402));
endmodule


