

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(n369), .B(n368), .ZN(n532) );
  INV_X1 U325 ( .A(KEYINPUT64), .ZN(n412) );
  INV_X1 U326 ( .A(KEYINPUT96), .ZN(n456) );
  XNOR2_X1 U327 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n343) );
  XNOR2_X1 U328 ( .A(n344), .B(n343), .ZN(n358) );
  INV_X1 U329 ( .A(n418), .ZN(n419) );
  INV_X1 U330 ( .A(KEYINPUT24), .ZN(n426) );
  INV_X1 U331 ( .A(KEYINPUT48), .ZN(n368) );
  XNOR2_X1 U332 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U333 ( .A(n320), .B(n430), .ZN(n321) );
  XNOR2_X1 U334 ( .A(n429), .B(n428), .ZN(n433) );
  XNOR2_X1 U335 ( .A(n322), .B(n321), .ZN(n325) );
  XNOR2_X1 U336 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U337 ( .A(n413), .B(n412), .ZN(n573) );
  XNOR2_X1 U338 ( .A(n459), .B(n458), .ZN(n574) );
  XOR2_X1 U339 ( .A(n581), .B(KEYINPUT41), .Z(n552) );
  XNOR2_X1 U340 ( .A(KEYINPUT38), .B(n480), .ZN(n504) );
  XNOR2_X1 U341 ( .A(n452), .B(n451), .ZN(n453) );
  INV_X1 U342 ( .A(G36GAT), .ZN(n481) );
  XNOR2_X1 U343 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n482), .B(n481), .ZN(G1329GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n293) );
  XNOR2_X1 U346 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n292) );
  XNOR2_X1 U347 ( .A(n293), .B(n292), .ZN(n307) );
  XOR2_X1 U348 ( .A(G99GAT), .B(G85GAT), .Z(n323) );
  XOR2_X1 U349 ( .A(G50GAT), .B(G162GAT), .Z(n418) );
  XOR2_X1 U350 ( .A(n323), .B(n418), .Z(n295) );
  NAND2_X1 U351 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U352 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U353 ( .A(KEYINPUT9), .B(G106GAT), .Z(n297) );
  XNOR2_X1 U354 ( .A(G134GAT), .B(G92GAT), .ZN(n296) );
  XOR2_X1 U355 ( .A(n297), .B(n296), .Z(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n305) );
  XOR2_X1 U357 ( .A(KEYINPUT69), .B(KEYINPUT8), .Z(n301) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(G29GAT), .ZN(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U360 ( .A(KEYINPUT7), .B(n302), .ZN(n342) );
  INV_X1 U361 ( .A(n342), .ZN(n303) );
  XOR2_X1 U362 ( .A(G36GAT), .B(G190GAT), .Z(n382) );
  XNOR2_X1 U363 ( .A(n303), .B(n382), .ZN(n304) );
  XNOR2_X1 U364 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U365 ( .A(n307), .B(n306), .Z(n558) );
  INV_X1 U366 ( .A(n558), .ZN(n546) );
  XOR2_X1 U367 ( .A(G78GAT), .B(KEYINPUT13), .Z(n309) );
  XNOR2_X1 U368 ( .A(G71GAT), .B(G64GAT), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n309), .B(n308), .ZN(n311) );
  INV_X1 U370 ( .A(G57GAT), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n348) );
  XOR2_X1 U372 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n313) );
  XNOR2_X1 U373 ( .A(G120GAT), .B(KEYINPUT74), .ZN(n312) );
  XNOR2_X1 U374 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n348), .B(n314), .ZN(n322) );
  XOR2_X1 U376 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n316) );
  NAND2_X1 U377 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U378 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n317), .B(KEYINPUT33), .ZN(n320) );
  XOR2_X1 U380 ( .A(KEYINPUT72), .B(G106GAT), .Z(n319) );
  XNOR2_X1 U381 ( .A(G148GAT), .B(G204GAT), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n430) );
  XOR2_X1 U383 ( .A(G176GAT), .B(G92GAT), .Z(n383) );
  XNOR2_X1 U384 ( .A(n383), .B(n323), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n581) );
  XOR2_X1 U386 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n327) );
  XNOR2_X1 U387 ( .A(KEYINPUT70), .B(KEYINPUT67), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n340) );
  XOR2_X1 U389 ( .A(G8GAT), .B(G197GAT), .Z(n329) );
  XNOR2_X1 U390 ( .A(G50GAT), .B(G36GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U392 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n331) );
  XNOR2_X1 U393 ( .A(G169GAT), .B(G22GAT), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U395 ( .A(n333), .B(n332), .Z(n338) );
  XOR2_X1 U396 ( .A(G15GAT), .B(G1GAT), .Z(n350) );
  XOR2_X1 U397 ( .A(G141GAT), .B(G113GAT), .Z(n335) );
  NAND2_X1 U398 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n350), .B(n336), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U402 ( .A(n340), .B(n339), .Z(n341) );
  XOR2_X1 U403 ( .A(n342), .B(n341), .Z(n550) );
  INV_X1 U404 ( .A(n550), .ZN(n575) );
  NOR2_X1 U405 ( .A1(n552), .A2(n575), .ZN(n344) );
  XOR2_X1 U406 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n346) );
  XNOR2_X1 U407 ( .A(KEYINPUT12), .B(KEYINPUT75), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n357) );
  XNOR2_X1 U410 ( .A(G8GAT), .B(G183GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n349), .B(G211GAT), .ZN(n381) );
  XOR2_X1 U412 ( .A(n381), .B(n350), .Z(n352) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U415 ( .A(n353), .B(KEYINPUT76), .Z(n355) );
  XOR2_X1 U416 ( .A(G22GAT), .B(G155GAT), .Z(n417) );
  XNOR2_X1 U417 ( .A(G127GAT), .B(n417), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n357), .B(n356), .ZN(n585) );
  XNOR2_X1 U420 ( .A(n585), .B(KEYINPUT114), .ZN(n571) );
  NAND2_X1 U421 ( .A1(n358), .A2(n571), .ZN(n359) );
  NOR2_X1 U422 ( .A1(n558), .A2(n359), .ZN(n360) );
  XNOR2_X1 U423 ( .A(KEYINPUT47), .B(n360), .ZN(n367) );
  INV_X1 U424 ( .A(n581), .ZN(n479) );
  INV_X1 U425 ( .A(KEYINPUT36), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n361), .B(n558), .ZN(n588) );
  NOR2_X1 U427 ( .A1(n588), .A2(n585), .ZN(n362) );
  XOR2_X1 U428 ( .A(KEYINPUT45), .B(n362), .Z(n363) );
  NOR2_X1 U429 ( .A1(n479), .A2(n363), .ZN(n364) );
  XNOR2_X1 U430 ( .A(KEYINPUT116), .B(n364), .ZN(n365) );
  NAND2_X1 U431 ( .A1(n365), .A2(n575), .ZN(n366) );
  NAND2_X1 U432 ( .A1(n367), .A2(n366), .ZN(n369) );
  XOR2_X1 U433 ( .A(KEYINPUT79), .B(KEYINPUT17), .Z(n371) );
  XNOR2_X1 U434 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U436 ( .A(G169GAT), .B(n372), .Z(n449) );
  XOR2_X1 U437 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n374) );
  XNOR2_X1 U438 ( .A(G204GAT), .B(G64GAT), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n380) );
  XOR2_X1 U440 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n376) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(G218GAT), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n425) );
  XOR2_X1 U443 ( .A(n425), .B(KEYINPUT91), .Z(n378) );
  NAND2_X1 U444 ( .A1(G226GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n382), .B(n381), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U450 ( .A(n449), .B(n387), .Z(n522) );
  NOR2_X1 U451 ( .A1(n532), .A2(n522), .ZN(n388) );
  XNOR2_X1 U452 ( .A(KEYINPUT54), .B(n388), .ZN(n411) );
  XOR2_X1 U453 ( .A(KEYINPUT86), .B(G155GAT), .Z(n390) );
  XNOR2_X1 U454 ( .A(G1GAT), .B(G148GAT), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U456 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n392) );
  XNOR2_X1 U457 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U459 ( .A(n394), .B(n393), .Z(n401) );
  XOR2_X1 U460 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n396) );
  XNOR2_X1 U461 ( .A(G141GAT), .B(KEYINPUT84), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n431) );
  XOR2_X1 U463 ( .A(G85GAT), .B(n431), .Z(n398) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(G57GAT), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U466 ( .A(G162GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U468 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n403) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U471 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U472 ( .A(G120GAT), .B(G134GAT), .Z(n407) );
  XNOR2_X1 U473 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n406) );
  XNOR2_X1 U474 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U475 ( .A(G113GAT), .B(n408), .Z(n435) );
  XNOR2_X1 U476 ( .A(n435), .B(KEYINPUT87), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n520) );
  NAND2_X1 U478 ( .A1(n411), .A2(n520), .ZN(n413) );
  XOR2_X1 U479 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n415) );
  XNOR2_X1 U480 ( .A(KEYINPUT82), .B(KEYINPUT81), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n422) );
  XNOR2_X1 U482 ( .A(G211GAT), .B(G78GAT), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U485 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n425), .B(KEYINPUT85), .ZN(n427) );
  XOR2_X1 U489 ( .A(n431), .B(n430), .Z(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n472) );
  NAND2_X1 U491 ( .A1(n573), .A2(n472), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n434), .B(KEYINPUT55), .ZN(n450) );
  INV_X1 U493 ( .A(n435), .ZN(n443) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XOR2_X1 U495 ( .A(G71GAT), .B(G176GAT), .Z(n437) );
  XNOR2_X1 U496 ( .A(G190GAT), .B(G183GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U498 ( .A(G43GAT), .B(G99GAT), .Z(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U502 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n445) );
  XNOR2_X1 U503 ( .A(G15GAT), .B(KEYINPUT80), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n535) );
  NAND2_X1 U507 ( .A1(n450), .A2(n535), .ZN(n562) );
  NOR2_X1 U508 ( .A1(n546), .A2(n562), .ZN(n454) );
  XNOR2_X1 U509 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n452) );
  INV_X1 U510 ( .A(G190GAT), .ZN(n451) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n455) );
  XNOR2_X1 U512 ( .A(n522), .B(n455), .ZN(n470) );
  INV_X1 U513 ( .A(n470), .ZN(n460) );
  NOR2_X1 U514 ( .A1(n535), .A2(n472), .ZN(n459) );
  XNOR2_X1 U515 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n457) );
  NAND2_X1 U516 ( .A1(n460), .A2(n574), .ZN(n461) );
  XNOR2_X1 U517 ( .A(KEYINPUT98), .B(n461), .ZN(n466) );
  INV_X1 U518 ( .A(n535), .ZN(n525) );
  OR2_X1 U519 ( .A1(n525), .A2(n522), .ZN(n462) );
  XOR2_X1 U520 ( .A(KEYINPUT99), .B(n462), .Z(n463) );
  NAND2_X1 U521 ( .A1(n463), .A2(n472), .ZN(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n467), .B(KEYINPUT100), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n468), .A2(n520), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n469), .B(KEYINPUT101), .ZN(n476) );
  NOR2_X1 U527 ( .A1(n520), .A2(n470), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT94), .B(n471), .Z(n533) );
  XOR2_X1 U529 ( .A(KEYINPUT28), .B(n472), .Z(n494) );
  NOR2_X1 U530 ( .A1(n533), .A2(n494), .ZN(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT95), .B(n473), .ZN(n474) );
  NOR2_X1 U532 ( .A1(n535), .A2(n474), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n485) );
  NOR2_X1 U534 ( .A1(n588), .A2(n485), .ZN(n477) );
  NAND2_X1 U535 ( .A1(n585), .A2(n477), .ZN(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT37), .B(n478), .ZN(n519) );
  NOR2_X1 U537 ( .A1(n575), .A2(n479), .ZN(n488) );
  NAND2_X1 U538 ( .A1(n519), .A2(n488), .ZN(n480) );
  NOR2_X1 U539 ( .A1(n522), .A2(n504), .ZN(n482) );
  XNOR2_X1 U540 ( .A(KEYINPUT16), .B(KEYINPUT77), .ZN(n484) );
  NOR2_X1 U541 ( .A1(n558), .A2(n585), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n486) );
  NOR2_X1 U543 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U544 ( .A(n487), .B(KEYINPUT102), .ZN(n506) );
  NAND2_X1 U545 ( .A1(n488), .A2(n506), .ZN(n495) );
  NOR2_X1 U546 ( .A1(n520), .A2(n495), .ZN(n489) );
  XOR2_X1 U547 ( .A(KEYINPUT34), .B(n489), .Z(n490) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n490), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n522), .A2(n495), .ZN(n491) );
  XOR2_X1 U550 ( .A(G8GAT), .B(n491), .Z(G1325GAT) );
  NOR2_X1 U551 ( .A1(n525), .A2(n495), .ZN(n493) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  INV_X1 U554 ( .A(n494), .ZN(n537) );
  NOR2_X1 U555 ( .A1(n537), .A2(n495), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1327GAT) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  NOR2_X1 U559 ( .A1(n520), .A2(n504), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n501) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n503) );
  NOR2_X1 U564 ( .A1(n525), .A2(n504), .ZN(n502) );
  XOR2_X1 U565 ( .A(n503), .B(n502), .Z(G1330GAT) );
  NOR2_X1 U566 ( .A1(n537), .A2(n504), .ZN(n505) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n505), .Z(G1331GAT) );
  XOR2_X1 U568 ( .A(n552), .B(KEYINPUT107), .Z(n565) );
  NOR2_X1 U569 ( .A1(n565), .A2(n550), .ZN(n518) );
  NAND2_X1 U570 ( .A1(n518), .A2(n506), .ZN(n515) );
  NOR2_X1 U571 ( .A1(n515), .A2(n520), .ZN(n510) );
  XOR2_X1 U572 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n508) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NOR2_X1 U576 ( .A1(n522), .A2(n515), .ZN(n511) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n525), .A2(n515), .ZN(n513) );
  XNOR2_X1 U579 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U582 ( .A1(n537), .A2(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n529) );
  NOR2_X1 U586 ( .A1(n520), .A2(n529), .ZN(n521) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n521), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n529), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U591 ( .A1(n525), .A2(n529), .ZN(n526) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(KEYINPUT113), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n531) );
  NOR2_X1 U596 ( .A1(n537), .A2(n529), .ZN(n530) );
  XOR2_X1 U597 ( .A(n531), .B(n530), .Z(G1339GAT) );
  NOR2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U599 ( .A(KEYINPUT117), .B(n534), .Z(n549) );
  AND2_X1 U600 ( .A1(n535), .A2(n549), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT118), .B(n536), .ZN(n538) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n575), .A2(n545), .ZN(n539) );
  XOR2_X1 U604 ( .A(G113GAT), .B(n539), .Z(G1340GAT) );
  NOR2_X1 U605 ( .A1(n565), .A2(n545), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NOR2_X1 U608 ( .A1(n571), .A2(n545), .ZN(n543) );
  XNOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  NOR2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n574), .A2(n549), .ZN(n556) );
  INV_X1 U616 ( .A(n556), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n559), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n556), .ZN(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n585), .A2(n556), .ZN(n557) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT120), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  NOR2_X1 U628 ( .A1(n575), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1348GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n562), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n567) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(KEYINPUT122), .B(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n562), .ZN(n572) );
  XOR2_X1 U638 ( .A(G183GAT), .B(n572), .Z(G1350GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n587) );
  NOR2_X1 U640 ( .A1(n575), .A2(n587), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT125), .B(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n587), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n587), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

