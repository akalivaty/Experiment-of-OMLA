//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0003(.A(G1), .ZN(new_n204));
  INV_X1    g0004(.A(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(G20), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n207), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n210), .B(new_n215), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT66), .Z(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n230), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n240), .B(new_n244), .Z(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n213), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NOR3_X1   g0049(.A1(KEYINPUT70), .A2(G20), .A3(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n205), .A2(G33), .ZN(new_n255));
  NOR3_X1   g0055(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n254), .A2(new_n255), .B1(new_n205), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n247), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G13), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n259), .A2(new_n205), .A3(G1), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n247), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n205), .A2(G1), .ZN(new_n262));
  INV_X1    g0062(.A(G50), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n261), .A2(new_n264), .B1(new_n263), .B2(new_n260), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G223), .A3(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G222), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n268), .B1(new_n216), .B2(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n213), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n204), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n204), .A2(G274), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT69), .A2(G45), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT69), .A2(G45), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(G226), .A2(new_n280), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n275), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n266), .B1(new_n289), .B2(G169), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n288), .A2(G179), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n266), .B(KEYINPUT9), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(G190), .ZN(new_n294));
  XOR2_X1   g0094(.A(KEYINPUT72), .B(G200), .Z(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n292), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n251), .A2(new_n263), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n255), .A2(new_n303), .B1(new_n205), .B2(G68), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n247), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT75), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT75), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(new_n247), .C1(new_n302), .C2(new_n304), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT11), .ZN(new_n310));
  INV_X1    g0110(.A(new_n260), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n311), .A2(KEYINPUT12), .A3(G68), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT12), .ZN(new_n313));
  INV_X1    g0113(.A(G68), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n260), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n261), .ZN(new_n316));
  OAI21_X1  g0116(.A(G68), .B1(new_n205), .B2(G1), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n312), .A2(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n309), .B2(KEYINPUT11), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n232), .A2(G1698), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n267), .B(new_n323), .C1(G226), .C2(G1698), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n277), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n282), .A2(new_n286), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n280), .A2(G238), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n327), .A2(new_n328), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n329), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT13), .B1(new_n332), .B2(new_n326), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n322), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n331), .A2(new_n333), .A3(G179), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n334), .B2(new_n335), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n320), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n331), .A2(new_n333), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G200), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n331), .A2(new_n333), .A3(G190), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n310), .A2(new_n341), .A3(new_n319), .A4(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n301), .B1(new_n344), .B2(KEYINPUT77), .ZN(new_n345));
  OAI21_X1  g0145(.A(G77), .B1(new_n205), .B2(G1), .ZN(new_n346));
  INV_X1    g0146(.A(new_n216), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n316), .A2(new_n346), .B1(new_n347), .B2(new_n311), .ZN(new_n348));
  OR3_X1    g0148(.A1(KEYINPUT70), .A2(G20), .A3(G33), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n248), .ZN(new_n350));
  INV_X1    g0150(.A(new_n254), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n350), .A2(new_n351), .B1(new_n347), .B2(G20), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT15), .B(G87), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT71), .B1(new_n353), .B2(new_n255), .ZN(new_n354));
  OR3_X1    g0154(.A1(new_n353), .A2(KEYINPUT71), .A3(new_n255), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n348), .B1(new_n356), .B2(new_n247), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n329), .B1(new_n217), .B2(new_n279), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n267), .A2(G238), .A3(G1698), .ZN(new_n359));
  INV_X1    g0159(.A(G107), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n359), .B1(new_n360), .B2(new_n267), .C1(new_n270), .C2(new_n232), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n358), .B1(new_n361), .B2(new_n274), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n357), .B1(new_n362), .B2(new_n295), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(KEYINPUT73), .B1(G190), .B2(new_n362), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT73), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n357), .B(new_n365), .C1(new_n362), .C2(new_n295), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n362), .A2(G169), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n357), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT74), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n339), .A2(KEYINPUT77), .A3(new_n343), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n367), .A2(new_n376), .A3(new_n372), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  OR2_X1    g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NAND2_X1  g0180(.A1(KEYINPUT3), .A2(G33), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n205), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n380), .A2(KEYINPUT7), .A3(new_n205), .A4(new_n381), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n314), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(G58), .B(G68), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G20), .ZN(new_n388));
  INV_X1    g0188(.A(G159), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n251), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n379), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(KEYINPUT3), .A2(G33), .ZN(new_n392));
  NOR2_X1   g0192(.A1(KEYINPUT3), .A2(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT7), .B1(new_n394), .B2(new_n205), .ZN(new_n395));
  INV_X1    g0195(.A(new_n385), .ZN(new_n396));
  OAI21_X1  g0196(.A(G68), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n350), .A2(G159), .B1(new_n387), .B2(G20), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(KEYINPUT16), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n391), .A2(new_n399), .A3(new_n247), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n254), .A2(new_n262), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n316), .B1(KEYINPUT78), .B2(new_n401), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n401), .A2(KEYINPUT78), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n402), .A2(new_n403), .B1(new_n260), .B2(new_n254), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT79), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT79), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n400), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(G232), .A2(new_n280), .B1(new_n282), .B2(new_n286), .ZN(new_n409));
  OR2_X1    g0209(.A1(G223), .A2(G1698), .ZN(new_n410));
  INV_X1    g0210(.A(G226), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G1698), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n410), .B(new_n412), .C1(new_n392), .C2(new_n393), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G87), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n277), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G169), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n369), .B2(new_n417), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n406), .A2(new_n408), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT18), .ZN(new_n421));
  INV_X1    g0221(.A(G200), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n409), .B2(new_n416), .ZN(new_n423));
  INV_X1    g0223(.A(new_n286), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n277), .A2(new_n281), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n424), .A2(new_n425), .B1(new_n232), .B2(new_n279), .ZN(new_n426));
  INV_X1    g0226(.A(G190), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n426), .A2(new_n415), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(new_n400), .A3(new_n404), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT17), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n406), .A2(new_n432), .A3(new_n408), .A4(new_n419), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n421), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n345), .A2(new_n378), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n267), .A2(G264), .A3(G1698), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n267), .A2(G257), .A3(new_n269), .ZN(new_n438));
  INV_X1    g0238(.A(G303), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n437), .B(new_n438), .C1(new_n439), .C2(new_n267), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n274), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT5), .B(G41), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n204), .A2(G45), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(G270), .A3(new_n277), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n204), .A2(G45), .A3(G274), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n214), .B2(new_n276), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n447), .B1(new_n449), .B2(new_n442), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n204), .A2(G45), .A3(G274), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n442), .A2(new_n451), .A3(new_n447), .A4(new_n277), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(KEYINPUT89), .B(new_n446), .C1(new_n450), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n442), .A2(new_n277), .A3(new_n451), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n452), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT89), .B1(new_n458), .B2(new_n446), .ZN(new_n459));
  OAI211_X1 g0259(.A(G190), .B(new_n441), .C1(new_n455), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(G20), .B1(G33), .B2(G283), .ZN(new_n461));
  INV_X1    g0261(.A(G33), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G97), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT91), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT91), .ZN(new_n467));
  INV_X1    g0267(.A(G116), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n246), .A2(new_n213), .B1(G20), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT20), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n466), .A2(KEYINPUT20), .A3(new_n467), .A4(new_n469), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT90), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n311), .B2(G116), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n260), .A2(KEYINPUT90), .A3(new_n468), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n462), .A2(G1), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n260), .A2(new_n247), .A3(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n476), .A2(new_n477), .B1(new_n479), .B2(G116), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n441), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n446), .B1(new_n450), .B2(new_n453), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT89), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n483), .B1(new_n486), .B2(new_n454), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n460), .B(new_n482), .C1(new_n487), .C2(new_n422), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT21), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n481), .A2(G169), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(G179), .A3(new_n481), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n441), .B1(new_n455), .B2(new_n459), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(KEYINPUT21), .A3(G169), .A4(new_n481), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n488), .A2(new_n491), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n205), .A2(G107), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT23), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT23), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n205), .B2(G107), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n462), .A2(new_n468), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n497), .A2(new_n499), .B1(new_n205), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n205), .B(G87), .C1(new_n392), .C2(new_n393), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n502), .A2(KEYINPUT22), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(KEYINPUT22), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT24), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(KEYINPUT24), .B(new_n501), .C1(new_n503), .C2(new_n504), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n247), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n479), .A2(G107), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n259), .A2(G1), .ZN(new_n511));
  OR2_X1    g0311(.A1(KEYINPUT92), .A2(KEYINPUT25), .ZN(new_n512));
  NAND2_X1  g0312(.A1(KEYINPUT92), .A2(KEYINPUT25), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n511), .A2(new_n496), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n511), .A2(new_n496), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n510), .B(new_n514), .C1(new_n513), .C2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G257), .B(G1698), .C1(new_n392), .C2(new_n393), .ZN(new_n519));
  OAI211_X1 g0319(.A(G250), .B(new_n269), .C1(new_n392), .C2(new_n393), .ZN(new_n520));
  INV_X1    g0320(.A(G294), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n519), .B(new_n520), .C1(new_n462), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n274), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n274), .B1(new_n444), .B2(new_n442), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G264), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n458), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT93), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(G169), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n522), .A2(new_n274), .B1(new_n524), .B2(G264), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(G179), .A3(new_n458), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n527), .B1(new_n526), .B2(G169), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n518), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n526), .A2(G190), .ZN(new_n534));
  AOI21_X1  g0334(.A(G200), .B1(new_n529), .B2(new_n458), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n509), .B(new_n517), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n538));
  NOR2_X1   g0338(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n539));
  INV_X1    g0339(.A(G97), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(G107), .ZN(new_n541));
  XNOR2_X1  g0341(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n542));
  XNOR2_X1  g0342(.A(G97), .B(G107), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(G20), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n350), .A2(G77), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n360), .B1(new_n384), .B2(new_n385), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n247), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT83), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n311), .A2(G97), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n479), .B2(G97), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n548), .B2(new_n551), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n457), .A2(new_n452), .B1(new_n524), .B2(G257), .ZN(new_n555));
  OAI211_X1 g0355(.A(G244), .B(new_n269), .C1(new_n392), .C2(new_n393), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT4), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G283), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n462), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G250), .A2(G1698), .ZN(new_n561));
  NAND2_X1  g0361(.A1(KEYINPUT4), .A2(G244), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(G1698), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n267), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n274), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT84), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n555), .A2(new_n566), .A3(new_n567), .A4(new_n369), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n555), .A2(new_n369), .A3(new_n566), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT84), .ZN(new_n570));
  AOI21_X1  g0370(.A(G169), .B1(new_n555), .B2(new_n566), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n548), .A2(new_n551), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n445), .A2(G257), .A3(new_n277), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n450), .B2(new_n453), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n277), .B1(new_n558), .B2(new_n564), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n573), .B1(G190), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n555), .A2(new_n566), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT82), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n555), .A2(KEYINPUT82), .A3(new_n566), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(G200), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n554), .A2(new_n572), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n205), .B1(new_n325), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G87), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n540), .A3(new_n360), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n205), .B(G68), .C1(new_n392), .C2(new_n393), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n585), .B1(new_n255), .B2(new_n540), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n247), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n353), .A2(new_n260), .ZN(new_n594));
  INV_X1    g0394(.A(new_n353), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n479), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n277), .A2(G250), .A3(new_n443), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G238), .A2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n217), .B2(G1698), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n500), .B1(new_n600), .B2(new_n267), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n598), .B1(new_n601), .B2(new_n277), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT85), .B1(new_n274), .B2(new_n448), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT85), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n451), .A2(new_n277), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(G169), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n598), .ZN(new_n608));
  INV_X1    g0408(.A(G238), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n269), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n217), .A2(G1698), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n610), .B(new_n611), .C1(new_n392), .C2(new_n393), .ZN(new_n612));
  INV_X1    g0412(.A(new_n500), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n608), .B1(new_n614), .B2(new_n274), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n603), .A2(new_n605), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(G179), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n607), .A2(KEYINPUT86), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT86), .B1(new_n607), .B2(new_n617), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n597), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n614), .A2(new_n274), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(new_n616), .A3(G190), .A4(new_n598), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT87), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT87), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n615), .A2(new_n624), .A3(G190), .A4(new_n616), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT88), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n623), .A2(new_n628), .A3(new_n625), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n479), .A2(G87), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n593), .A2(new_n594), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n615), .A2(new_n616), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n296), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n627), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n584), .A2(new_n620), .A3(new_n634), .ZN(new_n635));
  NOR4_X1   g0435(.A1(new_n436), .A2(new_n495), .A3(new_n537), .A4(new_n635), .ZN(G372));
  XNOR2_X1  g0436(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n405), .A2(new_n419), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n405), .A2(new_n419), .ZN(new_n639));
  INV_X1    g0439(.A(new_n637), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n339), .A2(new_n372), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n431), .A2(new_n343), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n638), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n299), .A2(new_n300), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n292), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n607), .A2(new_n617), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n597), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n626), .A2(new_n633), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n572), .A2(new_n573), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n634), .A2(new_n572), .A3(new_n620), .A4(new_n554), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n651), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n533), .A2(new_n491), .A3(new_n492), .A4(new_n494), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n626), .A2(new_n633), .B1(new_n647), .B2(new_n597), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n536), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n584), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n654), .A2(new_n648), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n646), .B1(new_n436), .B2(new_n660), .ZN(G369));
  NAND3_X1  g0461(.A1(new_n491), .A2(new_n494), .A3(new_n492), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n511), .A2(new_n205), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n482), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n495), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n669), .B1(new_n509), .B2(new_n517), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n537), .A2(new_n675), .B1(new_n533), .B2(new_n669), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n662), .A2(new_n669), .ZN(new_n678));
  INV_X1    g0478(.A(new_n537), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n533), .A2(new_n668), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n677), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n208), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n588), .A2(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n211), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  NOR4_X1   g0490(.A1(new_n635), .A2(new_n495), .A3(new_n537), .A4(new_n668), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  OAI211_X1 g0492(.A(G179), .B(new_n441), .C1(new_n455), .C2(new_n459), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n602), .A2(new_n606), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n577), .A2(new_n529), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n692), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n523), .A2(new_n525), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n579), .A2(new_n697), .A3(new_n632), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n487), .A3(KEYINPUT30), .A4(G179), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n694), .A2(G179), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n493), .A2(new_n526), .A3(new_n579), .A4(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n668), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n691), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G330), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n653), .A2(KEYINPUT26), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n648), .A3(new_n658), .A4(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n714), .B2(new_n669), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n659), .A2(new_n711), .A3(new_n669), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n710), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n690), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n259), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n204), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n685), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n674), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n672), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n208), .A2(new_n267), .ZN(new_n725));
  INV_X1    g0525(.A(G355), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n725), .A2(new_n726), .B1(G116), .B2(new_n208), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n208), .A2(new_n394), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT95), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n283), .A2(new_n285), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n730), .B1(new_n212), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n244), .A2(G45), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n727), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT96), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n213), .B1(G20), .B2(new_n321), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n722), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n427), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n369), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n205), .A2(G179), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G190), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n389), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT32), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n746), .A2(new_n540), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n394), .B(new_n752), .C1(new_n751), .C2(new_n750), .ZN(new_n753));
  NAND2_X1  g0553(.A1(G20), .A2(G179), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT97), .Z(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(new_n427), .A3(G200), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n753), .B1(new_n263), .B2(new_n756), .C1(new_n314), .C2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n296), .A2(G190), .A3(new_n747), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n755), .A2(new_n743), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G87), .A2(new_n760), .B1(new_n762), .B2(G58), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n755), .A2(new_n748), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n296), .A2(new_n427), .A3(new_n747), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT98), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT98), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n763), .B1(new_n216), .B2(new_n764), .C1(new_n769), .C2(new_n360), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n559), .ZN(new_n771));
  INV_X1    g0571(.A(new_n756), .ZN(new_n772));
  INV_X1    g0572(.A(new_n757), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT33), .B(G317), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G326), .A2(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n749), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n267), .B1(new_n776), .B2(G329), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n521), .B2(new_n746), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n762), .B2(G322), .ZN(new_n779));
  INV_X1    g0579(.A(new_n764), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G303), .A2(new_n760), .B1(new_n780), .B2(G311), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n775), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n758), .A2(new_n770), .B1(new_n771), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n784));
  INV_X1    g0584(.A(new_n739), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n783), .B2(KEYINPUT99), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n742), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n738), .B(KEYINPUT100), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n672), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n724), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  NOR2_X1   g0591(.A1(new_n357), .A2(new_n669), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT102), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n367), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n372), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n372), .A2(new_n668), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n660), .B2(new_n668), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n367), .A2(new_n793), .A3(new_n372), .A4(new_n669), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n659), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n710), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n722), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n710), .A2(new_n802), .A3(new_n799), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n394), .B1(new_n776), .B2(G132), .ZN(new_n807));
  INV_X1    g0607(.A(G58), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n746), .B2(new_n808), .C1(new_n759), .C2(new_n263), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n810), .A2(new_n756), .B1(new_n757), .B2(new_n252), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT101), .Z(new_n812));
  AOI22_X1  g0612(.A1(G143), .A2(new_n762), .B1(new_n780), .B2(G159), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT34), .Z(new_n815));
  INV_X1    g0615(.A(new_n769), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n809), .B(new_n815), .C1(G68), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(G87), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G283), .A2(new_n773), .B1(new_n772), .B2(G303), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n394), .B1(new_n749), .B2(new_n820), .C1(new_n746), .C2(new_n540), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n762), .B2(G294), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G107), .A2(new_n760), .B1(new_n780), .B2(G116), .ZN(new_n823));
  AND4_X1   g0623(.A1(new_n818), .A2(new_n819), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n739), .B1(new_n817), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n722), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n739), .A2(new_n736), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n303), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n796), .B1(new_n794), .B2(new_n372), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n825), .B(new_n828), .C1(new_n737), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n806), .A2(new_n830), .ZN(G384));
  NOR2_X1   g0631(.A1(new_n719), .A2(new_n204), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT40), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT107), .B1(new_n691), .B2(new_n707), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n320), .A2(new_n668), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n339), .A2(new_n343), .A3(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n320), .B(new_n668), .C1(new_n336), .C2(new_n338), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n798), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n554), .A2(new_n572), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n578), .A2(new_n583), .ZN(new_n841));
  AND4_X1   g0641(.A1(new_n840), .A2(new_n634), .A3(new_n841), .A4(new_n620), .ZN(new_n842));
  INV_X1    g0642(.A(new_n495), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n842), .A2(new_n843), .A3(new_n679), .A4(new_n669), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT107), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n844), .A2(new_n845), .A3(new_n705), .A4(new_n706), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n834), .A2(new_n839), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n666), .B1(new_n400), .B2(new_n404), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n434), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n666), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n406), .A2(new_n408), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n430), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n420), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n639), .A2(new_n430), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n855), .B2(new_n848), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n849), .A2(KEYINPUT38), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT38), .B1(new_n849), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n833), .B1(new_n847), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n862));
  INV_X1    g0662(.A(new_n854), .ZN(new_n863));
  INV_X1    g0663(.A(new_n855), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n852), .B1(new_n864), .B2(new_n851), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n641), .A2(new_n638), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n851), .B1(new_n868), .B2(new_n431), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n862), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n849), .A2(KEYINPUT38), .A3(new_n857), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n833), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n872), .A2(new_n839), .A3(new_n834), .A4(new_n846), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n861), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n435), .A2(new_n834), .A3(new_n846), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n709), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n874), .B2(new_n875), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n870), .A2(new_n871), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n339), .A2(new_n668), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n849), .A2(new_n857), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n871), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n871), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n836), .A2(new_n837), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n796), .B(KEYINPUT104), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n890), .B1(new_n802), .B2(new_n892), .ZN(new_n893));
  AOI211_X1 g0693(.A(KEYINPUT105), .B(new_n891), .C1(new_n659), .C2(new_n801), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n888), .B(new_n889), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n867), .A2(new_n666), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n887), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n435), .B1(new_n715), .B2(new_n716), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n646), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n897), .B(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n832), .B1(new_n877), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n900), .B2(new_n877), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n213), .A2(new_n205), .A3(new_n468), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT35), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n905), .B2(new_n904), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT36), .Z(new_n908));
  OAI21_X1  g0708(.A(new_n212), .B1(new_n808), .B2(new_n314), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n909), .A2(new_n216), .B1(G50), .B2(new_n314), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(G1), .A3(new_n259), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT103), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n902), .A2(new_n913), .ZN(G367));
  NAND2_X1  g0714(.A1(new_n668), .A2(new_n631), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n656), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n648), .A2(new_n915), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT43), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n572), .A2(new_n573), .A3(new_n668), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT108), .Z(new_n924));
  INV_X1    g0724(.A(new_n573), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n584), .B1(new_n925), .B2(new_n669), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n680), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT42), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n929), .B(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n928), .A2(new_n533), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n668), .B1(new_n932), .B2(new_n840), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n921), .B(new_n922), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n933), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n929), .B(KEYINPUT42), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n935), .A2(new_n936), .A3(new_n920), .A4(new_n919), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n677), .A2(new_n928), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n934), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n677), .B2(new_n928), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n685), .B(KEYINPUT41), .Z(new_n942));
  NOR2_X1   g0742(.A1(new_n682), .A2(new_n927), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT44), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n682), .A2(new_n927), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT45), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n677), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n717), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n680), .B1(new_n676), .B2(new_n678), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n673), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n944), .A2(new_n677), .A3(new_n947), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n942), .B1(new_n956), .B2(new_n717), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n939), .B(new_n941), .C1(new_n957), .C2(new_n721), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n816), .A2(new_n347), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n267), .B1(new_n749), .B2(new_n810), .C1(new_n746), .C2(new_n314), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G58), .B2(new_n760), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G50), .A2(new_n780), .B1(new_n762), .B2(G150), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G143), .A2(new_n772), .B1(new_n773), .B2(G159), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n959), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n816), .A2(G97), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n760), .A2(KEYINPUT46), .A3(G116), .ZN(new_n966));
  INV_X1    g0766(.A(G317), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n394), .B1(new_n749), .B2(new_n967), .C1(new_n746), .C2(new_n360), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n780), .B2(G283), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT46), .B1(new_n760), .B2(G116), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G294), .B2(new_n773), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n965), .A2(new_n966), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n756), .A2(new_n820), .B1(new_n761), .B2(new_n439), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT109), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n964), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n739), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n918), .A2(new_n788), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n729), .A2(new_n229), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n979), .B(new_n740), .C1(new_n208), .C2(new_n353), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n977), .A2(new_n722), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n958), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT110), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n958), .A2(KEYINPUT110), .A3(new_n981), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(G387));
  NOR2_X1   g0787(.A1(new_n953), .A2(new_n720), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT111), .Z(new_n989));
  NOR2_X1   g0789(.A1(new_n676), .A2(new_n788), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n729), .B1(new_n235), .B2(new_n732), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n687), .B2(new_n725), .ZN(new_n992));
  OR3_X1    g0792(.A1(new_n254), .A2(KEYINPUT50), .A3(G50), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT50), .B1(new_n254), .B2(G50), .ZN(new_n994));
  AOI21_X1  g0794(.A(G45), .B1(G68), .B2(G77), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n993), .A2(new_n687), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n992), .A2(new_n996), .B1(new_n360), .B2(new_n684), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n722), .B1(new_n997), .B2(new_n741), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n216), .A2(new_n759), .B1(new_n761), .B2(new_n263), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n394), .B1(new_n776), .B2(G150), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n746), .B2(new_n353), .C1(new_n764), .C2(new_n314), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n999), .B(new_n1001), .C1(new_n351), .C2(new_n773), .ZN(new_n1002));
  OR3_X1    g0802(.A1(new_n756), .A2(KEYINPUT112), .A3(new_n389), .ZN(new_n1003));
  OAI21_X1  g0803(.A(KEYINPUT112), .B1(new_n756), .B2(new_n389), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n965), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n267), .B1(new_n776), .B2(G326), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n759), .A2(new_n521), .B1(new_n746), .B2(new_n559), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G303), .A2(new_n780), .B1(new_n762), .B2(G317), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n772), .A2(G322), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(new_n820), .C2(new_n757), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1006), .B1(new_n468), .B2(new_n769), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1005), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n990), .B(new_n998), .C1(new_n1017), .C2(new_n739), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n989), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n954), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n951), .A2(new_n953), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n685), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(new_n1022), .ZN(G393));
  AND2_X1   g0823(.A1(new_n956), .A2(new_n685), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n950), .A2(new_n955), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n1020), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n950), .A2(new_n721), .A3(new_n955), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n928), .A2(new_n738), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n394), .B1(new_n776), .B2(G143), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n745), .A2(G77), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n314), .B2(new_n759), .C1(new_n254), .C2(new_n764), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G50), .B2(new_n773), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n756), .A2(new_n252), .B1(new_n761), .B2(new_n389), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT51), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n818), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n267), .B1(new_n776), .B2(G322), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n746), .B2(new_n468), .C1(new_n759), .C2(new_n559), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G294), .B2(new_n780), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n439), .B2(new_n757), .C1(new_n360), .C2(new_n769), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n756), .A2(new_n967), .B1(new_n761), .B2(new_n820), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT52), .Z(new_n1043));
  OAI21_X1  g0843(.A(new_n1037), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT113), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n739), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n740), .B1(new_n540), .B2(new_n208), .C1(new_n730), .C2(new_n239), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1029), .A2(new_n1046), .A3(new_n722), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT114), .B1(new_n1028), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1028), .A2(KEYINPUT114), .A3(new_n1048), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1027), .B1(new_n1049), .B2(new_n1051), .ZN(G390));
  NAND4_X1  g0852(.A1(new_n834), .A2(new_n839), .A3(G330), .A4(new_n846), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n889), .B1(new_n893), .B2(new_n894), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1055), .A2(new_n881), .B1(new_n880), .B2(new_n886), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n658), .A2(new_n648), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n713), .B1(new_n653), .B2(KEYINPUT26), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n669), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n797), .B1(new_n1059), .B2(new_n798), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n889), .B(KEYINPUT115), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(new_n881), .A3(new_n878), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1054), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(G330), .B(new_n829), .C1(new_n691), .C2(new_n707), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1066), .A2(new_n838), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n648), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n657), .A2(new_n584), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n655), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n800), .B1(new_n1071), .B2(new_n654), .ZN(new_n1072));
  OAI21_X1  g0872(.A(KEYINPUT105), .B1(new_n1072), .B2(new_n891), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n802), .A2(new_n890), .A3(new_n892), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n882), .B1(new_n1075), .B2(new_n889), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n880), .A2(new_n886), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1063), .B(new_n1068), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1065), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n435), .A2(G330), .A3(new_n834), .A4(new_n846), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n898), .A3(new_n646), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1067), .A2(new_n1060), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n834), .A2(G330), .A3(new_n829), .A4(new_n846), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1061), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1066), .A2(new_n838), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1053), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1075), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1082), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1080), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1065), .A2(new_n1079), .A3(new_n1091), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n685), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1065), .A2(new_n1079), .A3(new_n721), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n827), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n722), .B1(new_n351), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n816), .A2(G68), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1031), .B(new_n394), .C1(new_n521), .C2(new_n749), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G87), .B2(new_n760), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G97), .A2(new_n780), .B1(new_n762), .B2(G116), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G107), .A2(new_n773), .B1(new_n772), .B2(G283), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n267), .B1(new_n769), .B2(new_n263), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1106));
  INV_X1    g0906(.A(G128), .ZN(new_n1107));
  INV_X1    g0907(.A(G132), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n756), .A2(new_n1107), .B1(new_n761), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT118), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1106), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n773), .A2(G137), .B1(new_n780), .B2(new_n1114), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n1115), .A2(KEYINPUT116), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n759), .A2(new_n252), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(KEYINPUT116), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n745), .A2(G159), .B1(new_n776), .B2(G125), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1104), .B1(new_n1112), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1098), .B1(new_n1122), .B2(new_n739), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1078), .B2(new_n737), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1096), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1095), .A2(new_n1125), .ZN(G378));
  INV_X1    g0926(.A(new_n1082), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1094), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n266), .A2(new_n850), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n301), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n301), .A2(new_n1129), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OR3_X1    g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1134), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AND4_X1   g0937(.A1(G330), .A2(new_n861), .A3(new_n873), .A4(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n834), .A2(new_n839), .A3(new_n846), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n709), .B1(new_n1139), .B2(new_n872), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1137), .B1(new_n1140), .B2(new_n861), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n897), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n861), .A2(new_n873), .A3(G330), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1137), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n887), .A2(new_n895), .A3(new_n896), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1140), .A2(new_n861), .A3(new_n1137), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1128), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT57), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1151), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n686), .B1(new_n1153), .B2(new_n1128), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1138), .A2(new_n1141), .A3(new_n897), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1146), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n721), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n722), .B1(G50), .B2(new_n1097), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n267), .A2(G41), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G50), .B(new_n1160), .C1(new_n462), .C2(new_n284), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n816), .A2(G58), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1160), .B1(new_n559), .B2(new_n749), .C1(new_n746), .C2(new_n314), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n360), .A2(new_n761), .B1(new_n764), .B2(new_n353), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n347), .C2(new_n760), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G97), .A2(new_n773), .B1(new_n772), .B2(G116), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1162), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT58), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1161), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G125), .A2(new_n772), .B1(new_n773), .B2(G132), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n760), .A2(new_n1114), .B1(G150), .B2(new_n745), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G128), .A2(new_n762), .B1(new_n780), .B2(G137), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G33), .B(G41), .C1(new_n776), .C2(G124), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n389), .C2(new_n769), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1169), .B1(new_n1168), .B2(new_n1167), .C1(new_n1174), .C2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1159), .B1(new_n1178), .B2(new_n739), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n1137), .B2(new_n737), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT119), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1158), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1155), .A2(new_n1183), .ZN(G375));
  AOI22_X1  g0984(.A1(new_n1086), .A2(new_n1083), .B1(new_n1089), .B2(new_n1075), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(new_n720), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT121), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n468), .A2(new_n757), .B1(new_n756), .B2(new_n521), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G107), .A2(new_n780), .B1(new_n762), .B2(G283), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n394), .B1(new_n749), .B2(new_n439), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n595), .B2(new_n745), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1189), .B(new_n1191), .C1(new_n540), .C2(new_n759), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1188), .B(new_n1192), .C1(new_n816), .C2(G77), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n267), .B1(new_n749), .B2(new_n1107), .C1(new_n746), .C2(new_n263), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G150), .B2(new_n780), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1162), .B(new_n1195), .C1(new_n389), .C2(new_n759), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(KEYINPUT120), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n762), .A2(G137), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n1108), .B2(new_n756), .C1(new_n757), .C2(new_n1113), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1196), .B2(KEYINPUT120), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1193), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n722), .B1(G68), .B2(new_n1097), .C1(new_n1201), .C2(new_n785), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1085), .B2(new_n736), .ZN(new_n1203));
  OR3_X1    g1003(.A1(new_n1186), .A2(new_n1187), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1187), .B1(new_n1186), .B2(new_n1203), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1185), .A2(new_n1082), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1091), .A2(new_n942), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1204), .A2(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(G381));
  INV_X1    g1009(.A(G378), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1049), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1211), .A2(new_n1050), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1212));
  INV_X1    g1012(.A(G384), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n986), .A2(new_n1210), .A3(new_n1208), .A4(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(G375), .ZN(G407));
  NAND2_X1  g1017(.A1(new_n667), .A2(G213), .ZN(new_n1218));
  OR3_X1    g1018(.A1(G375), .A2(G378), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(G213), .A3(new_n1219), .ZN(G409));
  AOI221_X4 g1020(.A(new_n1182), .B1(new_n1095), .B2(new_n1125), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT122), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n942), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1222), .B1(new_n1223), .B2(new_n1128), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1158), .A2(new_n1180), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1128), .A3(new_n1222), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G378), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1218), .B1(new_n1221), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1206), .B1(new_n1091), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT123), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1087), .A2(new_n1090), .A3(new_n1082), .A4(KEYINPUT60), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT124), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1185), .A2(new_n1235), .A3(KEYINPUT60), .A4(new_n1082), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n686), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT123), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1206), .B(new_n1238), .C1(new_n1091), .C2(new_n1230), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1232), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1240), .A2(new_n1241), .A3(G384), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G384), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1243));
  INV_X1    g1043(.A(G2897), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1242), .A2(new_n1243), .B1(new_n1244), .B2(new_n1218), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1213), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1240), .A2(new_n1241), .A3(G384), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1218), .A2(new_n1244), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1245), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT61), .B1(new_n1229), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1155), .A2(G378), .A3(new_n1183), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1227), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1254), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1253), .B1(G378), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT62), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1218), .A4(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1218), .B(new_n1258), .C1(new_n1221), .C2(new_n1228), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1252), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G390), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1212), .A2(KEYINPUT126), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n984), .A2(new_n985), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(G393), .B(new_n790), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n982), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1268), .B2(G390), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n982), .A2(new_n1212), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(G390), .A2(new_n958), .A3(new_n981), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1266), .A2(new_n1269), .B1(new_n1272), .B2(new_n1267), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1262), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(KEYINPUT61), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1251), .A2(KEYINPUT125), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT125), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1245), .A2(new_n1250), .A3(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(new_n1229), .A3(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1256), .A2(KEYINPUT63), .A3(new_n1218), .A4(new_n1258), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1260), .A2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1275), .A2(new_n1279), .A3(new_n1280), .A4(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1274), .A2(new_n1283), .ZN(G405));
  INV_X1    g1084(.A(KEYINPUT127), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G378), .B1(new_n1155), .B2(new_n1183), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1253), .A3(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1258), .B1(new_n1221), .B2(new_n1286), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1272), .A2(new_n1267), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1285), .B1(new_n1291), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1273), .A2(new_n1289), .A3(new_n1290), .A4(KEYINPUT127), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(G402));
endmodule


