//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT82), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT4), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G127gat), .ZN(new_n212));
  INV_X1    g011(.A(G127gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G113gat), .B(G120gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n216), .B(new_n217), .C1(KEYINPUT1), .C2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G120gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G113gat), .ZN(new_n221));
  INV_X1    g020(.A(G113gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G120gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT71), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT71), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n221), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  XNOR2_X1  g028(.A(G127gat), .B(G134gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n219), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT2), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT81), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT81), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT2), .ZN(new_n238));
  NAND2_X1  g037(.A1(G141gat), .A2(G148gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n234), .A2(new_n236), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(G155gat), .A2(G162gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(G141gat), .A2(G148gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(new_n233), .ZN(new_n246));
  XNOR2_X1  g045(.A(G155gat), .B(G162gat), .ZN(new_n247));
  INV_X1    g046(.A(G155gat), .ZN(new_n248));
  INV_X1    g047(.A(G162gat), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT2), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n246), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n210), .B1(new_n232), .B2(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n246), .A2(new_n247), .A3(new_n250), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT81), .B(KEYINPUT2), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n247), .B1(new_n246), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT3), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n244), .A2(new_n258), .A3(new_n251), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n232), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n254), .A2(new_n256), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n225), .A2(new_n229), .A3(new_n230), .A4(new_n228), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n262), .A4(new_n219), .ZN(new_n263));
  AND4_X1   g062(.A1(new_n209), .A2(new_n253), .A3(new_n260), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n253), .A2(new_n260), .A3(new_n263), .ZN(new_n266));
  INV_X1    g065(.A(new_n209), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n261), .A2(new_n219), .A3(new_n262), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n232), .A2(new_n252), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n209), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n271));
  OAI22_X1  g070(.A1(new_n266), .A2(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n207), .B1(new_n265), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT84), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT6), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n268), .A2(new_n269), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n271), .B1(new_n276), .B2(new_n267), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n264), .A2(new_n277), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n266), .A2(new_n271), .A3(new_n267), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n206), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT84), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n272), .A3(new_n207), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n275), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n265), .A2(new_n272), .A3(KEYINPUT6), .A4(new_n207), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n286));
  XNOR2_X1  g085(.A(G211gat), .B(G218gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G211gat), .A2(G218gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT75), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G197gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G204gat), .ZN(new_n294));
  INV_X1    g093(.A(G204gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G197gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n288), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n298), .ZN(new_n300));
  XNOR2_X1  g099(.A(G197gat), .B(G204gat), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n300), .A2(new_n287), .A3(new_n301), .A4(new_n292), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304));
  OR2_X1    g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT64), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n308), .B2(new_n307), .ZN(new_n310));
  INV_X1    g109(.A(G169gat), .ZN(new_n311));
  INV_X1    g110(.A(G176gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(KEYINPUT65), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT65), .ZN(new_n316));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(KEYINPUT23), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n321), .B1(KEYINPUT23), .B2(new_n317), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n304), .B1(new_n310), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n305), .A2(new_n306), .ZN(new_n325));
  INV_X1    g124(.A(new_n307), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n304), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(new_n319), .A3(new_n322), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT26), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n330), .A3(new_n320), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n317), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT69), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT69), .B1(new_n331), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT27), .B(G183gat), .ZN(new_n336));
  INV_X1    g135(.A(G190gat), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n336), .A2(KEYINPUT28), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT27), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(new_n337), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT28), .B1(new_n343), .B2(KEYINPUT67), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n340), .A2(new_n342), .A3(new_n345), .A4(new_n337), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n338), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n335), .B1(new_n347), .B2(KEYINPUT68), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT68), .ZN(new_n349));
  AOI211_X1 g148(.A(new_n349), .B(new_n338), .C1(new_n346), .C2(new_n344), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n329), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n352), .B(KEYINPUT76), .Z(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n344), .A2(new_n346), .ZN(new_n355));
  INV_X1    g154(.A(new_n338), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n349), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n347), .A2(KEYINPUT68), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n335), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n360), .B2(new_n329), .ZN(new_n361));
  INV_X1    g160(.A(new_n352), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n303), .B(new_n354), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n299), .A2(new_n302), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n353), .B1(new_n351), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n352), .B1(new_n360), .B2(new_n329), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT77), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n363), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n286), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n374), .A2(new_n286), .A3(new_n375), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n285), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n351), .A2(new_n365), .ZN(new_n379));
  INV_X1    g178(.A(new_n353), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n351), .A2(new_n362), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n303), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n362), .B1(new_n351), .B2(new_n365), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n380), .B1(new_n360), .B2(new_n329), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n384), .A2(new_n385), .A3(new_n364), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n372), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n363), .A2(new_n368), .A3(KEYINPUT30), .A4(new_n373), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(KEYINPUT78), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n363), .A2(new_n368), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT30), .A4(new_n373), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT79), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT79), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n389), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n378), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT85), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT86), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n299), .A2(new_n302), .A3(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(KEYINPUT86), .B(new_n288), .C1(new_n297), .C2(new_n298), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n365), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n261), .B1(new_n403), .B2(new_n258), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n303), .B1(new_n365), .B2(new_n259), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n399), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT29), .B1(new_n261), .B2(new_n258), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(new_n303), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(KEYINPUT87), .ZN(new_n410));
  INV_X1    g209(.A(new_n398), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT29), .B1(new_n299), .B2(new_n302), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n252), .B1(new_n412), .B2(KEYINPUT3), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n409), .A2(new_n410), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G22gat), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n406), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n415), .B1(new_n406), .B2(new_n414), .ZN(new_n417));
  OAI21_X1  g216(.A(G78gat), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n406), .A2(new_n414), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G22gat), .ZN(new_n420));
  INV_X1    g219(.A(G78gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n414), .A3(new_n415), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT31), .B(G50gat), .ZN(new_n424));
  INV_X1    g223(.A(G106gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n418), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n418), .B2(new_n423), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n266), .A2(new_n267), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n430), .B(KEYINPUT39), .C1(new_n267), .C2(new_n276), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n206), .C1(KEYINPUT39), .C2(new_n430), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT40), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT88), .B1(new_n278), .B2(new_n279), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT88), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n265), .A2(new_n272), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n207), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n433), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n376), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n374), .A2(new_n286), .A3(new_n375), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n440), .B1(new_n443), .B2(new_n393), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT37), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n363), .A2(new_n368), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n364), .B(new_n354), .C1(new_n361), .C2(new_n362), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n303), .B1(new_n366), .B2(new_n367), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT37), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT38), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n446), .A2(new_n449), .A3(new_n450), .A4(new_n372), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n438), .A2(new_n275), .A3(new_n281), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n284), .A4(new_n374), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n446), .A2(new_n372), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT37), .B1(new_n383), .B2(new_n386), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n450), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n429), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  OAI22_X1  g256(.A1(new_n397), .A2(new_n429), .B1(new_n444), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n232), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n351), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G227gat), .ZN(new_n461));
  INV_X1    g260(.A(G233gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n232), .B(new_n329), .C1(new_n348), .C2(new_n350), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G15gat), .B(G43gat), .Z(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n471), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n465), .B(KEYINPUT32), .C1(new_n467), .C2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT34), .ZN(new_n476));
  INV_X1    g275(.A(new_n463), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n232), .B1(new_n360), .B2(new_n329), .ZN(new_n478));
  INV_X1    g277(.A(new_n464), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT73), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT34), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n463), .B1(new_n460), .B2(new_n464), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT73), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n476), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT74), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n475), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n474), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT74), .B1(new_n491), .B2(new_n487), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n487), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT72), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n485), .B1(new_n484), .B2(new_n476), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n484), .A2(new_n476), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n491), .A2(new_n497), .B1(new_n500), .B2(new_n486), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n475), .A2(KEYINPUT72), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n492), .A2(new_n490), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n496), .B1(new_n503), .B2(new_n494), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n458), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n489), .B1(new_n475), .B2(new_n488), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n491), .A2(new_n487), .A3(KEYINPUT74), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n429), .B(new_n495), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT89), .B(KEYINPUT35), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n452), .B2(new_n284), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n443), .A2(new_n393), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n394), .A2(new_n396), .ZN(new_n513));
  INV_X1    g312(.A(new_n378), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n503), .A2(new_n513), .A3(new_n514), .A4(new_n429), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n512), .B1(new_n515), .B2(KEYINPUT35), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT90), .B1(new_n505), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n396), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n395), .B1(new_n389), .B2(new_n392), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n285), .B(new_n443), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n502), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n493), .A2(new_n521), .A3(new_n429), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT35), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n512), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n429), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n443), .A2(new_n393), .ZN(new_n528));
  INV_X1    g327(.A(new_n440), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n453), .A2(new_n456), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(new_n429), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n493), .A2(new_n521), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n527), .A2(new_n532), .A3(new_n534), .A4(new_n496), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n525), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(G197gat), .ZN(new_n539));
  XOR2_X1   g338(.A(KEYINPUT11), .B(G169gat), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT12), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G29gat), .ZN(new_n544));
  INV_X1    g343(.A(G36gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT14), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(G29gat), .B2(G36gat), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n546), .B(new_n548), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  XNOR2_X1  g351(.A(G43gat), .B(G50gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OR3_X1    g353(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559));
  INV_X1    g358(.A(G1gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT16), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(G1gat), .B2(new_n559), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G8gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n554), .A2(KEYINPUT17), .A3(new_n555), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n558), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n556), .A2(new_n564), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT18), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT91), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(KEYINPUT91), .A3(new_n571), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n556), .B(new_n564), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n568), .B(KEYINPUT13), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n567), .A2(KEYINPUT18), .A3(new_n568), .A4(new_n569), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT92), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n543), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n580), .B(KEYINPUT92), .Z(new_n583));
  AND3_X1   g382(.A1(new_n572), .A2(new_n542), .A3(new_n578), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT7), .ZN(new_n588));
  XNOR2_X1  g387(.A(G99gat), .B(G106gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(G99gat), .A2(G106gat), .ZN(new_n590));
  INV_X1    g389(.A(G85gat), .ZN(new_n591));
  INV_X1    g390(.A(G92gat), .ZN(new_n592));
  AOI22_X1  g391(.A1(KEYINPUT8), .A2(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n589), .B1(new_n588), .B2(new_n593), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n556), .A2(new_n596), .B1(KEYINPUT41), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n594), .A2(new_n595), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n558), .A2(new_n566), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT97), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n597), .A2(KEYINPUT41), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n607), .A2(KEYINPUT97), .A3(new_n613), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(G57gat), .A2(G64gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(G57gat), .A2(G64gat), .ZN(new_n619));
  AND2_X1   g418(.A1(G71gat), .A2(G78gat), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(KEYINPUT9), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(KEYINPUT93), .B2(new_n620), .ZN(new_n622));
  NOR2_X1   g421(.A1(G71gat), .A2(G78gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n626), .B(new_n621), .C1(KEYINPUT93), .C2(new_n620), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G127gat), .B(G155gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT20), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G183gat), .B(G211gat), .Z(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  AOI21_X1  g435(.A(new_n564), .B1(KEYINPUT21), .B2(new_n628), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n636), .B(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT98), .B1(new_n628), .B2(new_n596), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(new_n628), .B2(new_n596), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n601), .A2(KEYINPUT98), .A3(new_n625), .A4(new_n627), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G230gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n462), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n648), .A2(KEYINPUT100), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT10), .B1(new_n642), .B2(new_n643), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n628), .A2(new_n596), .A3(KEYINPUT10), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n628), .A2(new_n596), .A3(KEYINPUT99), .A4(KEYINPUT10), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n647), .B1(new_n650), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n648), .A2(KEYINPUT100), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n649), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n661), .B(new_n662), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n658), .A2(new_n659), .A3(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n617), .A2(new_n640), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n517), .A2(new_n537), .A3(new_n586), .A4(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n285), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n560), .ZN(G1324gat));
  NAND3_X1  g471(.A1(new_n517), .A2(new_n537), .A3(new_n586), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n528), .A3(new_n669), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(KEYINPUT102), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(G8gat), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  OR3_X1    g479(.A1(new_n675), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n676), .B2(new_n677), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n678), .B(new_n681), .C1(new_n682), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g482(.A(new_n504), .ZN(new_n684));
  OAI21_X1  g483(.A(G15gat), .B1(new_n670), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n493), .A2(new_n495), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n669), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n685), .B1(new_n673), .B2(new_n688), .ZN(G1326gat));
  NOR2_X1   g488(.A1(new_n670), .A2(new_n429), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  NAND3_X1  g491(.A1(new_n517), .A2(new_n537), .A3(new_n617), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT44), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT104), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT104), .B1(new_n523), .B2(new_n524), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n535), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n617), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT103), .B1(new_n582), .B2(new_n585), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n582), .A2(KEYINPUT103), .A3(new_n585), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n640), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n668), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n700), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n285), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n617), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n673), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n285), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n544), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n710), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n712), .A2(KEYINPUT45), .A3(new_n544), .A4(new_n714), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n709), .A2(new_n716), .A3(new_n717), .ZN(G1328gat));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  INV_X1    g518(.A(new_n528), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(G36gat), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n719), .B1(new_n713), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n712), .A2(KEYINPUT106), .A3(new_n721), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n708), .B2(new_n720), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n723), .A2(new_n725), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(KEYINPUT46), .ZN(new_n730));
  AOI211_X1 g529(.A(KEYINPUT107), .B(new_n724), .C1(new_n723), .C2(new_n725), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n726), .B(new_n727), .C1(new_n730), .C2(new_n731), .ZN(G1329gat));
  OAI21_X1  g531(.A(G43gat), .B1(new_n708), .B2(new_n684), .ZN(new_n733));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n712), .A2(new_n734), .A3(new_n687), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1330gat));
  OAI21_X1  g539(.A(G50gat), .B1(new_n708), .B2(new_n429), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n713), .A2(G50gat), .A3(new_n429), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n741), .A2(new_n743), .A3(new_n745), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1331gat));
  NOR4_X1   g548(.A1(new_n705), .A2(new_n617), .A3(new_n640), .A4(new_n667), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n697), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n714), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  INV_X1    g552(.A(new_n751), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n720), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  NAND2_X1  g558(.A1(new_n751), .A2(new_n687), .ZN(new_n760));
  AOI21_X1  g559(.A(G71gat), .B1(new_n760), .B2(KEYINPUT109), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(KEYINPUT109), .B2(new_n760), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n751), .A2(G71gat), .A3(new_n504), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT50), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n762), .A2(new_n766), .A3(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1334gat));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n526), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G78gat), .ZN(G1335gat));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n705), .A2(new_n706), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n668), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n700), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n771), .B1(new_n775), .B2(new_n285), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n773), .B1(new_n694), .B2(new_n699), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(KEYINPUT110), .A3(new_n714), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(G85gat), .A3(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n697), .A2(new_n617), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT51), .B1(new_n780), .B2(new_n772), .ZN(new_n781));
  AND4_X1   g580(.A1(KEYINPUT51), .A2(new_n697), .A3(new_n617), .A4(new_n772), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n668), .A2(new_n591), .A3(new_n714), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n779), .B1(new_n783), .B2(new_n784), .ZN(G1336gat));
  OAI21_X1  g584(.A(KEYINPUT111), .B1(new_n775), .B2(new_n720), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n777), .A2(new_n787), .A3(new_n528), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(G92gat), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n781), .A2(new_n782), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n720), .A2(new_n667), .A3(G92gat), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n791), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n783), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n592), .B1(new_n777), .B2(new_n528), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT52), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n775), .B2(new_n684), .ZN(new_n799));
  INV_X1    g598(.A(G99gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n687), .A2(new_n668), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n783), .B2(new_n801), .ZN(G1338gat));
  NOR3_X1   g601(.A1(new_n667), .A2(G106gat), .A3(new_n429), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n781), .B2(new_n782), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n425), .B1(new_n777), .B2(new_n526), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g606(.A(KEYINPUT112), .B(new_n425), .C1(new_n777), .C2(new_n526), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT53), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n805), .A2(KEYINPUT53), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n804), .A2(KEYINPUT113), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n803), .C1(new_n781), .C2(new_n782), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n809), .A2(new_n814), .ZN(G1339gat));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816));
  INV_X1    g615(.A(new_n703), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT10), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n644), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n655), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n820), .A3(new_n646), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(KEYINPUT54), .A3(new_n656), .ZN(new_n822));
  XNOR2_X1  g621(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n647), .B(new_n823), .C1(new_n650), .C2(new_n655), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n664), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n649), .A2(new_n657), .A3(new_n656), .A4(new_n663), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n664), .A4(new_n824), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n817), .A2(new_n830), .A3(new_n701), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n576), .A2(new_n577), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT116), .Z(new_n833));
  NAND2_X1  g632(.A1(new_n567), .A2(new_n569), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(G229gat), .A3(G233gat), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(KEYINPUT115), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n838), .A2(new_n541), .B1(new_n583), .B2(new_n584), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n839), .A2(new_n665), .A3(new_n666), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n816), .B1(new_n831), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n615), .A2(new_n616), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(new_n665), .A3(new_n666), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT117), .B(new_n843), .C1(new_n704), .C2(new_n830), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n830), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n617), .A2(new_n846), .A3(new_n839), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n706), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NOR4_X1   g647(.A1(new_n705), .A2(new_n617), .A3(new_n640), .A4(new_n668), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n508), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n528), .A2(new_n285), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n586), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n222), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n522), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n850), .A2(new_n714), .A3(new_n856), .A4(new_n720), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(new_n704), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n855), .B1(new_n858), .B2(new_n222), .ZN(G1340gat));
  OAI21_X1  g658(.A(new_n220), .B1(new_n857), .B2(new_n667), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n668), .A2(G120gat), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n853), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT118), .ZN(G1341gat));
  OAI21_X1  g662(.A(G127gat), .B1(new_n853), .B2(new_n640), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n706), .A2(new_n213), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n857), .B2(new_n865), .ZN(G1342gat));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n714), .A3(new_n856), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n842), .A2(new_n528), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n211), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n867), .A2(KEYINPUT56), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G134gat), .B1(new_n853), .B2(new_n842), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT56), .B1(new_n867), .B2(new_n869), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G1343gat));
  NOR2_X1   g672(.A1(new_n504), .A2(new_n429), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n850), .A2(new_n714), .A3(new_n720), .A4(new_n874), .ZN(new_n875));
  OR3_X1    g674(.A1(new_n875), .A2(G141gat), .A3(new_n854), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n684), .A2(new_n852), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n843), .B1(new_n854), .B2(new_n830), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n842), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n706), .B1(new_n880), .B2(new_n847), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n526), .B1(new_n881), .B2(new_n849), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n878), .B1(new_n882), .B2(KEYINPUT57), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n884), .B(new_n526), .C1(new_n848), .C2(new_n849), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT120), .B1(new_n886), .B2(new_n854), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G141gat), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n886), .A2(KEYINPUT120), .A3(new_n854), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n876), .B(new_n877), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n883), .A2(new_n885), .A3(new_n705), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n891), .A2(KEYINPUT119), .A3(G141gat), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n875), .A2(G141gat), .A3(new_n854), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT119), .B1(new_n891), .B2(G141gat), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n890), .B1(new_n895), .B2(new_n877), .ZN(G1344gat));
  NOR3_X1   g695(.A1(new_n886), .A2(KEYINPUT59), .A3(new_n667), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT59), .B1(new_n875), .B2(new_n667), .ZN(new_n898));
  INV_X1    g697(.A(G148gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT57), .B(new_n526), .C1(new_n848), .C2(new_n849), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n669), .A2(new_n854), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n526), .B1(new_n903), .B2(new_n881), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n884), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n902), .A2(new_n901), .ZN(new_n908));
  AOI211_X1 g707(.A(new_n667), .B(new_n878), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n900), .B1(new_n909), .B2(new_n910), .ZN(G1345gat));
  OAI21_X1  g710(.A(G155gat), .B1(new_n886), .B2(new_n640), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n706), .A2(new_n248), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n875), .B2(new_n913), .ZN(G1346gat));
  NOR2_X1   g713(.A1(new_n848), .A2(new_n849), .ZN(new_n915));
  INV_X1    g714(.A(new_n874), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n868), .A2(new_n249), .ZN(new_n917));
  NOR4_X1   g716(.A1(new_n915), .A2(new_n285), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT122), .ZN(new_n919));
  OAI21_X1  g718(.A(G162gat), .B1(new_n886), .B2(new_n842), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1347gat));
  NAND2_X1  g720(.A1(new_n856), .A2(new_n528), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT123), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n285), .B(new_n923), .C1(new_n848), .C2(new_n849), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n705), .A2(new_n311), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT124), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n528), .A2(new_n285), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT125), .Z(new_n929));
  NAND3_X1  g728(.A1(new_n850), .A2(new_n851), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n854), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n927), .A2(KEYINPUT126), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1348gat));
  OAI21_X1  g735(.A(G176gat), .B1(new_n930), .B2(new_n667), .ZN(new_n937));
  INV_X1    g736(.A(new_n924), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n312), .A3(new_n668), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1349gat));
  OAI21_X1  g739(.A(G183gat), .B1(new_n930), .B2(new_n640), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n336), .A3(new_n706), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n938), .A2(new_n337), .A3(new_n617), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n850), .A2(new_n851), .A3(new_n617), .A4(new_n929), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n946), .A2(new_n947), .A3(G190gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n946), .B2(G190gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT127), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n952), .B(new_n945), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1351gat));
  NOR2_X1   g753(.A1(new_n915), .A2(new_n714), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n916), .A2(new_n720), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n705), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n929), .A2(new_n684), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n960), .B1(new_n907), .B2(new_n908), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n854), .A2(new_n293), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1352gat));
  NAND4_X1  g762(.A1(new_n955), .A2(new_n295), .A3(new_n668), .A4(new_n956), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT62), .Z(new_n965));
  INV_X1    g764(.A(new_n960), .ZN(new_n966));
  INV_X1    g765(.A(new_n908), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n668), .B(new_n966), .C1(new_n967), .C2(new_n906), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n965), .B1(new_n295), .B2(new_n969), .ZN(G1353gat));
  OR3_X1    g769(.A1(new_n957), .A2(G211gat), .A3(new_n640), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n706), .B(new_n966), .C1(new_n967), .C2(new_n906), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  INV_X1    g774(.A(G218gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n976), .A3(new_n617), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n617), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n977), .B1(new_n979), .B2(new_n976), .ZN(G1355gat));
endmodule


