//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1193, new_n1194, new_n1195,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  AND3_X1   g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT67), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n219), .B(new_n220), .C1(new_n215), .C2(new_n216), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT69), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n209), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(G250), .B1(G257), .B2(G264), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT0), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n230), .A2(G50), .A3(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n207), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n228), .A2(KEYINPUT0), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n229), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  OAI21_X1  g0039(.A(new_n239), .B1(KEYINPUT1), .B2(new_n222), .ZN(new_n240));
  NOR2_X1   g0040(.A1(new_n224), .A2(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  INV_X1    g0042(.A(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT2), .B(G226), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G264), .B(G270), .Z(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT70), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(G68), .B(G77), .Z(new_n255));
  XOR2_X1   g0055(.A(G50), .B(G58), .Z(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n254), .B(new_n257), .Z(G351));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n234), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n207), .B1(new_n201), .B2(new_n203), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n207), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n262), .A2(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n260), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G13), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n269), .A2(new_n207), .A3(G1), .ZN(new_n270));
  INV_X1    g0070(.A(G50), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n270), .A2(new_n260), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n206), .A2(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n268), .B(new_n272), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G222), .A2(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G223), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n234), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n283), .B(new_n287), .C1(G77), .C2(new_n279), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(new_n284), .B2(new_n285), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT71), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(new_n294), .B2(new_n206), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G41), .A2(G45), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n296), .A2(KEYINPUT71), .A3(G1), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n290), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n286), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G226), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n288), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n277), .A2(new_n278), .B1(G200), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n303), .B1(new_n278), .B2(new_n277), .C1(new_n304), .C2(new_n302), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT10), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n302), .A2(G179), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT72), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n277), .A3(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT75), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n275), .A2(G77), .ZN(new_n314));
  INV_X1    g0114(.A(new_n270), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n274), .A2(new_n314), .B1(G77), .B2(new_n315), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n262), .A2(new_n266), .B1(new_n207), .B2(new_n202), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT15), .B(G87), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n263), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n260), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT74), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(KEYINPUT74), .B(new_n260), .C1(new_n317), .C2(new_n319), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n316), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(G232), .A2(G1698), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n281), .A2(G238), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n279), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(new_n287), .C1(G107), .C2(new_n279), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n300), .A2(G244), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n298), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n309), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n329), .A2(new_n333), .A3(new_n330), .A4(new_n298), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n325), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n330), .A2(new_n298), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n336), .A2(KEYINPUT73), .A3(G190), .A4(new_n329), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT73), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n331), .B2(G200), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n331), .A2(new_n304), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n324), .B(new_n337), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n312), .A2(new_n313), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n313), .B1(new_n312), .B2(new_n342), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n262), .B1(new_n206), .B2(G20), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(new_n273), .B1(new_n270), .B2(new_n262), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G33), .ZN(new_n348));
  INV_X1    g0148(.A(G33), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT7), .B1(new_n351), .B2(new_n207), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  AOI211_X1 g0153(.A(new_n353), .B(G20), .C1(new_n348), .C2(new_n350), .ZN(new_n354));
  OAI21_X1  g0154(.A(G68), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G58), .ZN(new_n356));
  INV_X1    g0156(.A(G68), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(G20), .B1(new_n358), .B2(new_n203), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n265), .A2(G159), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n355), .A2(KEYINPUT16), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n260), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT78), .B1(new_n349), .B2(KEYINPUT3), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT78), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(new_n347), .A3(G33), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n367), .A3(new_n350), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n353), .A2(G20), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n353), .B1(new_n279), .B2(G20), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G68), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT16), .B1(new_n373), .B2(new_n362), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n346), .B1(new_n364), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT81), .ZN(new_n376));
  INV_X1    g0176(.A(G223), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(G1698), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT79), .B1(new_n279), .B2(new_n378), .ZN(new_n379));
  AND4_X1   g0179(.A1(KEYINPUT79), .A2(new_n378), .A3(new_n348), .A4(new_n350), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n348), .A2(new_n350), .A3(G226), .A4(G1698), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G87), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n286), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n286), .A2(G232), .A3(new_n299), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n298), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n376), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n378), .A2(new_n348), .A3(new_n350), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT79), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n378), .A2(new_n348), .A3(new_n350), .A4(KEYINPUT79), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n391), .A2(new_n383), .A3(new_n382), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n287), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n298), .A2(new_n386), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(KEYINPUT81), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(G200), .B1(new_n388), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n387), .B1(new_n287), .B2(new_n393), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n304), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT82), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G200), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n394), .A2(KEYINPUT81), .A3(new_n395), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT81), .B1(new_n394), .B2(new_n395), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT82), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n399), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n375), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g0208(.A(KEYINPUT83), .B(KEYINPUT17), .Z(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(KEYINPUT83), .A2(KEYINPUT17), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n411), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  AOI21_X1  g0214(.A(G169), .B1(new_n388), .B2(new_n396), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n394), .A2(new_n333), .A3(new_n395), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT80), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT80), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n398), .A2(new_n418), .A3(new_n333), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n414), .B1(new_n421), .B2(new_n375), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(new_n398), .B2(new_n333), .ZN(new_n423));
  AND4_X1   g0223(.A1(new_n418), .A2(new_n394), .A3(new_n333), .A4(new_n395), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n309), .B1(new_n403), .B2(new_n404), .ZN(new_n426));
  AND4_X1   g0226(.A1(new_n414), .A2(new_n425), .A3(new_n375), .A4(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n413), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n299), .B(KEYINPUT71), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n290), .A2(new_n430), .B1(new_n300), .B2(G238), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G97), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n243), .A2(G1698), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G226), .B2(G1698), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n432), .B1(new_n434), .B2(new_n351), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n287), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT13), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G169), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT14), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT14), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n441), .A3(G169), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT13), .ZN(new_n443));
  OR3_X1    g0243(.A1(new_n437), .A2(KEYINPUT76), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n437), .B1(KEYINPUT76), .B2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G179), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n270), .A2(new_n357), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT12), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n273), .A2(G68), .A3(new_n275), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n263), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT77), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n452), .A2(new_n453), .B1(new_n271), .B2(new_n266), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n260), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT11), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n450), .B(new_n451), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n456), .A2(new_n457), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n448), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n438), .A2(G200), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n460), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n304), .B1(new_n444), .B2(new_n445), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  NOR4_X1   g0268(.A1(new_n343), .A2(new_n344), .A3(new_n429), .A4(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n265), .A2(G77), .ZN(new_n471));
  XOR2_X1   g0271(.A(new_n471), .B(KEYINPUT84), .Z(new_n472));
  INV_X1    g0272(.A(G97), .ZN(new_n473));
  INV_X1    g0273(.A(G107), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT6), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(KEYINPUT6), .B2(new_n473), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT85), .B(G107), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n476), .B(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n472), .B1(new_n478), .B2(new_n207), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n474), .B1(new_n370), .B2(new_n371), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n260), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n315), .A2(G97), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n273), .B1(G1), .B2(new_n349), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n482), .B1(new_n484), .B2(G97), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n293), .A2(G1), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G257), .A3(new_n286), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n290), .A2(new_n489), .A3(new_n488), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(KEYINPUT87), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT87), .B1(new_n491), .B2(new_n492), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n281), .A2(G244), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n351), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G283), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n499), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n287), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(KEYINPUT86), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT86), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n503), .B2(new_n287), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n496), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G200), .ZN(new_n509));
  INV_X1    g0309(.A(new_n495), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n493), .A3(new_n504), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT88), .B1(new_n512), .B2(G190), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT88), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n511), .A2(new_n514), .A3(new_n304), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n487), .B(new_n509), .C1(new_n513), .C2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n496), .B(new_n333), .C1(new_n505), .C2(new_n507), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n511), .A2(new_n309), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n486), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n279), .A2(new_n207), .A3(G68), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT19), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n207), .B1(new_n432), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G87), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(new_n473), .A3(new_n474), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n521), .B1(new_n263), .B2(new_n473), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n260), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n318), .A2(new_n270), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT89), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n528), .A2(KEYINPUT89), .A3(new_n529), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n532), .A2(new_n533), .B1(G87), .B2(new_n484), .ZN(new_n534));
  INV_X1    g0334(.A(G250), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n489), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n290), .A2(new_n489), .B1(new_n536), .B2(new_n286), .ZN(new_n537));
  MUX2_X1   g0337(.A(G238), .B(G244), .S(G1698), .Z(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(new_n279), .B1(G33), .B2(G116), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n539), .B2(new_n286), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n304), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(G200), .B2(new_n540), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n528), .A2(KEYINPUT89), .A3(new_n529), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT89), .B1(new_n528), .B2(new_n529), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n543), .A2(new_n544), .B1(new_n318), .B2(new_n483), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n540), .A2(G179), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n309), .B2(new_n540), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n534), .A2(new_n542), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n516), .A2(new_n519), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n281), .A2(G250), .ZN(new_n550));
  INV_X1    g0350(.A(G294), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n351), .A2(new_n550), .B1(new_n349), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n279), .A2(G257), .A3(G1698), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT93), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n279), .A2(KEYINPUT93), .A3(G257), .A4(G1698), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n557), .A2(new_n286), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n490), .A2(G264), .A3(new_n286), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n558), .A2(new_n333), .A3(new_n492), .A4(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n492), .B(new_n559), .C1(new_n557), .C2(new_n286), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n309), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n279), .A2(new_n207), .A3(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT22), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT22), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n279), .A2(new_n565), .A3(new_n207), .A4(G87), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n474), .A3(G20), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT92), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n568), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n572), .B2(new_n571), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g0375(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n576), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n567), .A2(new_n578), .A3(new_n574), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n577), .A2(new_n579), .B1(new_n234), .B2(new_n259), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT25), .B1(new_n270), .B2(new_n474), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n474), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n483), .A2(new_n474), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n560), .B(new_n562), .C1(new_n580), .C2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n273), .B(G116), .C1(G1), .C2(new_n349), .ZN(new_n586));
  INV_X1    g0386(.A(G116), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n270), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n259), .A2(new_n234), .B1(G20), .B2(new_n587), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n501), .B(new_n207), .C1(G33), .C2(new_n473), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT20), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n589), .A2(KEYINPUT20), .A3(new_n590), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n586), .B(new_n588), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n351), .A2(new_n594), .ZN(new_n595));
  MUX2_X1   g0395(.A(G257), .B(G264), .S(G1698), .Z(new_n596));
  OAI211_X1 g0396(.A(new_n595), .B(new_n287), .C1(new_n351), .C2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n490), .A2(G270), .A3(new_n286), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n492), .A3(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n593), .A2(KEYINPUT21), .A3(new_n599), .A4(G169), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n599), .A2(new_n333), .ZN(new_n601));
  INV_X1    g0401(.A(new_n593), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n599), .A2(G169), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT21), .B1(new_n604), .B2(new_n593), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n585), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n599), .A2(G200), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n602), .B(new_n608), .C1(new_n304), .C2(new_n599), .ZN(new_n609));
  XOR2_X1   g0409(.A(new_n609), .B(KEYINPUT90), .Z(new_n610));
  NAND2_X1  g0410(.A1(new_n577), .A2(new_n579), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n260), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n561), .A2(new_n304), .ZN(new_n613));
  INV_X1    g0413(.A(new_n584), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n561), .A2(G200), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n612), .A2(new_n613), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n470), .A2(new_n549), .A3(new_n607), .A4(new_n617), .ZN(G372));
  NAND2_X1  g0418(.A1(new_n545), .A2(new_n547), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n607), .A2(new_n616), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n549), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n534), .A2(new_n542), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n619), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n622), .B1(new_n624), .B2(new_n519), .ZN(new_n625));
  INV_X1    g0425(.A(new_n519), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n548), .A3(KEYINPUT26), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n469), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n462), .B1(new_n466), .B2(new_n335), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n631), .A2(new_n413), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT94), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n422), .B2(new_n427), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n421), .A2(new_n414), .A3(new_n375), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n426), .A2(new_n375), .A3(new_n419), .A4(new_n417), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT18), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n637), .A3(KEYINPUT94), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n306), .B1(new_n632), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(new_n311), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n630), .A2(new_n641), .ZN(G369));
  NAND3_X1  g0442(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n602), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n606), .B1(new_n610), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT96), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT95), .B1(new_n602), .B2(new_n649), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G330), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n648), .B1(new_n580), .B2(new_n584), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n616), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n585), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n585), .A2(new_n648), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n585), .A2(new_n648), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n606), .A2(new_n648), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n664), .B1(new_n658), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(G399));
  NOR2_X1   g0467(.A1(new_n226), .A2(G41), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n524), .A2(G116), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G1), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n232), .B2(new_n669), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT97), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n628), .A2(new_n674), .ZN(new_n675));
  OAI221_X1 g0475(.A(new_n619), .B1(new_n627), .B2(new_n674), .C1(new_n549), .C2(new_n620), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n649), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n677), .A2(KEYINPUT29), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n629), .A2(new_n679), .A3(new_n649), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NOR4_X1   g0482(.A1(new_n617), .A2(new_n549), .A3(new_n607), .A4(new_n648), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n558), .A2(new_n559), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n601), .A2(new_n540), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(new_n512), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT30), .A4(new_n512), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n599), .A2(new_n540), .A3(new_n333), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n508), .A2(new_n561), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n648), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT31), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n684), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n682), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n673), .B1(new_n699), .B2(G1), .ZN(G364));
  NOR2_X1   g0500(.A1(new_n269), .A2(G20), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n206), .B1(new_n701), .B2(G45), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n668), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n654), .B2(G330), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(G330), .B2(new_n654), .ZN(new_n706));
  NOR2_X1   g0506(.A1(G13), .A2(G33), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G20), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT100), .Z(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n284), .B1(new_n207), .B2(G169), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT101), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n225), .A2(new_n351), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT99), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n257), .A2(G45), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT98), .Z(new_n718));
  AOI211_X1 g0518(.A(new_n716), .B(new_n718), .C1(new_n293), .C2(new_n233), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n225), .A2(new_n279), .ZN(new_n720));
  INV_X1    g0520(.A(G355), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n720), .A2(new_n721), .B1(G116), .B2(new_n225), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n714), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n304), .A2(G179), .A3(G200), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n207), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n473), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n207), .A2(new_n333), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G200), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n304), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n726), .B1(G50), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT32), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n207), .A2(G179), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G190), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G159), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n732), .A2(new_n304), .A3(G200), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n730), .B1(new_n731), .B2(new_n736), .C1(new_n474), .C2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n732), .A2(G190), .A3(G200), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G87), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n731), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n728), .A2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n741), .B(new_n742), .C1(new_n744), .C2(new_n357), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n727), .A2(new_n733), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n727), .A2(G190), .A3(new_n402), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n279), .B1(new_n746), .B2(new_n202), .C1(new_n356), .C2(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n738), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n747), .ZN(new_n750));
  INV_X1    g0550(.A(new_n734), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n750), .A2(G322), .B1(new_n751), .B2(G329), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n752), .B(new_n351), .C1(new_n753), .C2(new_n746), .ZN(new_n754));
  INV_X1    g0554(.A(G317), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n743), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n729), .A2(G326), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n758), .B(new_n759), .C1(new_n594), .C2(new_n739), .ZN(new_n760));
  INV_X1    g0560(.A(G283), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n725), .A2(new_n551), .B1(new_n737), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n754), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n713), .B1(new_n749), .B2(new_n763), .ZN(new_n764));
  AND3_X1   g0564(.A1(new_n723), .A2(new_n764), .A3(new_n704), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n654), .B2(new_n710), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n706), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(G396));
  INV_X1    g0568(.A(new_n704), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n713), .A2(new_n707), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(new_n202), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT105), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n332), .A2(new_n334), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n324), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n649), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n325), .A2(new_n648), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n341), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n772), .B(new_n775), .C1(new_n777), .C2(new_n774), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n774), .B1(new_n341), .B2(new_n776), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n335), .A2(new_n648), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT105), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n746), .A2(new_n587), .B1(new_n734), .B2(new_n753), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G294), .B2(new_n750), .ZN(new_n784));
  INV_X1    g0584(.A(new_n729), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n785), .A2(new_n594), .B1(new_n737), .B2(new_n523), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n726), .B(new_n786), .C1(G283), .C2(new_n743), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n351), .B1(new_n739), .B2(new_n474), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT102), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  AND4_X1   g0591(.A1(new_n784), .A2(new_n787), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n746), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n750), .A2(G143), .B1(new_n793), .B2(G159), .ZN(new_n794));
  INV_X1    g0594(.A(G137), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n794), .B1(new_n744), .B2(new_n264), .C1(new_n795), .C2(new_n785), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT34), .ZN(new_n797));
  INV_X1    g0597(.A(new_n737), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G68), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n271), .B2(new_n739), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n800), .A2(KEYINPUT103), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(KEYINPUT103), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n279), .B1(new_n734), .B2(new_n803), .C1(new_n725), .C2(new_n356), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n792), .B1(new_n797), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT104), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n713), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n806), .A2(KEYINPUT104), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n771), .B1(new_n782), .B2(new_n708), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n629), .A2(new_n649), .ZN(new_n811));
  INV_X1    g0611(.A(new_n782), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n649), .B(new_n782), .C1(new_n621), .C2(new_n628), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n697), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n697), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n704), .B(new_n816), .C1(KEYINPUT106), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(KEYINPUT106), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n810), .B1(new_n819), .B2(new_n820), .ZN(G384));
  NOR2_X1   g0621(.A1(new_n701), .A2(new_n206), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT39), .ZN(new_n823));
  INV_X1    g0623(.A(new_n375), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n646), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT37), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n636), .A2(new_n826), .ZN(new_n827));
  OR3_X1    g0627(.A1(new_n408), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n636), .A2(KEYINPUT94), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n425), .A2(new_n633), .A3(new_n426), .A4(new_n375), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n831), .A2(new_n408), .A3(new_n825), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n828), .B1(new_n832), .B2(new_n826), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n408), .A2(new_n412), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n375), .B(new_n409), .C1(new_n401), .C2(new_n407), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n634), .B(new_n638), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n833), .A2(KEYINPUT110), .B1(new_n825), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT110), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n828), .B(new_n838), .C1(new_n832), .C2(new_n826), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT38), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n408), .A2(new_n825), .A3(new_n827), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT108), .ZN(new_n842));
  INV_X1    g0642(.A(new_n346), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n351), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n371), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n361), .B1(new_n845), .B2(G68), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n260), .B1(new_n846), .B2(KEYINPUT16), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT107), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n847), .A2(new_n848), .B1(KEYINPUT16), .B2(new_n846), .ZN(new_n849));
  OAI211_X1 g0649(.A(KEYINPUT107), .B(new_n260), .C1(new_n846), .C2(KEYINPUT16), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n843), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n851), .A2(new_n415), .A3(new_n420), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n842), .B1(new_n408), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n397), .A2(KEYINPUT82), .A3(new_n400), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n406), .B1(new_n405), .B2(new_n399), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n824), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n851), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n421), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n856), .A2(new_n858), .A3(KEYINPUT108), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n851), .A2(new_n646), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n853), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n841), .B1(new_n862), .B2(KEYINPUT37), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n861), .B1(new_n413), .B2(new_n428), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n823), .B1(new_n840), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n448), .A2(new_n461), .A3(new_n649), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n828), .ZN(new_n871));
  INV_X1    g0671(.A(new_n865), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT39), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n867), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n814), .A2(new_n775), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n462), .B(new_n467), .C1(new_n460), .C2(new_n649), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n461), .B(new_n648), .C1(new_n448), .C2(new_n466), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n871), .B2(new_n872), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(new_n866), .ZN(new_n884));
  INV_X1    g0684(.A(new_n639), .ZN(new_n885));
  INV_X1    g0685(.A(new_n646), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(KEYINPUT109), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT109), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n881), .B1(new_n873), .B2(new_n874), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n887), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n876), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT111), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n876), .A2(new_n889), .A3(new_n892), .A4(KEYINPUT111), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n469), .B1(new_n678), .B2(new_n681), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n641), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT112), .Z(new_n900));
  XNOR2_X1  g0700(.A(new_n897), .B(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT31), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n694), .B(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n880), .B(new_n782), .C1(new_n904), .C2(new_n683), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n902), .B(new_n906), .C1(new_n883), .C2(new_n866), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n408), .A2(new_n825), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n829), .A2(new_n830), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n826), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT110), .B1(new_n910), .B2(new_n841), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n836), .A2(new_n825), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(new_n839), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n864), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n905), .B1(new_n914), .B2(new_n873), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n907), .B1(new_n915), .B2(new_n902), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n469), .A2(new_n696), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(G330), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n822), .B1(new_n901), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n901), .B2(new_n920), .ZN(new_n922));
  INV_X1    g0722(.A(new_n478), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n923), .A2(KEYINPUT35), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(KEYINPUT35), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n924), .A2(G116), .A3(new_n235), .A4(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT36), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n232), .A2(new_n202), .A3(new_n358), .ZN(new_n928));
  INV_X1    g0728(.A(new_n201), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n357), .ZN(new_n930));
  OAI211_X1 g0730(.A(G1), .B(new_n269), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n922), .A2(new_n927), .A3(new_n931), .ZN(G367));
  OAI21_X1  g0732(.A(new_n714), .B1(new_n225), .B2(new_n318), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n716), .A2(new_n249), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n704), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT115), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n534), .A2(new_n649), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n548), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n619), .B2(new_n937), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n351), .B1(new_n734), .B2(new_n755), .C1(new_n747), .C2(new_n594), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n740), .A2(KEYINPUT46), .A3(G116), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT46), .B1(new_n740), .B2(G116), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n744), .A2(new_n551), .B1(new_n737), .B2(new_n473), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(G311), .B2(new_n729), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n725), .A2(new_n474), .B1(new_n746), .B2(new_n761), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT116), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(KEYINPUT116), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n737), .A2(new_n202), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n351), .B(new_n951), .C1(G137), .C2(new_n751), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n356), .B2(new_n739), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n743), .A2(G159), .B1(new_n929), .B2(new_n793), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(KEYINPUT118), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(KEYINPUT118), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(G143), .A2(new_n729), .B1(new_n750), .B2(G150), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n357), .B2(new_n725), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT117), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n943), .A2(new_n950), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT47), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n713), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n962), .A2(KEYINPUT47), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n936), .B1(new_n939), .B2(new_n710), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n516), .B(new_n519), .C1(new_n487), .C2(new_n649), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n626), .A2(new_n648), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n666), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT45), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n969), .A2(new_n666), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT44), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n662), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT114), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n660), .B(new_n665), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n655), .B(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(new_n698), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n662), .A2(new_n974), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n699), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT113), .B(KEYINPUT41), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n668), .B(new_n983), .Z(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n703), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n969), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n663), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n967), .A2(new_n585), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n648), .B1(new_n989), .B2(new_n519), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n660), .A2(new_n969), .A3(new_n665), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n990), .B1(KEYINPUT42), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(KEYINPUT42), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n992), .A2(new_n993), .B1(KEYINPUT43), .B2(new_n939), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n988), .B(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n966), .B1(new_n986), .B2(new_n997), .ZN(G387));
  OAI22_X1  g0798(.A1(new_n720), .A2(new_n670), .B1(G107), .B2(new_n225), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n246), .A2(new_n293), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n262), .A2(G50), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT50), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n670), .ZN(new_n1003));
  AOI211_X1 g0803(.A(G45), .B(new_n1003), .C1(G68), .C2(G77), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n716), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n999), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n714), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n704), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT119), .Z(new_n1009));
  OAI22_X1  g0809(.A1(new_n746), .A2(new_n357), .B1(new_n734), .B2(new_n264), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n351), .B(new_n1010), .C1(G50), .C2(new_n750), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n740), .A2(G77), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n318), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n725), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n262), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1013), .A2(new_n1014), .B1(new_n743), .B2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n729), .A2(G159), .B1(new_n798), .B2(G97), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1011), .A2(new_n1012), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n279), .B1(new_n751), .B2(G326), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n725), .A2(new_n761), .B1(new_n739), .B2(new_n551), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n750), .A2(G317), .B1(new_n793), .B2(G303), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n729), .A2(G322), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n753), .C2(new_n744), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1024), .B2(new_n1023), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT49), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1019), .B1(new_n587), .B2(new_n737), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1018), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n713), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1009), .B(new_n1031), .C1(new_n660), .C2(new_n710), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n978), .A2(new_n698), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n668), .B1(new_n978), .B2(new_n698), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1032), .B1(new_n702), .B2(new_n978), .C1(new_n1033), .C2(new_n1034), .ZN(G393));
  AND2_X1   g0835(.A1(new_n980), .A2(new_n975), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n668), .B1(new_n1036), .B2(new_n979), .C1(new_n981), .C2(new_n976), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G150), .A2(new_n729), .B1(new_n750), .B2(G159), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT51), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n740), .A2(G68), .B1(new_n751), .B2(G143), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT120), .Z(new_n1041));
  NOR2_X1   g0841(.A1(new_n744), .A2(new_n201), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n279), .B1(new_n746), .B2(new_n262), .C1(new_n523), .C2(new_n737), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n725), .A2(new_n202), .ZN(new_n1044));
  OR3_X1    g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1039), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G317), .A2(new_n729), .B1(new_n750), .B2(G311), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT52), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n279), .B1(new_n751), .B2(G322), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n551), .B2(new_n746), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n744), .A2(new_n594), .B1(new_n737), .B2(new_n474), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n725), .A2(new_n587), .B1(new_n739), .B2(new_n761), .ZN(new_n1052));
  NOR4_X1   g0852(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n713), .B1(new_n1046), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n254), .A2(new_n716), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n714), .B1(new_n473), .B2(new_n225), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1054), .B(new_n704), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n987), .B2(new_n711), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1036), .B2(new_n703), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1037), .A2(new_n1059), .ZN(G390));
  NAND2_X1  g0860(.A1(new_n867), .A2(new_n875), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n881), .A2(new_n868), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n868), .B(KEYINPUT121), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n775), .B1(new_n677), .B2(new_n812), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n880), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n914), .A2(new_n873), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n812), .B1(new_n684), .B2(new_n695), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1069), .A2(G330), .A3(new_n880), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1063), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1061), .A2(new_n1062), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT122), .ZN(new_n1073));
  OAI211_X1 g0873(.A(G330), .B(new_n782), .C1(new_n904), .C2(new_n683), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n880), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1069), .A2(KEYINPUT122), .A3(G330), .A4(new_n880), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1071), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n469), .A2(G330), .A3(new_n696), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n898), .A2(new_n1080), .A3(new_n641), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n877), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1070), .A2(new_n1082), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(new_n1065), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1081), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1079), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1087), .B(new_n1071), .C1(new_n1072), .C2(new_n1078), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n668), .A3(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1071), .B(new_n703), .C1(new_n1072), .C2(new_n1078), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1061), .A2(new_n707), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n770), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n704), .B1(new_n1094), .B2(new_n1015), .ZN(new_n1095));
  INV_X1    g0895(.A(G125), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n279), .B1(new_n734), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n744), .A2(new_n795), .B1(new_n201), .B2(new_n737), .ZN(new_n1098));
  INV_X1    g0898(.A(G128), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n785), .A2(new_n1099), .B1(new_n735), .B2(new_n725), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT54), .B(G143), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n747), .A2(new_n803), .B1(new_n746), .B2(new_n1101), .ZN(new_n1102));
  OR4_X1    g0902(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n740), .A2(G150), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT53), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1044), .B1(G283), .B2(new_n729), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n474), .B2(new_n744), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n747), .A2(new_n587), .B1(new_n734), .B2(new_n551), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n279), .B(new_n1108), .C1(G97), .C2(new_n793), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n741), .A3(new_n799), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1103), .A2(new_n1105), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1095), .B1(new_n1111), .B2(new_n713), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1093), .A2(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1092), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1091), .A2(new_n1114), .ZN(G378));
  NAND2_X1  g0915(.A1(new_n277), .A2(new_n886), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n312), .B(new_n1116), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1118));
  XNOR2_X1  g0918(.A(new_n1117), .B(new_n1118), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n916), .A2(G330), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n916), .B2(G330), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n897), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n895), .B(new_n896), .C1(new_n1121), .C2(new_n1120), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(KEYINPUT123), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1081), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1090), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT123), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n897), .A2(new_n1122), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT57), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1090), .B2(new_n1126), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n669), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1125), .A2(new_n703), .A3(new_n1129), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n704), .B1(new_n1094), .B2(new_n929), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n798), .A2(G58), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n744), .B2(new_n473), .C1(new_n587), .C2(new_n785), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n292), .B(new_n351), .C1(new_n734), .C2(new_n761), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n747), .A2(new_n474), .B1(new_n746), .B2(new_n318), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1012), .B1(new_n357), .B2(new_n725), .ZN(new_n1143));
  OR4_X1    g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT58), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(G50), .B1(new_n349), .B2(new_n292), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n279), .B2(G41), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n744), .A2(new_n803), .B1(new_n785), .B2(new_n1096), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n750), .A2(G128), .B1(new_n793), .B2(G137), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n739), .B2(new_n1101), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(G150), .C2(new_n1014), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n798), .A2(G159), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G33), .B(G41), .C1(new_n751), .C2(G124), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1149), .B1(new_n1145), .B2(new_n1144), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1138), .B1(new_n1160), .B2(new_n713), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1119), .B2(new_n708), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1137), .A2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1136), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(G375));
  NAND3_X1  g0965(.A1(new_n1084), .A2(new_n1081), .A3(new_n1086), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1088), .A2(new_n985), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n702), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1075), .A2(new_n707), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n704), .B1(new_n1094), .B2(G68), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n744), .A2(new_n587), .B1(new_n785), .B2(new_n551), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G97), .B2(new_n740), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n747), .A2(new_n761), .B1(new_n746), .B2(new_n474), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n279), .B(new_n1173), .C1(G303), .C2(new_n751), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n951), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n279), .B1(new_n734), .B2(new_n1099), .C1(new_n264), .C2(new_n746), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1139), .B1(new_n271), .B2(new_n725), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(G159), .C2(new_n740), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT124), .Z(new_n1180));
  NAND2_X1  g0980(.A1(new_n729), .A2(G132), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n795), .B2(new_n747), .C1(new_n744), .C2(new_n1101), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1176), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1170), .B1(new_n1183), .B2(new_n713), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1168), .B1(new_n1169), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1167), .A2(new_n1185), .ZN(G381));
  OR4_X1    g0986(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1187), .A2(G387), .A3(G381), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1091), .A2(new_n1114), .A3(KEYINPUT125), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT125), .B1(new_n1091), .B2(new_n1114), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1164), .A3(new_n1191), .ZN(G407));
  NAND2_X1  g0992(.A1(new_n647), .A2(G213), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1164), .A2(new_n1191), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(G407), .A2(G213), .A3(new_n1195), .ZN(G409));
  NAND3_X1  g0996(.A1(new_n1136), .A2(G378), .A3(new_n1163), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1134), .A2(new_n703), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1162), .B(new_n1198), .C1(new_n1130), .C2(new_n984), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1191), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1193), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1088), .A2(KEYINPUT60), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1203), .A2(new_n1166), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n668), .B1(new_n1203), .B2(new_n1166), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1185), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(G384), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(G384), .B(new_n1185), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1194), .A2(G2897), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT61), .B1(new_n1202), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT63), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1202), .B2(new_n1210), .ZN(new_n1219));
  INV_X1    g1019(.A(G390), .ZN(new_n1220));
  OR2_X1    g1020(.A1(G387), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(G393), .B(G396), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G387), .A2(new_n1220), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1221), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1221), .A2(KEYINPUT126), .A3(new_n1226), .A4(new_n1224), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1194), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1210), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(KEYINPUT63), .A3(new_n1232), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1217), .A2(new_n1219), .A3(new_n1230), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT62), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1231), .A2(new_n1235), .A3(new_n1232), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT61), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n1231), .B2(new_n1215), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1235), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1234), .B1(new_n1240), .B2(new_n1230), .ZN(G405));
  AOI211_X1 g1041(.A(new_n1190), .B(new_n1189), .C1(new_n1136), .C2(new_n1163), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1197), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1242), .A2(new_n1243), .A3(new_n1232), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT127), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1228), .A2(new_n1246), .A3(new_n1229), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1223), .A2(new_n1224), .B1(new_n1226), .B2(new_n1221), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1229), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT127), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1232), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1245), .A2(new_n1247), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1251), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1246), .B(new_n1253), .C1(new_n1254), .C2(new_n1244), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1255), .ZN(G402));
endmodule


