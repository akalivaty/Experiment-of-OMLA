//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n601, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT65), .Z(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n451), .B(new_n452), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(new_n463), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n476));
  INV_X1    g051(.A(G136), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n469), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n463), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n478), .B1(G124), .B2(new_n483), .ZN(G162));
  NAND4_X1  g059(.A1(new_n479), .A2(new_n481), .A3(G126), .A4(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT69), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n461), .A2(new_n487), .A3(G126), .A4(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n479), .A2(new_n481), .A3(G138), .A4(new_n463), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n461), .A2(new_n492), .A3(G138), .A4(new_n463), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n489), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  XOR2_X1   g077(.A(KEYINPUT70), .B(G651), .Z(new_n503));
  OR2_X1    g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(KEYINPUT70), .A2(KEYINPUT71), .A3(G651), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(KEYINPUT6), .C1(KEYINPUT70), .C2(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT71), .A3(G651), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n506), .A2(G88), .A3(new_n501), .A4(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n506), .A2(G50), .A3(G543), .A4(new_n508), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT72), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT72), .B1(new_n509), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n506), .A2(new_n501), .A3(new_n508), .ZN(new_n517));
  INV_X1    g092(.A(G89), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n501), .B(KEYINPUT73), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n506), .A2(G543), .A3(new_n508), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n522), .A2(new_n524), .A3(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  AOI22_X1  g104(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n503), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n532), .A2(new_n525), .B1(new_n517), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT5), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT5), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT73), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n536), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT75), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n546), .B(new_n536), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  INV_X1    g122(.A(new_n503), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n517), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT76), .B(G81), .ZN(new_n551));
  AOI22_X1  g126(.A1(G43), .A2(new_n526), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n526), .A2(G53), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(G651), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n501), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G91), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n563), .A2(new_n564), .B1(new_n517), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n562), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G49), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n570), .A2(new_n525), .B1(new_n517), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n542), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n572), .B1(new_n574), .B2(G651), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G288));
  NAND4_X1  g151(.A1(new_n506), .A2(G48), .A3(G543), .A4(new_n508), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n506), .A2(G86), .A3(new_n501), .A4(new_n508), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n503), .ZN(G305));
  AOI22_X1  g155(.A1(G47), .A2(new_n526), .B1(new_n550), .B2(G85), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n503), .ZN(G290));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NOR2_X1   g159(.A1(G171), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT77), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n541), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n526), .A2(G54), .B1(G651), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OR3_X1    g166(.A1(new_n517), .A2(KEYINPUT10), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT10), .B1(new_n517), .B2(new_n591), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n586), .B1(G868), .B2(new_n595), .ZN(G284));
  OAI21_X1  g171(.A(new_n586), .B1(G868), .B2(new_n595), .ZN(G321));
  NAND2_X1  g172(.A1(G299), .A2(new_n584), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(G168), .B2(new_n584), .ZN(G297));
  OAI21_X1  g174(.A(new_n598), .B1(G168), .B2(new_n584), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n553), .A2(new_n584), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n594), .A2(G559), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT78), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n605), .B2(new_n584), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g182(.A1(new_n482), .A2(G2105), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G135), .ZN(new_n609));
  OAI21_X1  g184(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n463), .A2(G111), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G123), .B2(new_n483), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT79), .Z(new_n614));
  XOR2_X1   g189(.A(KEYINPUT80), .B(G2096), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n461), .A2(new_n467), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(G156));
  XOR2_X1   g196(.A(KEYINPUT81), .B(G2438), .Z(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT15), .B(G2435), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G1341), .B(G1348), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n629), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G14), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(G401));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  XOR2_X1   g212(.A(G2067), .B(G2678), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n637), .B1(new_n641), .B2(KEYINPUT18), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2096), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2100), .Z(new_n644));
  AND2_X1   g219(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n639), .A2(new_n640), .ZN(new_n646));
  AOI21_X1  g221(.A(KEYINPUT18), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(G227));
  XNOR2_X1  g223(.A(G1961), .B(G1966), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT83), .ZN(new_n650));
  XOR2_X1   g225(.A(G1956), .B(G2474), .Z(new_n651));
  AND2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT20), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n650), .A2(new_n651), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(new_n655), .ZN(new_n659));
  OR3_X1    g234(.A1(new_n652), .A2(new_n658), .A3(new_n655), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1991), .B(G1996), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1981), .B(G1986), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G229));
  NAND2_X1  g243(.A1(new_n483), .A2(G119), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n608), .A2(G131), .ZN(new_n670));
  OAI21_X1  g245(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n463), .A2(G107), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n669), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  MUX2_X1   g248(.A(G25), .B(new_n673), .S(G29), .Z(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT35), .B(G1991), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  MUX2_X1   g251(.A(G24), .B(G290), .S(G16), .Z(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT85), .B(G1986), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G22), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G166), .B2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(G1971), .Z(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(G23), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n575), .B2(new_n680), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT86), .B(KEYINPUT33), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(G6), .B(G305), .S(G16), .Z(new_n689));
  XOR2_X1   g264(.A(KEYINPUT32), .B(G1981), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n683), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(KEYINPUT34), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n694), .A2(new_n693), .A3(KEYINPUT34), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n693), .B2(KEYINPUT34), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n676), .B(new_n679), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT88), .B(KEYINPUT36), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n680), .A2(KEYINPUT23), .A3(G20), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT23), .ZN(new_n701));
  INV_X1    g276(.A(G20), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G16), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT9), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n561), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(new_n566), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n700), .B(new_n703), .C1(new_n706), .C2(new_n680), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1956), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(G28), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(G28), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(KEYINPUT24), .A2(G34), .ZN(new_n714));
  NOR2_X1   g289(.A1(KEYINPUT24), .A2(G34), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n714), .A2(new_n715), .A3(G29), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n473), .B2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G2084), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n713), .B1(new_n717), .B2(new_n718), .C1(new_n614), .C2(new_n712), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n712), .A2(G26), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n483), .A2(G128), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n608), .A2(G140), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n463), .A2(G116), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n721), .B(new_n722), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n720), .B1(new_n725), .B2(G29), .ZN(new_n726));
  MUX2_X1   g301(.A(new_n720), .B(new_n726), .S(KEYINPUT28), .Z(new_n727));
  INV_X1    g302(.A(G2067), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n719), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT31), .B(G11), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n595), .A2(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G4), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G1348), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n730), .A2(new_n731), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT27), .B(G1996), .ZN(new_n738));
  AOI22_X1  g313(.A1(G129), .A2(new_n483), .B1(new_n608), .B2(G141), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n467), .A2(G105), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT91), .Z(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(new_n712), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n712), .B2(G32), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n708), .B(new_n737), .C1(new_n738), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G16), .A2(G19), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n554), .B2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT89), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G1341), .Z(new_n752));
  NOR2_X1   g327(.A1(new_n747), .A2(new_n738), .ZN(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G35), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G162), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2090), .ZN(new_n757));
  NOR2_X1   g332(.A1(G27), .A2(G29), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G164), .B2(G29), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G2078), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n759), .A2(G2078), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n753), .A2(new_n757), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n680), .A2(G21), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G168), .B2(new_n680), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G1966), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT92), .B1(G5), .B2(G16), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g343(.A1(KEYINPUT92), .A2(G5), .A3(G16), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n768), .B(new_n769), .C1(G171), .C2(G16), .ZN(new_n770));
  OAI22_X1  g345(.A1(new_n765), .A2(new_n766), .B1(G1961), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n766), .B2(new_n765), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n748), .A2(new_n752), .A3(new_n762), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n699), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n717), .A2(new_n718), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n467), .A2(G103), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT25), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n608), .A2(G139), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n777), .B(new_n778), .C1(new_n463), .C2(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G33), .B(new_n780), .S(G29), .Z(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G2072), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n697), .A2(new_n698), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n774), .A2(new_n775), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n770), .A2(G1961), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT93), .Z(new_n786));
  NOR2_X1   g361(.A1(new_n784), .A2(new_n786), .ZN(G311));
  INV_X1    g362(.A(G311), .ZN(G150));
  AOI22_X1  g363(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(new_n503), .ZN(new_n790));
  INV_X1    g365(.A(G55), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT94), .B(G93), .ZN(new_n792));
  OAI22_X1  g367(.A1(new_n791), .A2(new_n525), .B1(new_n517), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G860), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT97), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT37), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(KEYINPUT95), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n790), .A2(new_n793), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n553), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n554), .A2(new_n800), .A3(new_n799), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT38), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n594), .A2(new_n601), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT96), .ZN(new_n810));
  INV_X1    g385(.A(G860), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n808), .B2(KEYINPUT39), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n797), .B1(new_n810), .B2(new_n812), .ZN(G145));
  MUX2_X1   g388(.A(new_n745), .B(new_n744), .S(new_n780), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(new_n618), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n673), .B(new_n725), .Z(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n483), .A2(G130), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n608), .A2(G142), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n463), .A2(G118), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n499), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n815), .A2(new_n816), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n817), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n823), .B1(new_n817), .B2(new_n824), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n614), .B(new_n473), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(G162), .Z(new_n829));
  NOR3_X1   g404(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT99), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n826), .B2(new_n827), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(KEYINPUT98), .B(new_n829), .C1(new_n826), .C2(new_n827), .ZN(new_n835));
  AOI21_X1  g410(.A(G37), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g413(.A1(new_n794), .A2(new_n584), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n804), .B(new_n605), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n706), .A2(new_n594), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n706), .B2(new_n594), .ZN(new_n845));
  NAND3_X1  g420(.A1(G299), .A2(KEYINPUT100), .A3(new_n595), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n841), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n849), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(KEYINPUT102), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n840), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n851), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(new_n840), .ZN(new_n859));
  XOR2_X1   g434(.A(G290), .B(G305), .Z(new_n860));
  XOR2_X1   g435(.A(new_n575), .B(G303), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT103), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT42), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n859), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n839), .B1(new_n865), .B2(new_n584), .ZN(G295));
  OAI21_X1  g441(.A(new_n839), .B1(new_n865), .B2(new_n584), .ZN(G331));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n868));
  XNOR2_X1  g443(.A(G286), .B(G171), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n869), .A2(new_n803), .A3(new_n802), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n803), .B2(new_n802), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n804), .A2(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT104), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n874), .A3(new_n851), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT105), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n870), .A2(new_n871), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n855), .A2(new_n856), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n862), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n872), .A2(new_n874), .A3(new_n880), .A4(new_n851), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n876), .A2(new_n878), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT107), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n876), .A2(new_n878), .A3(new_n881), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n862), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT106), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n888));
  AOI211_X1 g463(.A(new_n888), .B(G37), .C1(new_n884), .C2(new_n862), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n883), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n887), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n882), .B(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n885), .A2(KEYINPUT106), .A3(new_n886), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n894), .A2(new_n896), .A3(new_n892), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT108), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n872), .A2(new_n874), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n848), .A2(KEYINPUT41), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n858), .B1(new_n903), .B2(new_n877), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n849), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n862), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n896), .A2(new_n886), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n900), .B1(new_n907), .B2(KEYINPUT43), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n893), .A2(new_n899), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n896), .A2(new_n892), .A3(new_n886), .A4(new_n906), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n890), .B2(new_n892), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n900), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(G397));
  AOI21_X1  g488(.A(new_n497), .B1(new_n486), .B2(new_n488), .ZN(new_n914));
  AOI21_X1  g489(.A(G1384), .B1(new_n914), .B2(new_n494), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(KEYINPUT45), .ZN(new_n916));
  INV_X1    g491(.A(G40), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n464), .A2(new_n471), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(G1996), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n920), .A2(KEYINPUT46), .ZN(new_n921));
  INV_X1    g496(.A(new_n919), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n725), .B(new_n728), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n924), .B2(new_n744), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(KEYINPUT46), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT47), .Z(new_n928));
  NOR3_X1   g503(.A1(new_n919), .A2(G1986), .A3(G290), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT126), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT48), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n920), .A2(new_n745), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n932), .A2(KEYINPUT109), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(KEYINPUT109), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n744), .A2(G1996), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n919), .B1(new_n923), .B2(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  XOR2_X1   g512(.A(new_n673), .B(new_n675), .Z(new_n938));
  OAI21_X1  g513(.A(new_n937), .B1(new_n919), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n931), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n673), .A2(new_n675), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n941), .A2(KEYINPUT125), .ZN(new_n944));
  OAI22_X1  g519(.A1(new_n943), .A2(new_n944), .B1(G2067), .B2(new_n725), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n928), .B(new_n940), .C1(new_n922), .C2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT124), .ZN(new_n947));
  XOR2_X1   g522(.A(G290), .B(G1986), .Z(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(new_n919), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n939), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT111), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G303), .A2(G8), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n952), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n465), .A2(G40), .A3(new_n472), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n499), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n962), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n965), .B(G1384), .C1(new_n914), .C2(new_n494), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT110), .B1(new_n916), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G1971), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n964), .A2(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n915), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n918), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(G2090), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n961), .B(G8), .C1(new_n971), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(G305), .A2(G1981), .ZN(new_n978));
  NAND2_X1  g553(.A1(G73), .A2(G543), .ZN(new_n979));
  INV_X1    g554(.A(G61), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n979), .B1(new_n541), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n548), .ZN(new_n982));
  INV_X1    g557(.A(G1981), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n983), .A3(new_n577), .A4(new_n578), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT49), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n915), .B2(new_n918), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n978), .A2(KEYINPUT49), .A3(new_n984), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT112), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n987), .A2(new_n993), .A3(new_n989), .A4(new_n990), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n574), .A2(G651), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n526), .A2(G49), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n550), .A2(G87), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n997), .A2(G1976), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(new_n989), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n989), .A2(new_n1000), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n996), .B1(new_n575), .B2(G1976), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n995), .A2(new_n1002), .A3(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n977), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(new_n989), .B(KEYINPUT113), .Z(new_n1009));
  AOI211_X1 g584(.A(G1976), .B(G288), .C1(new_n992), .C2(new_n994), .ZN(new_n1010));
  INV_X1    g585(.A(new_n984), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT63), .ZN(new_n1015));
  OAI21_X1  g590(.A(G8), .B1(new_n971), .B2(new_n976), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n953), .A2(new_n954), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1007), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n915), .A2(KEYINPUT45), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n464), .A2(new_n917), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n966), .A2(new_n472), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n973), .B1(new_n499), .B2(new_n963), .ZN(new_n1022));
  AOI211_X1 g597(.A(KEYINPUT50), .B(G1384), .C1(new_n914), .C2(new_n494), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n962), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n766), .A2(new_n1021), .B1(new_n1024), .B2(new_n718), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(new_n988), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1018), .A2(G168), .A3(new_n977), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1015), .B1(new_n1027), .B2(KEYINPUT114), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1001), .B(new_n1005), .C1(new_n992), .C2(new_n994), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1029), .A2(new_n1030), .A3(new_n977), .A4(new_n1026), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT114), .B(new_n1015), .C1(new_n1031), .C2(G286), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1014), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n975), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(KEYINPUT117), .A3(new_n918), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1348), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n915), .A2(new_n918), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(G2067), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT118), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT117), .B1(new_n1037), .B2(new_n918), .ZN(new_n1043));
  NOR4_X1   g618(.A1(new_n1022), .A2(new_n1023), .A3(new_n1035), .A4(new_n962), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n734), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1041), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT60), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1042), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1042), .A2(new_n1048), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n594), .B1(new_n1051), .B2(KEYINPUT60), .ZN(new_n1052));
  AOI211_X1 g627(.A(new_n1049), .B(new_n595), .C1(new_n1042), .C2(new_n1048), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n968), .A2(new_n970), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(G1996), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT58), .B(G1341), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n915), .B2(new_n918), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n554), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1059), .B(KEYINPUT59), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT61), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT119), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT115), .B(G1956), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n975), .A2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT56), .B(G2072), .Z(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1055), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n562), .B2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(new_n706), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1062), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1071), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n1073), .A2(new_n1074), .B1(KEYINPUT119), .B2(new_n1061), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1075), .B2(new_n1062), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1054), .A2(new_n1060), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1042), .A2(new_n1048), .A3(new_n595), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1074), .B1(new_n1078), .B2(new_n1071), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1029), .A2(new_n1030), .A3(new_n977), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1055), .B2(G2078), .ZN(new_n1084));
  INV_X1    g659(.A(G1961), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n916), .A2(new_n969), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1083), .A2(G2078), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1087), .A2(new_n472), .A3(new_n1088), .A4(new_n1020), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1090), .A2(G171), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n471), .B(KEYINPUT122), .Z(new_n1093));
  NAND4_X1  g668(.A1(new_n1087), .A2(new_n1093), .A3(new_n1088), .A4(new_n1020), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1084), .A2(new_n1086), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1092), .B1(new_n1095), .B2(G171), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1082), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G286), .A2(G8), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1098), .B2(KEYINPUT120), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1098), .B(new_n1100), .C1(new_n1025), .C2(new_n988), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n520), .A2(new_n521), .B1(G51), .B2(new_n526), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n988), .B1(new_n1102), .B2(new_n524), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT51), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1021), .A2(new_n766), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1037), .A2(new_n718), .A3(new_n918), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(G8), .B(new_n1105), .C1(new_n1108), .C2(G286), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(G8), .A3(G286), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1101), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1101), .A2(new_n1109), .A3(KEYINPUT121), .A4(new_n1110), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1090), .A2(G171), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(G171), .B2(new_n1095), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1092), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1097), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1034), .B1(new_n1081), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1113), .A2(new_n1122), .A3(new_n1114), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1082), .A2(new_n1116), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1115), .A2(KEYINPUT62), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1123), .A2(KEYINPUT123), .A3(new_n1124), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n947), .B(new_n951), .C1(new_n1121), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1028), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1013), .B1(new_n1132), .B2(new_n1032), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1060), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1039), .A2(KEYINPUT118), .A3(new_n1041), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1046), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT60), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n595), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1051), .A2(KEYINPUT60), .A3(new_n594), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1134), .B1(new_n1140), .B2(new_n1050), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1079), .B1(new_n1141), .B2(new_n1076), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1130), .B(new_n1133), .C1(new_n1142), .C2(new_n1119), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT124), .B1(new_n1143), .B2(new_n950), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n946), .B1(new_n1131), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT127), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1147), .B(new_n946), .C1(new_n1131), .C2(new_n1144), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g724(.A(G229), .B1(new_n831), .B2(new_n836), .ZN(new_n1151));
  INV_X1    g725(.A(G319), .ZN(new_n1152));
  NOR2_X1   g726(.A1(new_n1152), .A2(G227), .ZN(new_n1153));
  NAND4_X1  g727(.A1(new_n911), .A2(new_n1151), .A3(new_n635), .A4(new_n1153), .ZN(G225));
  INV_X1    g728(.A(G225), .ZN(G308));
endmodule


