//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT73), .B(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(KEYINPUT22), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n202), .B1(new_n209), .B2(KEYINPUT29), .ZN(new_n210));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT2), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  INV_X1    g017(.A(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n211), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(KEYINPUT75), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT75), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(new_n220), .B2(new_n211), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n217), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT76), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(new_n213), .B2(G141gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n215), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n227), .B(new_n228), .C1(new_n215), .C2(G148gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n211), .B1(new_n220), .B2(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n210), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n209), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G228gat), .ZN(new_n238));
  INV_X1    g037(.A(G233gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n233), .A2(G228gat), .A3(G233gat), .A4(new_n236), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G78gat), .B(G106gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT31), .B(G50gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G22gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(KEYINPUT82), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n249), .B2(new_n245), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n242), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n250), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n240), .A2(new_n241), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G169gat), .ZN(new_n256));
  INV_X1    g055(.A(G176gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n260), .B2(KEYINPUT26), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n258), .A2(KEYINPUT26), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n261), .B2(new_n262), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT27), .B(G183gat), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n270), .A2(KEYINPUT66), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n271), .B1(new_n270), .B2(KEYINPUT66), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n266), .B(new_n267), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n267), .A2(KEYINPUT24), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT64), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(G169gat), .B2(G176gat), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(KEYINPUT23), .B2(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n277), .A2(KEYINPUT23), .ZN(new_n279));
  OR2_X1    g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(KEYINPUT24), .A3(new_n267), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n278), .A2(new_n279), .A3(new_n284), .A4(new_n281), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n283), .A2(new_n259), .B1(new_n285), .B2(KEYINPUT25), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT25), .ZN(new_n287));
  NOR4_X1   g086(.A1(new_n282), .A2(new_n284), .A3(new_n287), .A4(new_n260), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n274), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n289), .B2(new_n234), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n293), .A2(new_n294), .A3(new_n209), .ZN(new_n295));
  INV_X1    g094(.A(new_n209), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n285), .A2(KEYINPUT25), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n260), .B2(new_n282), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n283), .A2(KEYINPUT65), .A3(KEYINPUT25), .A4(new_n259), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n272), .A2(new_n273), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n263), .A2(new_n265), .B1(G183gat), .B2(G190gat), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n298), .A2(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n290), .B1(new_n302), .B2(KEYINPUT29), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n296), .B1(new_n303), .B2(new_n292), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT37), .B1(new_n295), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G8gat), .B(G36gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(G64gat), .B(G92gat), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n306), .B(new_n307), .Z(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n209), .B1(new_n293), .B2(new_n294), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n303), .A2(new_n296), .A3(new_n292), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT37), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n305), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT38), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n310), .A2(new_n311), .A3(new_n308), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT38), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n305), .A2(new_n317), .A3(new_n309), .A4(new_n313), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT79), .ZN(new_n320));
  XOR2_X1   g119(.A(G127gat), .B(G134gat), .Z(new_n321));
  INV_X1    g120(.A(G113gat), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT1), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT69), .B(G113gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G120gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n324), .B1(new_n322), .B2(new_n323), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n326), .A2(new_n328), .B1(new_n329), .B2(new_n321), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n221), .B(KEYINPUT75), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n333), .A2(new_n217), .B1(new_n229), .B2(new_n230), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT77), .B1(new_n334), .B2(new_n202), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n232), .A2(new_n336), .A3(KEYINPUT3), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n332), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n330), .A2(new_n225), .A3(new_n231), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n334), .A2(KEYINPUT4), .A3(new_n330), .ZN(new_n342));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n320), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n330), .B1(new_n334), .B2(new_n202), .ZN(new_n346));
  AOI211_X1 g145(.A(KEYINPUT77), .B(new_n202), .C1(new_n225), .C2(new_n231), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n336), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n343), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n350), .B1(new_n339), .B2(new_n340), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n349), .A2(KEYINPUT79), .A3(new_n342), .A4(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n331), .A2(new_n232), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n339), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n353), .B1(new_n355), .B2(new_n350), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n345), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT0), .ZN(new_n359));
  XNOR2_X1  g158(.A(G57gat), .B(G85gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(new_n339), .B2(new_n340), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n365), .A2(new_n349), .A3(new_n343), .A4(new_n353), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n357), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT81), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n357), .A2(new_n366), .ZN(new_n369));
  INV_X1    g168(.A(new_n361), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n357), .A2(new_n374), .A3(new_n361), .A4(new_n366), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n373), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n372), .A2(new_n373), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n255), .B1(new_n319), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT85), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n350), .B1(new_n338), .B2(new_n364), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n355), .A2(new_n350), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT39), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n382), .B(new_n350), .C1(new_n338), .C2(new_n364), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(KEYINPUT83), .A3(new_n361), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT83), .B1(new_n385), .B2(new_n361), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n379), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT40), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT84), .B1(new_n392), .B2(KEYINPUT85), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n391), .A2(new_n392), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n309), .B1(new_n295), .B2(new_n304), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT30), .A4(new_n308), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n316), .A2(KEYINPUT74), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT74), .B1(new_n316), .B2(new_n398), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n371), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT86), .B1(new_n394), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n395), .A2(new_n396), .ZN(new_n405));
  INV_X1    g204(.A(new_n401), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(new_n399), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n361), .B1(new_n357), .B2(new_n366), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n389), .A2(new_n393), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n385), .A2(new_n361), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n414), .A2(new_n386), .B1(new_n380), .B2(new_n383), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT85), .B1(new_n415), .B2(KEYINPUT84), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n411), .B1(new_n416), .B2(KEYINPUT40), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n409), .A2(new_n410), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n378), .B1(new_n404), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n376), .A2(new_n371), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n408), .B1(KEYINPUT81), .B2(new_n367), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n420), .B1(new_n421), .B2(KEYINPUT6), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n254), .B1(new_n422), .B2(new_n402), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT72), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT34), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n289), .A2(new_n330), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n274), .B(new_n331), .C1(new_n286), .C2(new_n288), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G227gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(new_n239), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n425), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  AOI211_X1 g231(.A(KEYINPUT34), .B(new_n430), .C1(new_n426), .C2(new_n427), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n426), .A2(new_n430), .A3(new_n427), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(KEYINPUT70), .A3(new_n436), .ZN(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G43gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n435), .B2(KEYINPUT32), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n435), .B(KEYINPUT32), .C1(new_n436), .C2(new_n443), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n424), .B(new_n434), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n440), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT70), .B1(new_n435), .B2(new_n436), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n434), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT72), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n434), .B(new_n446), .C1(new_n448), .C2(new_n449), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT71), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n445), .A2(KEYINPUT71), .A3(new_n434), .A4(new_n446), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT36), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n450), .A2(new_n451), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n460), .A2(KEYINPUT36), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n458), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n423), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n419), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n434), .B1(new_n445), .B2(new_n446), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(new_n254), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n458), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n377), .A2(new_n407), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n458), .A2(KEYINPUT88), .A3(new_n467), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n460), .A2(new_n424), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n466), .A2(KEYINPUT72), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n458), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT35), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n251), .A2(new_n478), .A3(new_n253), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n422), .A2(new_n402), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(KEYINPUT87), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n458), .A2(new_n475), .A3(new_n476), .ZN(new_n483));
  INV_X1    g282(.A(new_n479), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n377), .A2(new_n407), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(KEYINPUT35), .A2(new_n474), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n465), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G29gat), .ZN(new_n489));
  INV_X1    g288(.A(G36gat), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT89), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(G29gat), .A3(G36gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n494), .B(KEYINPUT91), .Z(new_n495));
  XNOR2_X1  g294(.A(G43gat), .B(G50gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n490), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n500), .A2(KEYINPUT90), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(KEYINPUT90), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n495), .A2(new_n497), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n500), .A2(new_n498), .ZN(new_n506));
  OAI211_X1 g305(.A(KEYINPUT15), .B(new_n496), .C1(new_n506), .C2(new_n494), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT17), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(G1gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(KEYINPUT16), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(new_n512), .B2(new_n511), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT92), .B(G8gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(KEYINPUT93), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(new_n514), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT93), .B1(new_n514), .B2(new_n515), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n505), .A2(KEYINPUT17), .A3(new_n507), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n510), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n508), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT18), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n522), .A2(KEYINPUT18), .A3(new_n523), .A4(new_n525), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n523), .B(KEYINPUT13), .Z(new_n530));
  NOR2_X1   g329(.A1(new_n524), .A2(new_n508), .ZN(new_n531));
  INV_X1    g330(.A(new_n508), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(new_n520), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n530), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G113gat), .B(G141gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(G197gat), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT11), .B(G169gat), .Z(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT12), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n540), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n528), .A2(new_n542), .A3(new_n529), .A4(new_n534), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G85gat), .ZN(new_n550));
  INV_X1    g349(.A(G92gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n546), .A2(new_n549), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n554), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n556), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(KEYINPUT96), .A3(new_n545), .ZN(new_n562));
  AND3_X1   g361(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n559), .B1(new_n555), .B2(new_n556), .ZN(new_n566));
  AOI22_X1  g365(.A1(KEYINPUT8), .A2(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n562), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n510), .A2(new_n521), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n532), .B2(new_n570), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  OAI22_X1  g376(.A1(new_n571), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n578), .B(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT95), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n576), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  XOR2_X1   g384(.A(new_n581), .B(new_n585), .Z(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  AND2_X1   g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G57gat), .B(G64gat), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G57gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(G64gat), .ZN(new_n595));
  INV_X1    g394(.A(G64gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(G57gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G71gat), .B(G78gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n592), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n593), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n520), .B1(new_n587), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n587), .ZN(new_n604));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n603), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT94), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G183gat), .B(G211gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n602), .A2(new_n560), .A3(new_n568), .ZN(new_n617));
  XOR2_X1   g416(.A(KEYINPUT99), .B(KEYINPUT10), .Z(new_n618));
  AOI21_X1  g417(.A(KEYINPUT98), .B1(new_n565), .B2(new_n567), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n593), .B(new_n601), .C1(new_n619), .C2(new_n557), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n554), .A2(new_n621), .A3(new_n557), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n617), .B(new_n618), .C1(new_n620), .C2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n569), .A2(KEYINPUT10), .A3(new_n593), .A4(new_n601), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n617), .B1(new_n620), .B2(new_n622), .ZN(new_n628));
  INV_X1    g427(.A(new_n626), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n586), .A2(new_n616), .A3(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n488), .A2(new_n544), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n422), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n402), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT42), .B1(new_n646), .B2(KEYINPUT100), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT16), .B(G8gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR4_X1   g449(.A1(new_n645), .A2(KEYINPUT100), .A3(KEYINPUT42), .A4(new_n648), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n645), .A2(new_n652), .A3(G8gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n645), .B2(G8gat), .ZN(new_n655));
  OAI22_X1  g454(.A1(new_n650), .A2(new_n651), .B1(new_n654), .B2(new_n655), .ZN(G1325gat));
  NOR2_X1   g455(.A1(new_n488), .A2(new_n544), .ZN(new_n657));
  INV_X1    g456(.A(new_n641), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n462), .B1(new_n477), .B2(KEYINPUT36), .ZN(new_n660));
  OAI21_X1  g459(.A(G15gat), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n483), .A2(G15gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n659), .B2(new_n662), .ZN(G1326gat));
  OAI21_X1  g462(.A(KEYINPUT102), .B1(new_n659), .B2(new_n255), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n642), .A2(new_n665), .A3(new_n254), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(G1327gat));
  NAND2_X1  g468(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n481), .A2(new_n486), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n419), .B2(new_n464), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n541), .A2(new_n543), .ZN(new_n674));
  INV_X1    g473(.A(new_n616), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n640), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n586), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n422), .A2(new_n489), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT45), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n586), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n465), .B2(new_n487), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n676), .A2(new_n544), .ZN(new_n686));
  INV_X1    g485(.A(new_n378), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n394), .A2(new_n403), .A3(KEYINPUT86), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n410), .B1(new_n409), .B2(new_n417), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n423), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n471), .A2(KEYINPUT103), .A3(new_n254), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n690), .A2(new_n694), .A3(new_n660), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n586), .B1(new_n695), .B2(new_n672), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n685), .B(new_n686), .C1(new_n696), .C2(KEYINPUT44), .ZN(new_n697));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697), .B2(new_n377), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n682), .A2(KEYINPUT104), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1328gat));
  NOR3_X1   g502(.A1(new_n678), .A2(G36gat), .A3(new_n407), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n697), .B2(new_n407), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1329gat));
  XNOR2_X1  g506(.A(new_n581), .B(new_n585), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n692), .B(new_n693), .C1(new_n459), .C2(new_n463), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n419), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n710), .B2(new_n487), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n683), .ZN(new_n712));
  INV_X1    g511(.A(new_n660), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n685), .A4(new_n686), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G43gat), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n483), .A2(G43gat), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n678), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n657), .A2(KEYINPUT105), .A3(new_n677), .A4(new_n717), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n715), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT47), .B1(new_n678), .B2(new_n718), .ZN(new_n724));
  INV_X1    g523(.A(G43gat), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n714), .B2(new_n726), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n711), .A2(new_n683), .B1(new_n673), .B2(new_n684), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n728), .A2(KEYINPUT106), .A3(new_n713), .A4(new_n686), .ZN(new_n729));
  AOI211_X1 g528(.A(KEYINPUT107), .B(new_n724), .C1(new_n727), .C2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n726), .B1(new_n697), .B2(new_n660), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(new_n729), .A3(G43gat), .ZN(new_n733));
  INV_X1    g532(.A(new_n724), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n723), .B1(new_n730), .B2(new_n735), .ZN(G1330gat));
  NOR2_X1   g535(.A1(new_n678), .A2(new_n255), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n254), .A2(G50gat), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n737), .A2(G50gat), .B1(new_n697), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1331gat));
  NAND2_X1  g540(.A1(new_n695), .A2(new_n672), .ZN(new_n742));
  NOR4_X1   g541(.A1(new_n708), .A2(new_n674), .A3(new_n675), .A4(new_n640), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n377), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(new_n594), .ZN(G1332gat));
  NOR2_X1   g545(.A1(new_n744), .A2(new_n407), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  INV_X1    g550(.A(G71gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n744), .B2(new_n483), .ZN(new_n753));
  INV_X1    g552(.A(new_n744), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n660), .A2(new_n752), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n754), .A2(KEYINPUT109), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT109), .B1(new_n754), .B2(new_n755), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g558(.A1(new_n754), .A2(new_n254), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g560(.A1(new_n674), .A2(new_n616), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n728), .A2(new_n639), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G85gat), .B1(new_n763), .B2(new_n377), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n696), .A2(new_n762), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n766), .A2(KEYINPUT110), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(KEYINPUT110), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n696), .A2(KEYINPUT110), .A3(new_n766), .A4(new_n762), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n377), .A2(G85gat), .A3(new_n640), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n764), .A2(new_n772), .ZN(G1336gat));
  NAND4_X1  g572(.A1(new_n728), .A2(new_n402), .A3(new_n639), .A4(new_n762), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n407), .A2(G92gat), .A3(new_n640), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n769), .A2(new_n770), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n765), .A2(KEYINPUT111), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT51), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n781), .A2(new_n777), .B1(G92gat), .B2(new_n774), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n782), .B2(new_n776), .ZN(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n763), .B2(new_n660), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n483), .A2(G99gat), .A3(new_n640), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n784), .A2(KEYINPUT112), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(G1338gat));
  NAND4_X1  g590(.A1(new_n728), .A2(new_n254), .A3(new_n639), .A4(new_n762), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G106gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n255), .A2(G106gat), .A3(new_n640), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n769), .A2(new_n770), .A3(new_n794), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AOI22_X1  g596(.A1(new_n781), .A2(new_n794), .B1(G106gat), .B2(new_n792), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(G1339gat));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n641), .A2(new_n674), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n625), .B2(new_n626), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n623), .A2(new_n629), .A3(new_n624), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT114), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n808), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n625), .A2(new_n803), .A3(new_n626), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n635), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n810), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  AND4_X1   g614(.A1(new_n808), .A2(new_n627), .A3(KEYINPUT54), .A4(new_n805), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n808), .B1(new_n804), .B2(new_n805), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT115), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n812), .A2(new_n635), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n816), .B2(new_n817), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT116), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n822), .A2(new_n826), .A3(new_n823), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n820), .A2(new_n825), .A3(new_n637), .A4(new_n827), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n531), .A2(new_n533), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n523), .B1(new_n522), .B2(new_n525), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n829), .A2(new_n530), .B1(new_n830), .B2(KEYINPUT117), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n830), .A2(KEYINPUT117), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n539), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n543), .ZN(new_n834));
  OR3_X1    g633(.A1(new_n586), .A2(new_n828), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n543), .A3(new_n639), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n828), .B2(new_n544), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n586), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n802), .B1(new_n839), .B2(new_n675), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n801), .B1(new_n840), .B2(new_n254), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n586), .A2(new_n828), .A3(new_n834), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n586), .A2(new_n837), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n675), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n802), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(KEYINPUT118), .A3(new_n255), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n483), .A2(new_n377), .A3(new_n402), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n544), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n840), .A2(new_n377), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n470), .A2(new_n473), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n402), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n544), .A2(new_n327), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n851), .B1(new_n855), .B2(new_n856), .ZN(G1340gat));
  INV_X1    g656(.A(new_n855), .ZN(new_n858));
  AOI21_X1  g657(.A(G120gat), .B1(new_n858), .B2(new_n639), .ZN(new_n859));
  INV_X1    g658(.A(new_n850), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n640), .A2(new_n323), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(G1341gat));
  OAI21_X1  g661(.A(G127gat), .B1(new_n850), .B2(new_n675), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n675), .A2(G127gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n855), .B2(new_n864), .ZN(G1342gat));
  NOR3_X1   g664(.A1(new_n855), .A2(G134gat), .A3(new_n586), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT56), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n850), .B2(new_n586), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n377), .A2(new_n402), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n660), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n872), .B1(new_n840), .B2(new_n255), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n636), .B1(new_n822), .B2(new_n823), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n811), .B1(new_n810), .B2(new_n814), .ZN(new_n876));
  AOI211_X1 g675(.A(KEYINPUT115), .B(new_n813), .C1(new_n807), .C2(new_n809), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n674), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n875), .B1(new_n820), .B2(new_n874), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n836), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n708), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n836), .B(KEYINPUT120), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n842), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n845), .B1(new_n885), .B2(new_n616), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n255), .A2(new_n872), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n871), .B1(new_n873), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(G141gat), .A3(new_n674), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n713), .A2(new_n402), .A3(new_n255), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n852), .A2(new_n674), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n215), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n890), .B(new_n893), .C1(KEYINPUT121), .C2(KEYINPUT58), .ZN(new_n894));
  NAND2_X1  g693(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n894), .B(new_n895), .ZN(G1344gat));
  NAND2_X1  g695(.A1(new_n852), .A2(new_n891), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n213), .A3(new_n639), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n889), .A2(new_n639), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n213), .A2(KEYINPUT59), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n902), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT122), .B(new_n904), .C1(new_n889), .C2(new_n639), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  INV_X1    g706(.A(new_n887), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n844), .B2(new_n845), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n881), .A2(new_n882), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n586), .A3(new_n884), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n616), .B1(new_n911), .B2(new_n835), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n254), .B1(new_n912), .B2(new_n802), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n909), .B1(new_n913), .B2(new_n872), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n660), .A2(new_n639), .A3(new_n870), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n914), .A2(KEYINPUT123), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(new_n213), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT123), .B1(new_n914), .B2(new_n915), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n907), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n899), .B1(new_n906), .B2(new_n919), .ZN(G1345gat));
  INV_X1    g719(.A(new_n889), .ZN(new_n921));
  OAI21_X1  g720(.A(G155gat), .B1(new_n921), .B2(new_n675), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n898), .A2(new_n218), .A3(new_n616), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  NAND3_X1  g723(.A1(new_n898), .A2(new_n219), .A3(new_n708), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT124), .ZN(new_n926));
  OAI21_X1  g725(.A(G162gat), .B1(new_n921), .B2(new_n586), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n840), .A2(new_n422), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n853), .A2(new_n407), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n674), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n422), .A2(new_n407), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n477), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT125), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n848), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n544), .A2(new_n256), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(G1348gat));
  AOI21_X1  g738(.A(new_n257), .B1(new_n937), .B2(new_n639), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n931), .A2(G176gat), .A3(new_n640), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n940), .A2(new_n941), .ZN(G1349gat));
  NAND3_X1  g741(.A1(new_n848), .A2(new_n616), .A3(new_n936), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(G183gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n932), .A2(new_n268), .A3(new_n616), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n269), .A3(new_n708), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n937), .A2(new_n708), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(G190gat), .ZN(new_n951));
  AOI211_X1 g750(.A(KEYINPUT61), .B(new_n269), .C1(new_n937), .C2(new_n708), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(G1351gat));
  NOR3_X1   g752(.A1(new_n713), .A2(new_n407), .A3(new_n255), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n929), .A2(new_n954), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n955), .A2(G197gat), .A3(new_n544), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n660), .A2(new_n934), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n914), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT126), .B1(new_n959), .B2(new_n544), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G197gat), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n959), .A2(KEYINPUT126), .A3(new_n544), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n956), .B1(new_n961), .B2(new_n962), .ZN(G1352gat));
  NOR3_X1   g762(.A1(new_n955), .A2(G204gat), .A3(new_n640), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT62), .ZN(new_n965));
  OAI21_X1  g764(.A(G204gat), .B1(new_n959), .B2(new_n640), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1353gat));
  NAND4_X1  g766(.A1(new_n929), .A2(new_n205), .A3(new_n616), .A4(new_n954), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n914), .A2(new_n675), .A3(new_n957), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n205), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n957), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT57), .B1(new_n886), .B2(new_n254), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n616), .B(new_n972), .C1(new_n973), .C2(new_n909), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT127), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n913), .A2(new_n872), .ZN(new_n977));
  INV_X1    g776(.A(new_n909), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n979), .A2(new_n970), .A3(new_n616), .A4(new_n972), .ZN(new_n980));
  AND4_X1   g779(.A1(KEYINPUT63), .A2(new_n975), .A3(new_n980), .A4(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n968), .B1(new_n976), .B2(new_n981), .ZN(G1354gat));
  NOR2_X1   g781(.A1(new_n586), .A2(new_n204), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n929), .A2(new_n708), .A3(new_n954), .ZN(new_n984));
  INV_X1    g783(.A(G218gat), .ZN(new_n985));
  AOI22_X1  g784(.A1(new_n958), .A2(new_n983), .B1(new_n984), .B2(new_n985), .ZN(G1355gat));
endmodule


