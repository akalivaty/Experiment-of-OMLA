//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(KEYINPUT67), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(KEYINPUT67), .ZN(new_n463));
  OAI21_X1  g038(.A(G101), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT66), .B1(new_n468), .B2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n460), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n460), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n474), .A2(new_n478), .ZN(G160));
  NAND4_X1  g054(.A1(new_n471), .A2(new_n467), .A3(G2105), .A4(new_n469), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n460), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n472), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G136), .ZN(G162));
  INV_X1    g061(.A(new_n480), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n460), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT68), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n488), .B2(new_n489), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n487), .A2(G126), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n471), .A2(new_n467), .A3(new_n469), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n475), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(KEYINPUT69), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(new_n493), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n488), .A2(new_n489), .A3(new_n492), .ZN(new_n505));
  INV_X1    g080(.A(G126), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n504), .A2(new_n505), .B1(new_n480), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n475), .B2(new_n499), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT73), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT70), .B(G651), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT72), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT70), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G651), .ZN(new_n529));
  AND4_X1   g104(.A1(new_n524), .A2(new_n527), .A3(new_n529), .A4(KEYINPUT6), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n523), .B(new_n517), .C1(new_n525), .C2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G88), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n527), .A2(new_n529), .A3(KEYINPUT6), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT71), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n527), .A2(new_n529), .A3(new_n524), .A4(KEYINPUT6), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G543), .A3(new_n523), .ZN(new_n537));
  INV_X1    g112(.A(G50), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n520), .B1(new_n531), .B2(new_n532), .C1(new_n537), .C2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  NAND2_X1  g115(.A1(new_n522), .A2(KEYINPUT72), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n522), .A2(KEYINPUT72), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n534), .A2(new_n535), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT74), .B(G89), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n543), .A2(new_n517), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n536), .A2(G51), .A3(G543), .A4(new_n523), .ZN(new_n546));
  AND2_X1   g121(.A1(G63), .A2(G651), .ZN(new_n547));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n517), .A2(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n545), .A2(new_n546), .A3(new_n551), .ZN(G168));
  XNOR2_X1  g127(.A(KEYINPUT75), .B(G52), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n536), .A2(G543), .A3(new_n523), .A4(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n536), .A2(G90), .A3(new_n523), .A4(new_n517), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n517), .A2(G64), .ZN(new_n556));
  NAND2_X1  g131(.A1(G77), .A2(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n519), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n554), .A2(new_n555), .A3(new_n560), .ZN(G171));
  NAND3_X1  g136(.A1(new_n543), .A2(G81), .A3(new_n517), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n543), .A2(G43), .A3(G543), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n519), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n537), .A2(new_n572), .B1(KEYINPUT76), .B2(KEYINPUT9), .ZN(new_n573));
  XNOR2_X1  g148(.A(KEYINPUT76), .B(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n543), .A2(G53), .A3(G543), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n531), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n517), .A2(G65), .ZN(new_n578));
  INV_X1    g153(.A(G78), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT77), .B1(new_n579), .B2(new_n512), .ZN(new_n580));
  OR3_X1    g155(.A1(new_n579), .A2(new_n512), .A3(KEYINPUT77), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n577), .A2(G91), .B1(G651), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n576), .A2(new_n583), .ZN(G299));
  NAND3_X1  g159(.A1(new_n554), .A2(new_n555), .A3(new_n560), .ZN(G301));
  NAND3_X1  g160(.A1(new_n545), .A2(new_n546), .A3(new_n551), .ZN(G286));
  NAND2_X1  g161(.A1(new_n577), .A2(G87), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n543), .A2(G49), .A3(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  NAND3_X1  g165(.A1(new_n543), .A2(G48), .A3(G543), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n519), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n591), .B(new_n593), .C1(new_n594), .C2(new_n531), .ZN(G305));
  NAND2_X1  g170(.A1(new_n577), .A2(G85), .ZN(new_n596));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI221_X1 g173(.A(new_n596), .B1(new_n597), .B2(new_n537), .C1(new_n519), .C2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n543), .A2(G54), .A3(G543), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n517), .A2(G66), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT79), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT78), .B1(new_n531), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n543), .A2(new_n609), .A3(G92), .A4(new_n517), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n608), .A2(new_n613), .A3(new_n610), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n606), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n600), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n600), .B1(new_n615), .B2(G868), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  XOR2_X1   g195(.A(G280), .B(KEYINPUT80), .Z(G297));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI22_X1  g200(.A1(new_n625), .A2(KEYINPUT81), .B1(G868), .B2(new_n566), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(KEYINPUT81), .B2(new_n625), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT82), .Z(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g204(.A(new_n461), .B(KEYINPUT67), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(new_n475), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n487), .A2(G123), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n637), .C1(new_n638), .C2(new_n472), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n634), .A2(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  XOR2_X1   g219(.A(new_n643), .B(new_n644), .Z(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT85), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT84), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT83), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n649), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n649), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT86), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(G2072), .A2(G2078), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n663), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n663), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n671), .A2(new_n664), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n667), .B(KEYINPUT88), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n663), .A2(new_n665), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n667), .B(KEYINPUT17), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  OAI221_X1 g252(.A(new_n670), .B1(new_n673), .B2(new_n674), .C1(new_n675), .C2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  MUX2_X1   g272(.A(G24), .B(G290), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT89), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(G1986), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G25), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n485), .A2(G131), .ZN(new_n703));
  INV_X1    g278(.A(G119), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n460), .A2(G107), .ZN(new_n705));
  OAI21_X1  g280(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n706));
  OAI22_X1  g281(.A1(new_n480), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n702), .B1(new_n709), .B2(new_n701), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n700), .A2(KEYINPUT90), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(G23), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n714), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G6), .B(G305), .S(G16), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT32), .B(G1981), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n718), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n699), .A2(G1986), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n713), .A2(new_n728), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  NOR2_X1   g309(.A1(G29), .A2(G32), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT26), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n630), .A2(G105), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n487), .A2(G129), .ZN(new_n741));
  INV_X1    g316(.A(G141), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n740), .B(new_n741), .C1(new_n742), .C2(new_n472), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT92), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT93), .Z(new_n745));
  AOI21_X1  g320(.A(new_n735), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT27), .B(G1996), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n566), .A2(G16), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G16), .B2(G19), .ZN(new_n750));
  INV_X1    g325(.A(G1341), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NOR2_X1   g328(.A1(G5), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G171), .B2(G16), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT97), .B(G1961), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n752), .B(new_n753), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n714), .A2(G20), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT23), .Z(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G299), .B2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  NAND2_X1  g336(.A1(G168), .A2(G16), .ZN(new_n762));
  NOR2_X1   g337(.A1(G16), .A2(G21), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(KEYINPUT94), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT94), .B2(new_n762), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1966), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n757), .A2(new_n761), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G29), .A2(G33), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT91), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n485), .A2(G139), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(new_n460), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT25), .Z(new_n774));
  NAND3_X1  g349(.A1(new_n770), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n769), .B1(new_n775), .B2(new_n701), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2072), .ZN(new_n777));
  AND2_X1   g352(.A1(KEYINPUT24), .A2(G34), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n701), .B1(KEYINPUT24), .B2(G34), .ZN(new_n779));
  OAI22_X1  g354(.A1(G160), .A2(new_n701), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G29), .A2(G35), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G162), .B2(G29), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT29), .B(G2090), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n777), .B1(G2084), .B2(new_n780), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n755), .A2(new_n756), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n701), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n701), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G2078), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n701), .A2(G26), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  INV_X1    g366(.A(G128), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n460), .A2(G116), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n480), .A2(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n485), .B2(G140), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n791), .B1(new_n796), .B2(new_n701), .ZN(new_n797));
  INV_X1    g372(.A(G2067), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT31), .B(G11), .Z(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT96), .B(G28), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT30), .ZN(new_n802));
  AOI21_X1  g377(.A(G29), .B1(new_n801), .B2(KEYINPUT30), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n639), .A2(new_n701), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n800), .B(new_n804), .C1(new_n805), .C2(KEYINPUT95), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(KEYINPUT95), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n780), .A2(G2084), .B1(new_n782), .B2(new_n783), .ZN(new_n808));
  AND4_X1   g383(.A1(new_n799), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n786), .A2(new_n789), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n714), .A2(G4), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n615), .B2(new_n714), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1348), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n748), .A2(new_n767), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n733), .A2(new_n734), .A3(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  NAND2_X1  g391(.A1(new_n615), .A2(G559), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT38), .Z(new_n818));
  NAND3_X1  g393(.A1(new_n543), .A2(G93), .A3(new_n517), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n543), .A2(G55), .A3(G543), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(new_n519), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n566), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n818), .B(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT98), .B(G860), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n823), .A2(new_n832), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT37), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(G145));
  INV_X1    g411(.A(new_n775), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n745), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n744), .A2(new_n775), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n494), .A2(new_n501), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n796), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n709), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n487), .A2(G130), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n460), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  INV_X1    g421(.A(G142), .ZN(new_n847));
  OAI221_X1 g422(.A(new_n844), .B1(new_n845), .B2(new_n846), .C1(new_n847), .C2(new_n472), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n632), .B(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n842), .B(new_n708), .ZN(new_n851));
  INV_X1    g426(.A(new_n849), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n840), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n850), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n855), .A2(new_n838), .A3(new_n839), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n639), .B(KEYINPUT99), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G160), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(G162), .Z(new_n860));
  AOI21_X1  g435(.A(G37), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n860), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n854), .A2(new_n856), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT100), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n861), .A2(new_n866), .A3(new_n863), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n865), .A2(KEYINPUT40), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT40), .B1(new_n865), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(G395));
  XNOR2_X1  g445(.A(new_n624), .B(new_n828), .ZN(new_n871));
  INV_X1    g446(.A(new_n606), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n608), .A2(new_n613), .A3(new_n610), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n613), .B1(new_n608), .B2(new_n610), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n619), .ZN(new_n876));
  OAI211_X1 g451(.A(G299), .B(new_n872), .C1(new_n874), .C2(new_n873), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n615), .B2(G299), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n875), .A2(new_n619), .A3(KEYINPUT101), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n615), .B2(G299), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n883), .A2(new_n884), .B1(new_n876), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n879), .B1(new_n886), .B2(new_n871), .ZN(new_n887));
  XOR2_X1   g462(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n888));
  OR2_X1    g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(G290), .B(G305), .ZN(new_n890));
  XNOR2_X1  g465(.A(G288), .B(G303), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n888), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n889), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n889), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(G868), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(G868), .B2(new_n823), .ZN(G295));
  OAI21_X1  g473(.A(new_n897), .B1(G868), .B2(new_n823), .ZN(G331));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  NAND2_X1  g477(.A1(G301), .A2(KEYINPUT103), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n554), .A2(new_n555), .A3(new_n904), .A4(new_n560), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(G286), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(G168), .A2(G171), .A3(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n828), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n906), .A2(new_n907), .A3(new_n824), .A4(new_n827), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(KEYINPUT104), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n828), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n907), .A4(new_n906), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n878), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n892), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n909), .A2(new_n910), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n883), .A2(new_n884), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n885), .A2(new_n876), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n902), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n915), .A2(new_n878), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n893), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n901), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n881), .A2(new_n885), .A3(new_n882), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n878), .A2(new_n884), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n914), .A3(new_n911), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n918), .A2(new_n878), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n892), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n922), .A2(new_n932), .A3(KEYINPUT43), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n900), .B1(new_n926), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n916), .B(new_n892), .C1(new_n886), .C2(new_n918), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n925), .A2(new_n901), .A3(new_n902), .A4(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(KEYINPUT44), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n922), .B2(new_n932), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n915), .B1(new_n928), .B2(new_n927), .ZN(new_n940));
  INV_X1    g515(.A(new_n931), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n893), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n942), .A2(KEYINPUT105), .A3(new_n902), .A4(new_n935), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(KEYINPUT43), .A3(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n937), .A2(new_n944), .A3(KEYINPUT106), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT106), .B1(new_n937), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n934), .B1(new_n945), .B2(new_n946), .ZN(G397));
  XNOR2_X1  g522(.A(KEYINPUT107), .B(G1384), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n841), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n485), .A2(G137), .ZN(new_n952));
  INV_X1    g527(.A(new_n478), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n952), .A2(new_n953), .A3(G40), .A4(new_n464), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(G290), .A2(G1986), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT109), .Z(new_n957));
  NAND2_X1  g532(.A1(G290), .A2(G1986), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n958), .B(KEYINPUT110), .Z(new_n959));
  OR2_X1    g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n745), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n796), .B(new_n798), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n744), .B2(G1996), .ZN(new_n964));
  OR2_X1    g539(.A1(new_n709), .A2(new_n711), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n709), .A2(new_n711), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n962), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n955), .B1(new_n960), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n720), .A2(G1976), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  INV_X1    g545(.A(G40), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n474), .A2(new_n971), .A3(new_n478), .ZN(new_n972));
  AOI21_X1  g547(.A(G1384), .B1(new_n494), .B2(new_n501), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT52), .ZN(new_n976));
  INV_X1    g551(.A(G1976), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT52), .B1(G288), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n969), .A2(new_n978), .A3(new_n974), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n974), .ZN(new_n981));
  NAND2_X1  g556(.A1(G305), .A2(G1981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n577), .A2(G86), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n591), .A4(new_n593), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n981), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n982), .A2(KEYINPUT49), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT111), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n992), .A3(new_n989), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n980), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(G303), .A2(G8), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n995), .B(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n510), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n972), .B1(new_n973), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G2090), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT45), .B(new_n948), .C1(new_n507), .C2(new_n508), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n972), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n502), .B2(new_n509), .ZN(new_n1008));
  INV_X1    g583(.A(new_n950), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1004), .A2(new_n1005), .B1(new_n717), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n998), .B1(new_n1011), .B2(new_n970), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1002), .B(new_n999), .C1(new_n507), .C2(new_n508), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n972), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1014), .B(new_n1005), .C1(new_n1008), .C2(new_n1002), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n972), .A2(new_n1006), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n1000), .B2(new_n950), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1017), .B2(G1971), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(G8), .A3(new_n997), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n994), .A2(new_n1012), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G2084), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1014), .B(new_n1021), .C1(new_n1008), .C2(new_n1002), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1024));
  INV_X1    g599(.A(new_n973), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n954), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1966), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G286), .A2(G8), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT124), .B(KEYINPUT51), .Z(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1022), .B1(new_n1034), .B2(G1966), .ZN(new_n1035));
  OAI211_X1 g610(.A(G8), .B(new_n1033), .C1(new_n1035), .C2(G286), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(G8), .A3(G286), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1032), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1020), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1008), .A2(new_n1002), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n972), .A2(new_n1013), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT118), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1961), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1014), .B(new_n1044), .C1(new_n1008), .C2(new_n1002), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n1010), .B2(G2078), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(G2078), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n953), .A2(G40), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(KEYINPUT125), .B2(new_n474), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n474), .A2(KEYINPUT125), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n951), .A2(new_n1051), .A3(new_n1006), .A4(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1046), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G171), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1024), .A2(new_n1027), .A3(new_n1049), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1046), .A2(new_n1056), .A3(new_n1048), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1055), .B(KEYINPUT54), .C1(G171), .C2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(G171), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1046), .A2(G301), .A3(new_n1048), .A4(new_n1053), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT54), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT126), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g638(.A(KEYINPUT126), .B(KEYINPUT54), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1039), .B(new_n1058), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT120), .B(G1996), .Z(new_n1066));
  NAND2_X1  g641(.A1(new_n1017), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n972), .A2(new_n973), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT58), .B(G1341), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n825), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT59), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1007), .B(new_n1073), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1017), .A2(KEYINPUT116), .A3(new_n1073), .ZN(new_n1077));
  INV_X1    g652(.A(G1956), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n576), .B2(KEYINPUT115), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G299), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n576), .B(new_n583), .C1(KEYINPUT115), .C2(KEYINPUT57), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1084), .A2(new_n1076), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1087), .A2(KEYINPUT117), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(KEYINPUT117), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1072), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1348), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1042), .A2(new_n1093), .A3(new_n1045), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n972), .A2(new_n798), .A3(new_n973), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT60), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(KEYINPUT123), .A3(new_n615), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1096), .B2(new_n875), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1086), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1087), .B1(new_n1107), .B2(KEYINPUT122), .ZN(new_n1108));
  OR3_X1    g683(.A1(new_n1080), .A2(new_n1085), .A3(KEYINPUT122), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(KEYINPUT61), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1098), .A2(new_n1104), .A3(new_n1100), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1092), .A2(new_n1106), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1087), .B(KEYINPUT117), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1102), .A2(new_n615), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1086), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1113), .A2(KEYINPUT119), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT119), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1065), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n1120));
  OAI211_X1 g695(.A(G8), .B(G168), .C1(new_n1023), .C2(new_n1028), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT113), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT113), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1035), .A2(new_n1123), .A3(G8), .A4(G168), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(new_n994), .A3(new_n1012), .A4(new_n1019), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT114), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n976), .A2(new_n979), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n988), .A2(new_n992), .A3(new_n989), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n992), .B1(new_n988), .B2(new_n989), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1129), .B(new_n1019), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1133));
  OAI22_X1  g708(.A1(new_n1133), .A2(G2090), .B1(G1971), .B2(new_n1017), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n997), .B1(new_n1134), .B2(G8), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT114), .B1(new_n1136), .B2(new_n1125), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1125), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1018), .A2(G8), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1120), .B1(new_n1139), .B2(new_n998), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n994), .A2(new_n1019), .A3(new_n1140), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n1128), .A2(new_n1137), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1032), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT62), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1059), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1032), .A2(new_n1036), .A3(new_n1146), .A4(new_n1037), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1144), .A2(new_n1136), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n977), .B(new_n720), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n985), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n974), .B(KEYINPUT112), .Z(new_n1151));
  INV_X1    g726(.A(new_n1019), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1150), .A2(new_n1151), .B1(new_n1152), .B2(new_n994), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1142), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n968), .B1(new_n1119), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n955), .B1(new_n744), .B2(new_n963), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n955), .A2(new_n961), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1158), .A2(KEYINPUT46), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(KEYINPUT46), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1157), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT47), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n796), .A2(new_n798), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n962), .A2(new_n964), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1163), .B1(new_n1164), .B2(new_n966), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1165), .A2(new_n955), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n967), .A2(new_n955), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n957), .A2(new_n955), .ZN(new_n1168));
  XOR2_X1   g743(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1169));
  XNOR2_X1  g744(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1162), .B(new_n1166), .C1(new_n1167), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1156), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g747(.A1(new_n660), .A2(G319), .ZN(new_n1174));
  NOR3_X1   g748(.A1(G229), .A2(G227), .A3(new_n1174), .ZN(new_n1175));
  AND3_X1   g749(.A1(new_n861), .A2(new_n866), .A3(new_n863), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n866), .B1(new_n861), .B2(new_n863), .ZN(new_n1177));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n926), .A2(new_n933), .ZN(new_n1179));
  NOR2_X1   g753(.A1(new_n1178), .A2(new_n1179), .ZN(G308));
  OR2_X1    g754(.A1(new_n1178), .A2(new_n1179), .ZN(G225));
endmodule


