//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G50), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n238), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G13), .ZN(new_n247));
  NOR3_X1   g0047(.A1(new_n247), .A2(new_n207), .A3(G1), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n241), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT12), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n241), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n207), .A2(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n213), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n248), .A2(new_n257), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n206), .A2(G20), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G68), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n250), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT11), .B1(new_n255), .B2(new_n257), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT14), .ZN(new_n266));
  AND2_X1   g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT66), .B1(new_n267), .B2(new_n213), .ZN(new_n268));
  AND2_X1   g0068(.A1(G1), .A2(G13), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n268), .A2(G274), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT67), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n273), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n268), .A2(new_n272), .A3(G274), .A4(new_n277), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT67), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n267), .A2(KEYINPUT66), .A3(new_n213), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n270), .B1(new_n269), .B2(new_n271), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n281), .A2(new_n282), .A3(new_n277), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n278), .A2(new_n280), .B1(G238), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G232), .A3(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G97), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT3), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(G226), .A4(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT69), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n285), .A2(KEYINPUT69), .A3(G226), .A4(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n269), .A2(new_n271), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT13), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n284), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n284), .B2(new_n302), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n266), .B(G169), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n278), .A2(new_n280), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n283), .A2(G238), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n300), .B1(new_n288), .B2(new_n298), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT13), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n284), .A2(new_n303), .A3(new_n302), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(G179), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n312), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n266), .B1(new_n315), .B2(G169), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n265), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(G200), .B1(new_n304), .B2(new_n305), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n311), .A2(G190), .A3(new_n312), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n318), .A2(new_n319), .A3(new_n264), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n259), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT8), .B(G58), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n260), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n247), .A2(G1), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G20), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n323), .A2(new_n326), .B1(new_n328), .B2(new_n325), .ZN(new_n329));
  INV_X1    g0129(.A(new_n257), .ZN(new_n330));
  AND2_X1   g0130(.A1(G58), .A2(G68), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n331), .A2(new_n201), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n291), .A2(KEYINPUT70), .A3(G33), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT70), .B1(new_n291), .B2(G33), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n290), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT7), .B1(new_n337), .B2(new_n207), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT71), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n241), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n291), .A2(G33), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT70), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n289), .B2(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n291), .A2(KEYINPUT70), .A3(G33), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n342), .B1(new_n347), .B2(G20), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n341), .A2(new_n348), .A3(KEYINPUT71), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n334), .B1(new_n340), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n330), .B1(new_n350), .B2(KEYINPUT16), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT73), .B1(new_n289), .B2(KEYINPUT3), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT73), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(new_n291), .A3(G33), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n355), .A3(new_n290), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n342), .B1(new_n356), .B2(new_n207), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n285), .A2(KEYINPUT7), .A3(G20), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n357), .A2(new_n241), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n352), .B1(new_n359), .B2(new_n334), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n329), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n279), .B(new_n274), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n281), .A2(new_n282), .ZN(new_n363));
  INV_X1    g0163(.A(new_n277), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(G232), .A3(new_n364), .ZN(new_n365));
  MUX2_X1   g0165(.A(G223), .B(G226), .S(G1698), .Z(new_n366));
  AOI22_X1  g0166(.A1(new_n347), .A2(new_n366), .B1(G33), .B2(G87), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n367), .B2(new_n300), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT74), .ZN(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AND4_X1   g0172(.A1(G232), .A2(new_n364), .A3(new_n268), .A4(new_n272), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n347), .A2(new_n366), .ZN(new_n374));
  INV_X1    g0174(.A(G87), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n289), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n373), .B1(new_n376), .B2(new_n301), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n307), .A3(new_n371), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT74), .ZN(new_n379));
  INV_X1    g0179(.A(G169), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n362), .B2(new_n368), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n372), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT18), .B1(new_n361), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n378), .B2(KEYINPUT74), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n370), .B1(new_n369), .B2(new_n371), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n349), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n348), .B2(KEYINPUT71), .ZN(new_n388));
  OAI211_X1 g0188(.A(KEYINPUT16), .B(new_n333), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(new_n257), .A3(new_n360), .ZN(new_n390));
  INV_X1    g0190(.A(new_n329), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n386), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n377), .A2(new_n307), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n369), .B2(G200), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n361), .A2(KEYINPUT17), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n390), .A2(new_n391), .A3(new_n397), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n383), .A2(new_n394), .A3(new_n398), .A4(new_n401), .ZN(new_n402));
  XOR2_X1   g0202(.A(KEYINPUT68), .B(G226), .Z(new_n403));
  OR2_X1    g0203(.A1(G222), .A2(G1698), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(G223), .B2(new_n293), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n300), .B1(new_n405), .B2(new_n285), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n290), .A2(new_n292), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n253), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n283), .A2(new_n403), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n307), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G190), .ZN(new_n412));
  INV_X1    g0212(.A(G150), .ZN(new_n413));
  INV_X1    g0213(.A(new_n251), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n324), .A2(new_n254), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n207), .B1(new_n201), .B2(new_n239), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n257), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n239), .B1(new_n206), .B2(G20), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n259), .A2(new_n418), .B1(new_n239), .B2(new_n248), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n417), .A2(KEYINPUT9), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT9), .B1(new_n417), .B2(new_n419), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n410), .A2(G200), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n412), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT10), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT10), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n412), .A2(new_n422), .A3(new_n426), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n285), .A2(G238), .A3(G1698), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n285), .A2(G232), .A3(new_n293), .ZN(new_n431));
  INV_X1    g0231(.A(G107), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n285), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n433), .A2(new_n301), .B1(new_n283), .B2(G244), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n434), .A2(new_n307), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n371), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n325), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n437));
  XOR2_X1   g0237(.A(KEYINPUT15), .B(G87), .Z(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(new_n207), .A3(G33), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n330), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n259), .A2(G77), .A3(new_n260), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(G77), .B2(new_n328), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n436), .B1(G169), .B2(new_n435), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n435), .A2(G190), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n440), .A2(new_n442), .ZN(new_n445));
  INV_X1    g0245(.A(G200), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n444), .B(new_n445), .C1(new_n446), .C2(new_n435), .ZN(new_n447));
  INV_X1    g0247(.A(new_n417), .ZN(new_n448));
  INV_X1    g0248(.A(new_n419), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n410), .B2(new_n380), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(G179), .B2(new_n410), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n443), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n322), .A2(new_n402), .A3(new_n429), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n248), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT83), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n206), .A2(G33), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n330), .A2(new_n328), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G116), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT75), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(KEYINPUT75), .A2(G33), .A3(G283), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n468), .B(new_n207), .C1(G33), .C2(new_n469), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n256), .A2(new_n213), .B1(G20), .B2(new_n455), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT20), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n470), .A2(KEYINPUT20), .A3(new_n471), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n463), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  MUX2_X1   g0275(.A(G257), .B(G264), .S(G1698), .Z(new_n476));
  AOI22_X1  g0276(.A1(new_n347), .A2(new_n476), .B1(G303), .B2(new_n407), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n300), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n268), .A2(G274), .A3(new_n272), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT76), .B1(new_n482), .B2(G41), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT76), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n275), .A3(KEYINPUT5), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n275), .A2(KEYINPUT5), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n206), .A2(G45), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT77), .B1(new_n481), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT77), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n206), .B(G45), .C1(new_n275), .C2(KEYINPUT5), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n483), .B2(new_n485), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n363), .A2(new_n492), .A3(new_n494), .A4(G274), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n276), .A2(G1), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n482), .A2(G41), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n275), .A2(KEYINPUT5), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AND4_X1   g0300(.A1(G270), .A2(new_n500), .A3(new_n268), .A4(new_n272), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n480), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(KEYINPUT82), .B(new_n501), .C1(new_n491), .C2(new_n495), .ZN(new_n504));
  OAI211_X1 g0304(.A(G190), .B(new_n479), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n492), .B1(new_n273), .B2(new_n494), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n481), .A2(new_n490), .A3(KEYINPUT77), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT82), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n496), .A2(new_n480), .A3(new_n502), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n478), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n475), .B(new_n505), .C1(new_n511), .C2(new_n446), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n347), .A2(new_n476), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n407), .A2(G303), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n371), .B1(new_n516), .B2(new_n301), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(new_n474), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n474), .A2(G169), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n511), .A2(new_n519), .A3(KEYINPUT21), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n479), .B1(new_n503), .B2(new_n504), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n473), .A2(new_n472), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n380), .B1(new_n523), .B2(new_n463), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n521), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n512), .B(new_n518), .C1(new_n520), .C2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AND4_X1   g0327(.A1(G257), .A2(new_n500), .A3(new_n268), .A4(new_n272), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n491), .B2(new_n495), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n293), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n468), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G244), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(G1698), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT4), .B1(new_n347), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n301), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n529), .A2(G190), .A3(new_n536), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n357), .A2(new_n432), .A3(new_n358), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n539), .A2(new_n469), .A3(G107), .ZN(new_n540));
  XNOR2_X1  g0340(.A(G97), .B(G107), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI22_X1  g0342(.A1(new_n542), .A2(new_n207), .B1(new_n253), .B2(new_n414), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n257), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n328), .A2(G97), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n461), .B2(G97), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n537), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n536), .ZN(new_n548));
  INV_X1    g0348(.A(new_n528), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n496), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT78), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT78), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n529), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n548), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n547), .B1(new_n554), .B2(new_n446), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n529), .A2(new_n552), .ZN(new_n556));
  AOI211_X1 g0356(.A(KEYINPUT78), .B(new_n528), .C1(new_n491), .C2(new_n495), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n371), .B(new_n536), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n529), .A2(new_n536), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(new_n380), .B1(new_n544), .B2(new_n546), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n438), .A2(new_n328), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n460), .A2(new_n375), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n347), .A2(new_n207), .A3(G68), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n287), .B2(new_n207), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G87), .A2(G97), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n567), .A2(KEYINPUT80), .A3(new_n432), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT80), .B1(new_n567), .B2(new_n432), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n565), .B1(new_n254), .B2(new_n469), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n564), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI211_X1 g0372(.A(new_n562), .B(new_n563), .C1(new_n572), .C2(new_n257), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n497), .A2(G250), .ZN(new_n574));
  OR2_X1    g0374(.A1(new_n488), .A2(G274), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n363), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n289), .A2(new_n455), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G238), .A2(G1698), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n533), .B2(G1698), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n577), .B1(new_n347), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n301), .B1(new_n580), .B2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT79), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n582), .B(new_n577), .C1(new_n347), .C2(new_n579), .ZN(new_n583));
  OAI211_X1 g0383(.A(G190), .B(new_n576), .C1(new_n581), .C2(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n573), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n576), .B1(new_n581), .B2(new_n583), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G200), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n562), .B1(new_n572), .B2(new_n257), .ZN(new_n588));
  XOR2_X1   g0388(.A(new_n438), .B(KEYINPUT81), .Z(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n461), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n586), .A2(new_n380), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n371), .B(new_n576), .C1(new_n581), .C2(new_n583), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n585), .A2(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n555), .A2(new_n561), .A3(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n248), .A2(KEYINPUT25), .A3(new_n432), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT25), .B1(new_n248), .B2(new_n432), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n595), .A2(new_n596), .B1(new_n460), .B2(new_n432), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n347), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT22), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n207), .A2(G87), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n407), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT23), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n432), .A3(G20), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n607), .B(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT24), .B1(new_n602), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n607), .B(KEYINPUT84), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT24), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n611), .A2(new_n612), .A3(new_n598), .A4(new_n601), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n597), .B1(new_n614), .B2(new_n257), .ZN(new_n615));
  MUX2_X1   g0415(.A(G250), .B(G257), .S(G1698), .Z(new_n616));
  NAND2_X1  g0416(.A1(new_n347), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(G294), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n289), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n500), .A2(new_n268), .A3(new_n272), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n621), .A2(new_n301), .B1(G264), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(new_n496), .A3(new_n371), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n500), .A2(new_n268), .A3(G264), .A4(new_n272), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n347), .B2(new_n616), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n300), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n495), .B2(new_n491), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n624), .B1(new_n628), .B2(G169), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n615), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(G200), .B1(new_n623), .B2(new_n496), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT85), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n623), .A2(new_n496), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n631), .A2(new_n632), .B1(new_n633), .B2(G190), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n628), .A2(KEYINPUT85), .A3(G200), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n615), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n594), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n454), .A2(new_n527), .A3(new_n638), .ZN(G372));
  INV_X1    g0439(.A(KEYINPUT86), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n428), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n425), .A2(KEYINPUT86), .A3(new_n427), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n398), .A2(new_n401), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n320), .A2(new_n443), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n317), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n383), .A2(new_n394), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n452), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n555), .A2(new_n636), .A3(new_n593), .A4(new_n561), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n518), .B(new_n630), .C1(new_n520), .C2(new_n525), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n558), .A2(new_n560), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(KEYINPUT26), .A3(new_n593), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n587), .A2(new_n573), .A3(new_n584), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n588), .A2(new_n590), .ZN(new_n657));
  INV_X1    g0457(.A(new_n576), .ZN(new_n658));
  INV_X1    g0458(.A(new_n577), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n533), .A2(G1698), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(G238), .B2(G1698), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n337), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n300), .B1(new_n662), .B2(new_n582), .ZN(new_n663));
  INV_X1    g0463(.A(new_n583), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n658), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n592), .B(new_n657), .C1(new_n665), .C2(G169), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n656), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n655), .B1(new_n561), .B2(new_n667), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n654), .A2(new_n668), .B1(new_n592), .B2(new_n591), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n652), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n454), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n649), .A2(new_n671), .ZN(G369));
  OAI21_X1  g0472(.A(new_n518), .B1(new_n520), .B2(new_n525), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n327), .A2(new_n207), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(G213), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n475), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n526), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n637), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n615), .B2(new_n680), .ZN(new_n687));
  INV_X1    g0487(.A(new_n630), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n679), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT21), .B1(new_n511), .B2(new_n519), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n522), .A2(new_n524), .A3(new_n521), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n679), .B1(new_n694), .B2(new_n518), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n686), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n688), .A2(new_n680), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n691), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n210), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n568), .A2(new_n569), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n455), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n702), .A2(new_n206), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n216), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(new_n702), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  INV_X1    g0508(.A(G330), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n536), .B1(new_n556), .B2(new_n557), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n633), .A2(new_n586), .A3(new_n371), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(new_n522), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n503), .A2(new_n504), .ZN(new_n714));
  OAI21_X1  g0514(.A(G179), .B1(new_n477), .B2(new_n300), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n627), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n665), .A2(new_n536), .A3(new_n529), .A4(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n713), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n623), .A2(new_n517), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n559), .A2(new_n719), .A3(new_n586), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(KEYINPUT30), .A3(new_n513), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n712), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT31), .B1(new_n722), .B2(new_n679), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n527), .A2(new_n638), .A3(new_n680), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n709), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n670), .B2(new_n680), .ZN(new_n729));
  AOI211_X1 g0529(.A(KEYINPUT29), .B(new_n679), .C1(new_n652), .C2(new_n669), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n708), .B1(new_n731), .B2(G1), .ZN(G364));
  NOR2_X1   g0532(.A1(new_n247), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n206), .B1(new_n733), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n702), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n685), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G330), .B2(new_n683), .ZN(new_n738));
  INV_X1    g0538(.A(new_n736), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n213), .B1(G20), .B2(new_n380), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(G20), .A2(G179), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT88), .Z(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G190), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G200), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT89), .Z(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G58), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT91), .B1(G179), .B2(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(KEYINPUT91), .A2(G179), .A3(G200), .ZN(new_n751));
  OAI211_X1 g0551(.A(G20), .B(new_n395), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G159), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(KEYINPUT92), .B(KEYINPUT32), .Z(new_n755));
  XNOR2_X1  g0555(.A(new_n754), .B(new_n755), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n743), .A2(new_n395), .A3(new_n446), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT90), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n757), .A2(KEYINPUT90), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n756), .B1(new_n762), .B2(G77), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n207), .A2(new_n446), .A3(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G190), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n446), .A2(G190), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n743), .A2(new_n766), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n285), .B1(new_n375), .B2(new_n765), .C1(new_n767), .C2(new_n241), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n750), .A2(new_n751), .ZN(new_n769));
  OAI21_X1  g0569(.A(G20), .B1(new_n769), .B2(new_n395), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n768), .B1(G97), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n764), .A2(new_n395), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT93), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT93), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n744), .A2(new_n446), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n775), .A2(G107), .B1(G50), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n748), .A2(new_n763), .A3(new_n771), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n762), .A2(G311), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n745), .A2(G322), .B1(G294), .B2(new_n770), .ZN(new_n780));
  INV_X1    g0580(.A(G303), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n407), .B1(new_n765), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n752), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(G329), .ZN(new_n784));
  INV_X1    g0584(.A(new_n767), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n782), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n775), .A2(G283), .B1(G326), .B2(new_n776), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n779), .A2(new_n780), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n741), .B1(new_n778), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n740), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n701), .A2(new_n407), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G355), .B1(new_n455), .B2(new_n701), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT87), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT87), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n245), .A2(new_n276), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n701), .A2(new_n347), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G45), .B2(new_n216), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n739), .B(new_n790), .C1(new_n794), .C2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n793), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n683), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n738), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  AOI21_X1  g0607(.A(new_n679), .B1(new_n652), .B2(new_n669), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n447), .B1(new_n445), .B2(new_n680), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n443), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n443), .A2(new_n679), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n808), .B(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n727), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n736), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n740), .A2(new_n791), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n739), .B1(new_n253), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n765), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n285), .B1(new_n819), .B2(G107), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  INV_X1    g0621(.A(G283), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n752), .C1(new_n767), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n775), .A2(G87), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G294), .A2(new_n745), .B1(new_n776), .B2(G303), .ZN(new_n825));
  INV_X1    g0625(.A(new_n770), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n824), .B(new_n825), .C1(new_n469), .C2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n823), .B(new_n827), .C1(G116), .C2(new_n762), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT94), .Z(new_n829));
  INV_X1    g0629(.A(new_n776), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n830), .A2(new_n831), .B1(new_n767), .B2(new_n413), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n762), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n746), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT34), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n775), .A2(G68), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n770), .A2(G58), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n783), .A2(G132), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n337), .B1(new_n819), .B2(G50), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT95), .Z(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n836), .B2(KEYINPUT34), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n829), .B1(new_n837), .B2(new_n844), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n818), .B1(new_n792), .B2(new_n812), .C1(new_n845), .C2(new_n741), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n816), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  INV_X1    g0648(.A(new_n542), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n455), .B(new_n215), .C1(new_n849), .C2(KEYINPUT35), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(KEYINPUT35), .B2(new_n849), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT36), .Z(new_n852));
  OR3_X1    g0652(.A1(new_n216), .A2(new_n253), .A3(new_n331), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n206), .B(G13), .C1(new_n853), .C2(new_n240), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n399), .B1(new_n361), .B2(new_n382), .ZN(new_n856));
  XNOR2_X1  g0656(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n361), .B2(new_n677), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT98), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n857), .ZN(new_n860));
  INV_X1    g0660(.A(new_n677), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(new_n392), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT98), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n386), .A2(new_n392), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .A4(new_n399), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n361), .A2(new_n677), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n860), .B1(new_n856), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n402), .A2(new_n867), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT100), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n402), .A2(KEYINPUT100), .A3(new_n867), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n333), .B1(new_n387), .B2(new_n388), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n352), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n329), .B1(new_n351), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT96), .B1(new_n880), .B2(new_n677), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n389), .A2(new_n257), .ZN(new_n882));
  INV_X1    g0682(.A(new_n352), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n350), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n391), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT96), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(new_n861), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n386), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n881), .A2(new_n887), .A3(new_n399), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n866), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n881), .A2(new_n887), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n402), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n876), .A2(new_n877), .A3(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n859), .A2(new_n865), .B1(new_n889), .B2(KEYINPUT37), .ZN(new_n896));
  INV_X1    g0696(.A(new_n893), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n875), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n894), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT39), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(G169), .B1(new_n304), .B2(new_n305), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT14), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n313), .A3(new_n306), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(new_n265), .A3(new_n680), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n265), .A2(new_n679), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n317), .A2(new_n321), .A3(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n265), .B(new_n679), .C1(new_n904), .C2(new_n320), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n670), .A2(new_n680), .A3(new_n812), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n912), .B1(new_n913), .B2(new_n811), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n899), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n861), .B1(new_n383), .B2(new_n394), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT99), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n899), .B2(new_n914), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT99), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n907), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n454), .B1(new_n729), .B2(new_n730), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n649), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n724), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR4_X1   g0727(.A1(new_n526), .A2(new_n594), .A3(new_n637), .A4(new_n679), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n812), .B(new_n911), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT40), .B1(new_n899), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n725), .A2(new_n726), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n932), .A2(KEYINPUT40), .A3(new_n812), .A4(new_n911), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n876), .B2(new_n894), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n932), .A2(new_n454), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n709), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n924), .A2(new_n938), .B1(new_n206), .B2(new_n733), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT101), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n924), .A2(new_n938), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n939), .A2(KEYINPUT101), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n855), .B1(new_n942), .B2(new_n943), .ZN(G367));
  AND2_X1   g0744(.A1(new_n544), .A2(new_n546), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n555), .B(new_n561), .C1(new_n945), .C2(new_n680), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n653), .A2(new_n679), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n691), .A2(KEYINPUT102), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n593), .B1(new_n573), .B2(new_n680), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n666), .A2(new_n573), .A3(new_n680), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT102), .B1(new_n691), .B2(new_n949), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n950), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n955), .B1(new_n950), .B2(new_n956), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n946), .A2(new_n630), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n679), .B1(new_n959), .B2(new_n561), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n948), .A2(new_n686), .A3(new_n695), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n961), .B2(KEYINPUT42), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n962), .A2(new_n963), .B1(KEYINPUT43), .B2(new_n953), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n957), .A2(new_n958), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(new_n957), .B2(new_n958), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n702), .B(KEYINPUT41), .Z(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n696), .B1(new_n690), .B2(new_n695), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n685), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n731), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n684), .B1(new_n687), .B2(new_n689), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT105), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT44), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(KEYINPUT103), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n698), .B2(new_n949), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(KEYINPUT103), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT104), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n981), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n699), .A2(KEYINPUT45), .A3(new_n948), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n698), .B2(new_n949), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n976), .A2(new_n982), .A3(new_n983), .A4(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n974), .A2(new_n975), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n989), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n973), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n731), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n970), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n968), .B1(new_n995), .B2(new_n734), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n951), .A2(new_n793), .A3(new_n952), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n800), .A2(new_n234), .ZN(new_n998));
  INV_X1    g0798(.A(new_n794), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n701), .B2(new_n438), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n739), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n407), .B1(new_n819), .B2(G58), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n831), .B2(new_n752), .C1(new_n767), .C2(new_n753), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G77), .B2(new_n775), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n770), .A2(G68), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n745), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n1006), .B2(new_n413), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1007), .A2(KEYINPUT106), .B1(new_n834), .B2(new_n830), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(KEYINPUT106), .B2(new_n1007), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1004), .B1(new_n239), .B2(new_n761), .C1(new_n1010), .C2(KEYINPUT107), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n746), .A2(new_n781), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT46), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n765), .B2(new_n455), .ZN(new_n1015));
  INV_X1    g0815(.A(G317), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1015), .B1(new_n1016), .B2(new_n752), .C1(new_n767), .C2(new_n618), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n762), .B2(G283), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n765), .A2(new_n1014), .A3(new_n455), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n347), .B(new_n1019), .C1(new_n775), .C2(G97), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n776), .A2(G311), .B1(G107), .B2(new_n770), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1011), .A2(new_n1012), .B1(new_n1013), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n997), .B(new_n1001), .C1(new_n1025), .C2(new_n741), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n996), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(G387));
  NOR2_X1   g0829(.A1(new_n972), .A2(new_n731), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1030), .A2(KEYINPUT111), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(KEYINPUT111), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n702), .B(KEYINPUT110), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1031), .A2(new_n973), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n795), .A2(new_n704), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(G107), .B2(new_n210), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n231), .A2(new_n276), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT109), .Z(new_n1038));
  AOI211_X1 g0838(.A(G45), .B(new_n704), .C1(G68), .C2(G77), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n324), .A2(G50), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n701), .B(new_n347), .C1(new_n1039), .C2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1036), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n736), .B1(new_n1043), .B2(new_n999), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n762), .A2(G68), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G159), .A2(new_n776), .B1(new_n589), .B2(new_n770), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n775), .A2(G97), .B1(G50), .B2(new_n745), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n347), .B1(new_n765), .B2(new_n253), .C1(new_n752), .C2(new_n413), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n325), .B2(new_n785), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n347), .B1(new_n783), .B2(G326), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n775), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n826), .A2(new_n822), .B1(new_n618), .B2(new_n765), .ZN(new_n1053));
  INV_X1    g0853(.A(G322), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n830), .A2(new_n1054), .B1(new_n767), .B2(new_n821), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n762), .B2(G303), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1016), .B2(new_n746), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT48), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1053), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1051), .B1(new_n455), .B2(new_n1052), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1050), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1044), .B1(new_n1064), .B2(new_n740), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n687), .A2(new_n689), .A3(new_n793), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1065), .A2(new_n1066), .B1(new_n972), .B2(new_n735), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1034), .A2(new_n1067), .ZN(G393));
  NAND2_X1  g0868(.A1(new_n991), .A2(new_n992), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n973), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n991), .A2(new_n992), .A3(new_n973), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n1033), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n800), .A2(new_n238), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1074), .B(new_n794), .C1(new_n469), .C2(new_n210), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n285), .B1(new_n819), .B2(G283), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n1054), .B2(new_n752), .C1(new_n767), .C2(new_n781), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1052), .A2(new_n432), .B1(new_n455), .B2(new_n826), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G294), .C2(new_n762), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G311), .A2(new_n745), .B1(new_n776), .B2(G317), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT52), .Z(new_n1081));
  OAI221_X1 g0881(.A(new_n347), .B1(new_n241), .B2(new_n765), .C1(new_n767), .C2(new_n239), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G143), .B2(new_n783), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n770), .A2(G77), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n824), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n325), .B2(new_n762), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G150), .A2(new_n776), .B1(new_n745), .B2(G159), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1079), .A2(new_n1081), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n736), .B(new_n1075), .C1(new_n1090), .C2(new_n741), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n949), .B2(new_n793), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1069), .B2(new_n735), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1073), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(KEYINPUT113), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT113), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1073), .A2(new_n1096), .A3(new_n1093), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(G390));
  INV_X1    g0898(.A(new_n1033), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n727), .A2(new_n454), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n922), .A2(new_n649), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n913), .A2(new_n811), .ZN(new_n1102));
  OAI211_X1 g0902(.A(G330), .B(new_n812), .C1(new_n927), .C2(new_n928), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1103), .A2(new_n912), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n911), .B1(new_n727), .B2(new_n812), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT114), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT114), .B1(new_n909), .B2(new_n910), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1103), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n811), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n808), .B2(new_n812), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n727), .A2(new_n812), .A3(new_n911), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(KEYINPUT116), .B(new_n1101), .C1(new_n1106), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT116), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1101), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n905), .B1(new_n1112), .B2(new_n912), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n895), .A2(new_n900), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1113), .A2(KEYINPUT115), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1109), .A2(new_n1107), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n906), .B1(new_n1124), .B2(new_n1102), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n876), .A2(new_n894), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1122), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1123), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1099), .B1(new_n1120), .B2(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1115), .A2(new_n1119), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT117), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1103), .A2(new_n912), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1112), .B1(new_n1136), .B2(new_n1113), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1118), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(KEYINPUT116), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1117), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1123), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1122), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1131), .B1(new_n1134), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n901), .A2(new_n792), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n817), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n736), .B1(new_n325), .B2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT118), .Z(new_n1152));
  NAND2_X1  g0952(.A1(new_n783), .A2(G125), .ZN(new_n1153));
  OR3_X1    g0953(.A1(new_n765), .A2(KEYINPUT53), .A3(new_n413), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT53), .B1(new_n765), .B2(new_n413), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n285), .B1(new_n831), .B2(new_n767), .C1(new_n1052), .C2(new_n239), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT54), .B(G143), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1156), .B(new_n1157), .C1(new_n762), .C2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n830), .A2(new_n1161), .B1(new_n753), .B2(new_n826), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G132), .B2(new_n745), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n838), .A2(new_n1084), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n455), .A2(new_n1006), .B1(new_n830), .B2(new_n822), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n752), .A2(new_n618), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n407), .B1(new_n375), .B2(new_n765), .C1(new_n767), .C2(new_n432), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(new_n762), .C2(G97), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1160), .A2(new_n1163), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1152), .B1(new_n1170), .B2(new_n741), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1149), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1146), .B2(new_n735), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1148), .A2(new_n1173), .ZN(G378));
  NAND2_X1  g0974(.A1(new_n775), .A2(G58), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n1005), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n432), .A2(new_n1006), .B1(new_n830), .B2(new_n455), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n762), .A2(new_n589), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n337), .A2(new_n275), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n767), .A2(new_n469), .B1(new_n253), .B2(new_n765), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G283), .C2(new_n783), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1178), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT58), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1180), .B(new_n239), .C1(G33), .C2(G41), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n745), .A2(G128), .B1(G150), .B2(new_n770), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n776), .A2(G125), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n785), .A2(G132), .B1(new_n819), .B2(new_n1159), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n762), .B2(G137), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n775), .A2(G159), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1184), .B(new_n1185), .C1(new_n1192), .C2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT119), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n740), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT120), .Z(new_n1200));
  NAND3_X1  g1000(.A1(new_n641), .A2(new_n452), .A3(new_n642), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n450), .A2(new_n677), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1202), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n641), .A2(new_n452), .A3(new_n642), .A4(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1203), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1206), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1208));
  OR3_X1    g1008(.A1(new_n1207), .A2(new_n1208), .A3(new_n792), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n739), .B1(new_n239), .B2(new_n817), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1200), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT121), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1207), .A2(new_n1208), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n935), .B2(G330), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(new_n931), .A2(new_n934), .A3(new_n1213), .A4(new_n709), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n921), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n896), .A2(new_n897), .A3(new_n875), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n875), .B2(new_n874), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n929), .B1(new_n898), .B2(new_n894), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1219), .A2(new_n933), .B1(new_n1220), .B2(KEYINPUT40), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1213), .B1(new_n1221), .B2(new_n709), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n901), .A2(new_n906), .B1(new_n918), .B2(new_n919), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n934), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n899), .A2(new_n930), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT40), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1227), .A3(G330), .A4(new_n1214), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1222), .A2(new_n917), .A3(new_n1223), .A4(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT122), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1217), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n921), .B(KEYINPUT122), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1211), .B1(new_n1233), .B2(new_n734), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1118), .B1(new_n1134), .B2(new_n1147), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1141), .A2(new_n1146), .A3(KEYINPUT117), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1101), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1217), .A2(new_n1229), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT57), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1033), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1235), .B1(new_n1238), .B2(new_n1244), .ZN(G375));
  NAND2_X1  g1045(.A1(new_n1117), .A2(new_n735), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1124), .A2(new_n792), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT123), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n761), .A2(new_n432), .B1(new_n455), .B2(new_n767), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT124), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n407), .B1(new_n765), .B2(new_n469), .C1(new_n752), .C2(new_n781), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G283), .A2(new_n745), .B1(new_n589), .B2(new_n770), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n618), .B2(new_n830), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1251), .B(new_n1253), .C1(G77), .C2(new_n775), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n337), .B1(new_n819), .B2(G159), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n1161), .B2(new_n752), .C1(new_n767), .C2(new_n1158), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1175), .B1(new_n239), .B2(new_n826), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(G150), .C2(new_n762), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n776), .A2(KEYINPUT125), .A3(G132), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT125), .ZN(new_n1260));
  INV_X1    g1060(.A(G132), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n830), .B2(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n747), .A2(G137), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1250), .A2(new_n1254), .B1(new_n1258), .B2(new_n1263), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n736), .B1(G68), .B2(new_n1150), .C1(new_n1264), .C2(new_n741), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1246), .B1(new_n1248), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1106), .A2(new_n1101), .A3(new_n1114), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1120), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n1269), .B2(new_n969), .ZN(G381));
  NOR4_X1   g1070(.A1(G387), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1271));
  INV_X1    g1071(.A(G378), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1243), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1099), .B1(new_n1236), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT57), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1241), .B2(new_n1233), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1234), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(G390), .A2(G381), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1271), .A2(new_n1272), .A3(new_n1277), .A4(new_n1278), .ZN(G407));
  INV_X1    g1079(.A(G213), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(G343), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1272), .A3(new_n1281), .ZN(new_n1282));
  XOR2_X1   g1082(.A(new_n1282), .B(KEYINPUT126), .Z(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1084(.A1(G390), .A2(new_n1028), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1095), .B(new_n1097), .C1(new_n996), .C2(new_n1027), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(new_n806), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1285), .A2(new_n1288), .A3(new_n1286), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G378), .B(new_n1235), .C1(new_n1238), .C2(new_n1244), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1241), .A2(new_n1233), .A3(new_n969), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1242), .A2(new_n735), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1296), .A2(new_n1211), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1272), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT127), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1281), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1268), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1033), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1269), .B2(KEYINPUT60), .ZN(new_n1306));
  OR3_X1    g1106(.A1(new_n1306), .A2(new_n847), .A3(new_n1266), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n847), .B1(new_n1306), .B2(new_n1266), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1236), .A2(new_n1237), .A3(new_n970), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G378), .B1(new_n1311), .B2(new_n1297), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1277), .B2(G378), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT127), .ZN(new_n1314));
  AND4_X1   g1114(.A1(new_n1293), .A2(new_n1302), .A3(new_n1310), .A4(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1281), .A2(G2897), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1309), .A2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1307), .A2(new_n1308), .A3(G2897), .A4(new_n1281), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1313), .B2(new_n1281), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n1281), .B(new_n1309), .C1(new_n1294), .C2(new_n1299), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1320), .B(new_n1321), .C1(new_n1322), .C2(new_n1293), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1292), .B1(new_n1315), .B2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1302), .A2(new_n1310), .A3(new_n1314), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1302), .A2(new_n1314), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1319), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1290), .A2(new_n1321), .A3(new_n1291), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1330), .B1(KEYINPUT63), .B2(new_n1322), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1327), .A2(new_n1329), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1324), .A2(new_n1332), .ZN(G405));
  XNOR2_X1  g1133(.A(new_n1277), .B(new_n1272), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1334), .A2(new_n1309), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1309), .ZN(new_n1336));
  OR3_X1    g1136(.A1(new_n1335), .A2(new_n1336), .A3(new_n1292), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1292), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


