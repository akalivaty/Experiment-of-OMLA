//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  AND2_X1   g001(.A1(KEYINPUT80), .A2(G107), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT80), .A2(G107), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G101), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT71), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G116), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(KEYINPUT71), .A3(G119), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n199), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT5), .ZN(new_n205));
  INV_X1    g019(.A(G113), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT5), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n199), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT70), .B1(new_n209), .B2(new_n206), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT2), .A3(G113), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n210), .A2(new_n212), .B1(new_n209), .B2(new_n206), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n205), .A2(new_n208), .B1(new_n213), .B2(new_n204), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(KEYINPUT79), .B(KEYINPUT3), .C1(new_n192), .C2(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n189), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n192), .A2(KEYINPUT3), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT80), .A2(G107), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT81), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G101), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n192), .A2(G107), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AND4_X1   g043(.A1(KEYINPUT82), .A2(new_n219), .A3(new_n223), .A4(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n217), .A2(new_n218), .B1(new_n190), .B2(new_n221), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT82), .B1(new_n231), .B2(new_n229), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n197), .B(new_n214), .C1(new_n230), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT85), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  INV_X1    g049(.A(new_n218), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT79), .B1(new_n195), .B2(KEYINPUT3), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n223), .B(new_n228), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n235), .B1(new_n238), .B2(G101), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n239), .B1(new_n230), .B2(new_n232), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n213), .B(new_n204), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n235), .A3(G101), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n224), .B1(new_n193), .B2(new_n195), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n219), .A2(new_n223), .A3(new_n229), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT82), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n231), .A2(KEYINPUT82), .A3(new_n229), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT85), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(new_n214), .ZN(new_n251));
  XNOR2_X1  g065(.A(G110), .B(G122), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n234), .A2(new_n243), .A3(new_n251), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT64), .A2(G143), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(G146), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT66), .B1(new_n256), .B2(G146), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n263), .A3(G146), .A4(new_n258), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n254), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n254), .ZN(new_n266));
  NOR2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n256), .B2(G146), .ZN(new_n270));
  INV_X1    g084(.A(G146), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n271), .A2(KEYINPUT65), .A3(G143), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT64), .A2(G143), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT64), .A2(G143), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n268), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n265), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G125), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT86), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G128), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(KEYINPUT1), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n274), .A2(new_n275), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n260), .B1(new_n283), .B2(G146), .ZN(new_n284));
  INV_X1    g098(.A(new_n264), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n273), .A2(new_n276), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT1), .B1(new_n256), .B2(G146), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n290), .A3(new_n279), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n294), .B(G125), .C1(new_n265), .C2(new_n277), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n286), .A2(new_n290), .A3(KEYINPUT88), .A4(new_n279), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n280), .A2(new_n293), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G224), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT7), .B1(new_n298), .B2(G953), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n252), .B(KEYINPUT8), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n249), .A2(new_n214), .ZN(new_n302));
  INV_X1    g116(.A(new_n233), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n253), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n299), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n280), .A2(new_n295), .A3(new_n291), .A4(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(G902), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n234), .A2(new_n243), .A3(new_n251), .ZN(new_n311));
  INV_X1    g125(.A(new_n252), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT6), .A3(new_n253), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n280), .A2(new_n295), .A3(new_n291), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n298), .A2(G953), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT87), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n315), .B(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT6), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n311), .A2(new_n319), .A3(new_n312), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n314), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G210), .B1(G237), .B2(G902), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n310), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n310), .B2(new_n321), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n187), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G478), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(KEYINPUT15), .ZN(new_n327));
  INV_X1    g141(.A(G902), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT9), .B(G234), .ZN(new_n329));
  INV_X1    g143(.A(G217), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n329), .A2(new_n330), .A3(G953), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT96), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n257), .A2(new_n258), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(new_n281), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n283), .A2(KEYINPUT96), .A3(G128), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT13), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(KEYINPUT13), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n281), .A2(G143), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G134), .ZN(new_n342));
  INV_X1    g156(.A(G134), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n336), .A2(new_n343), .A3(new_n340), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n198), .A2(G122), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n198), .A2(G122), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n190), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n191), .A2(new_n347), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n344), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n198), .A2(KEYINPUT14), .A3(G122), .ZN(new_n353));
  OAI211_X1 g167(.A(G107), .B(new_n353), .C1(new_n347), .C2(KEYINPUT14), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n336), .A2(new_n340), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G134), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n357), .B2(new_n344), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n331), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n344), .A2(new_n351), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(G134), .B2(new_n341), .ZN(new_n362));
  INV_X1    g176(.A(new_n331), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n362), .A2(new_n358), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n328), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT97), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n327), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n366), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n352), .A2(new_n359), .A3(new_n331), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n363), .B1(new_n362), .B2(new_n358), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT97), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n367), .B1(new_n373), .B2(new_n327), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G475), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT91), .ZN(new_n377));
  INV_X1    g191(.A(G237), .ZN(new_n378));
  INV_X1    g192(.A(G953), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G143), .A4(G214), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n378), .A2(new_n379), .A3(G214), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT90), .B(new_n380), .C1(new_n333), .C2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n380), .A2(KEYINPUT90), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT18), .A2(G131), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n377), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n380), .A2(KEYINPUT90), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n378), .A2(new_n379), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n283), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n383), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n391), .A2(KEYINPUT91), .A3(KEYINPUT18), .A4(G131), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G125), .B(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n271), .ZN(new_n395));
  INV_X1    g209(.A(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G125), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n279), .A2(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G146), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n385), .A2(new_n386), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT16), .ZN(new_n403));
  OR3_X1    g217(.A1(new_n279), .A2(KEYINPUT16), .A3(G140), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(G146), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(G146), .B1(new_n403), .B2(new_n404), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n391), .A2(KEYINPUT17), .A3(G131), .ZN(new_n409));
  INV_X1    g223(.A(G131), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n385), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n391), .A2(G131), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT95), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n408), .B(new_n409), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n414), .A2(new_n415), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n402), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G113), .B(G122), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(new_n192), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n420), .B(new_n402), .C1(new_n416), .C2(new_n417), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n376), .B1(new_n424), .B2(new_n328), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n394), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT92), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n399), .B1(new_n429), .B2(KEYINPUT19), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n430), .A3(new_n271), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT93), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT93), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n428), .A2(new_n430), .A3(new_n433), .A4(new_n271), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n406), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n411), .A2(new_n412), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n393), .A2(new_n401), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT94), .B1(new_n437), .B2(new_n420), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n436), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n402), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n421), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n423), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n444), .B1(new_n443), .B2(new_n445), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n426), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(G234), .A2(G237), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n450), .A2(G952), .A3(new_n379), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n450), .A2(G902), .A3(G953), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(G898), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR4_X1   g268(.A1(new_n325), .A2(new_n375), .A3(new_n449), .A4(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G221), .B1(new_n329), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G140), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n379), .A2(G227), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT11), .B1(new_n343), .B2(G137), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT11), .ZN(new_n463));
  INV_X1    g277(.A(G137), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(G134), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n462), .A2(new_n465), .B1(new_n343), .B2(G137), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G131), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n465), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n343), .A2(G137), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n410), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT68), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT68), .B1(new_n466), .B2(new_n410), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n247), .A2(new_n248), .ZN(new_n477));
  INV_X1    g291(.A(new_n282), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n262), .B2(new_n264), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n262), .A2(new_n264), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n281), .B1(new_n276), .B2(KEYINPUT1), .ZN(new_n481));
  OAI22_X1  g295(.A1(new_n479), .A2(KEYINPUT83), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n480), .A2(KEYINPUT83), .A3(new_n282), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n477), .B(new_n197), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n197), .B1(new_n230), .B2(new_n232), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n479), .B1(new_n289), .B2(new_n287), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n476), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT12), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT10), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n482), .A2(new_n483), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(new_n491), .B2(new_n485), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n486), .A2(new_n490), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n249), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n240), .A2(new_n278), .A3(new_n242), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n492), .A2(new_n476), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n461), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n495), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n475), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n496), .A3(new_n461), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT84), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT84), .ZN(new_n503));
  INV_X1    g317(.A(new_n496), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n488), .A2(KEYINPUT12), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n506));
  AOI211_X1 g320(.A(new_n506), .B(new_n476), .C1(new_n484), .C2(new_n487), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n504), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n503), .B(new_n500), .C1(new_n509), .C2(new_n461), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n502), .A2(G469), .A3(new_n510), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n484), .A2(new_n490), .B1(new_n493), .B2(new_n249), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n476), .B1(new_n512), .B2(new_n495), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n460), .B1(new_n513), .B2(new_n504), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n488), .A2(KEYINPUT12), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n496), .B(new_n461), .C1(new_n515), .C2(new_n507), .ZN(new_n516));
  AOI211_X1 g330(.A(G469), .B(G902), .C1(new_n514), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G469), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(new_n328), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n457), .B1(new_n511), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n455), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n480), .A2(new_n266), .ZN(new_n523));
  INV_X1    g337(.A(new_n268), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n287), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT67), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT67), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n265), .B2(new_n277), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n475), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n471), .A2(new_n472), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n466), .A2(KEYINPUT68), .A3(new_n410), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT69), .B1(new_n464), .B2(G134), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n343), .A3(G137), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n464), .A2(G134), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n530), .A2(new_n531), .B1(G131), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n286), .A2(new_n290), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT30), .B1(new_n529), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n475), .A2(new_n278), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n541), .A2(new_n539), .A3(KEYINPUT30), .ZN(new_n542));
  INV_X1    g356(.A(new_n241), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n539), .A3(new_n543), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n378), .A2(new_n379), .A3(G210), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT27), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT26), .B(G101), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT31), .B1(new_n544), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n529), .A2(new_n539), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT30), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n278), .A2(new_n475), .B1(new_n537), .B2(new_n538), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT30), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n241), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT31), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n545), .A4(new_n549), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n552), .A2(new_n241), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT28), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n555), .B2(new_n543), .ZN(new_n562));
  AND4_X1   g376(.A1(new_n561), .A2(new_n541), .A3(new_n539), .A4(new_n543), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n549), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n551), .A2(new_n559), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT32), .ZN(new_n568));
  NOR2_X1   g382(.A1(G472), .A2(G902), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n545), .A2(KEYINPUT28), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n555), .A2(new_n561), .A3(new_n543), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n541), .A2(new_n539), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n241), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n549), .A2(KEYINPUT29), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n328), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT72), .B1(new_n564), .B2(new_n565), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT72), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n574), .A2(new_n581), .A3(new_n560), .A4(new_n549), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n557), .A2(new_n545), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT29), .B1(new_n584), .B2(new_n565), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n579), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G472), .ZN(new_n587));
  OAI22_X1  g401(.A1(new_n570), .A2(new_n571), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI221_X1 g404(.A(KEYINPUT73), .B1(new_n586), .B2(new_n587), .C1(new_n570), .C2(new_n571), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n281), .A2(G119), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n201), .A2(G128), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n592), .B1(KEYINPUT74), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(KEYINPUT74), .B2(new_n593), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT24), .B(G110), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT23), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT75), .B1(new_n592), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n593), .A2(KEYINPUT76), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT75), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n601), .B(KEYINPUT23), .C1(new_n281), .C2(G119), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n281), .A2(G119), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT76), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n599), .A2(new_n600), .A3(new_n602), .A4(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n598), .B2(new_n603), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n597), .B1(new_n607), .B2(G110), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n405), .A3(new_n395), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(G110), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n595), .A2(new_n596), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n610), .B(new_n611), .C1(new_n407), .C2(new_n406), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT77), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n612), .A3(KEYINPUT77), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT22), .B(G137), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n379), .A2(G221), .A3(G234), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT78), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n615), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n609), .A2(new_n612), .A3(new_n619), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n328), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT25), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n621), .A2(KEYINPUT25), .A3(new_n328), .A4(new_n622), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n330), .B1(G234), .B2(new_n328), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n621), .A2(new_n622), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n628), .A2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n590), .A2(new_n591), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n522), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n225), .A2(new_n227), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n635), .B(new_n636), .Z(G3));
  AOI21_X1  g451(.A(new_n587), .B1(new_n567), .B2(new_n328), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n569), .B2(new_n567), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n521), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n325), .A2(KEYINPUT98), .ZN(new_n641));
  INV_X1    g455(.A(new_n322), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n314), .A2(new_n318), .A3(new_n320), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n307), .B(KEYINPUT89), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n253), .A2(new_n300), .A3(new_n304), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n328), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n642), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n310), .A2(new_n321), .A3(new_n322), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(new_n650), .A3(new_n187), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n641), .A2(new_n651), .ZN(new_n652));
  OR3_X1    g466(.A1(new_n360), .A2(new_n364), .A3(KEYINPUT33), .ZN(new_n653));
  OAI21_X1  g467(.A(KEYINPUT33), .B1(new_n360), .B2(new_n364), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(G478), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n326), .A2(new_n328), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n371), .B2(new_n326), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n449), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n454), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT99), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n652), .A2(new_n663), .A3(new_n660), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n640), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT100), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT34), .B(G104), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  AOI21_X1  g482(.A(new_n650), .B1(new_n649), .B2(new_n187), .ZN(new_n669));
  INV_X1    g483(.A(new_n187), .ZN(new_n670));
  AOI211_X1 g484(.A(KEYINPUT98), .B(new_n670), .C1(new_n647), .C2(new_n648), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n371), .A2(KEYINPUT97), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n366), .B(G902), .C1(new_n369), .C2(new_n370), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n327), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n367), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n425), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n454), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n446), .A2(KEYINPUT101), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n443), .A2(new_n445), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT20), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(KEYINPUT101), .A3(new_n446), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n677), .A2(new_n678), .A3(new_n679), .A4(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n640), .A2(new_n672), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT35), .B(G107), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G9));
  NAND2_X1  g500(.A1(new_n615), .A2(new_n616), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n620), .A2(KEYINPUT36), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n687), .B(new_n688), .Z(new_n689));
  AOI22_X1  g503(.A1(new_n627), .A2(new_n628), .B1(new_n689), .B2(new_n631), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n455), .A2(new_n521), .A3(new_n639), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT37), .B(G110), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G12));
  AND4_X1   g508(.A1(new_n590), .A2(new_n521), .A3(new_n591), .A4(new_n691), .ZN(new_n695));
  INV_X1    g509(.A(G900), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n451), .B1(new_n452), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n677), .A2(new_n679), .A3(new_n682), .A4(new_n698), .ZN(new_n699));
  AOI211_X1 g513(.A(KEYINPUT102), .B(new_n699), .C1(new_n641), .C2(new_n651), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  INV_X1    g515(.A(new_n699), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n701), .B1(new_n652), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n695), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  XOR2_X1   g519(.A(new_n649), .B(KEYINPUT38), .Z(new_n706));
  XOR2_X1   g520(.A(new_n697), .B(KEYINPUT39), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n521), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n570), .A2(new_n571), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n565), .B1(new_n557), .B2(new_n545), .ZN(new_n712));
  INV_X1    g526(.A(new_n576), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n545), .A2(new_n565), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n328), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(G472), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT103), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n691), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n187), .A3(new_n449), .A4(new_n375), .ZN(new_n719));
  OR4_X1    g533(.A1(new_n706), .A2(new_n709), .A3(new_n710), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n333), .ZN(G45));
  NAND4_X1  g535(.A1(new_n590), .A2(new_n521), .A3(new_n591), .A4(new_n691), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n449), .A2(new_n658), .A3(new_n698), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n652), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n271), .ZN(G48));
  NAND2_X1  g541(.A1(new_n662), .A2(new_n664), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n590), .A2(new_n591), .A3(new_n633), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n496), .A2(new_n461), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n505), .B2(new_n508), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n461), .B1(new_n499), .B2(new_n496), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n328), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G469), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n514), .A2(new_n516), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n518), .A3(new_n328), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n456), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT104), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n734), .A2(new_n739), .A3(new_n456), .A4(new_n736), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n738), .A2(KEYINPUT105), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT105), .B1(new_n738), .B2(new_n740), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n728), .A2(new_n729), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  AOI21_X1  g560(.A(new_n683), .B1(new_n641), .B2(new_n651), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n518), .B1(new_n735), .B2(new_n328), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n517), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n739), .B1(new_n750), .B2(new_n456), .ZN(new_n751));
  INV_X1    g565(.A(new_n740), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n738), .A2(KEYINPUT105), .A3(new_n740), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n729), .A2(new_n747), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G116), .ZN(G18));
  NOR3_X1   g570(.A1(new_n375), .A2(new_n449), .A3(new_n454), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n590), .A2(new_n591), .A3(new_n757), .A4(new_n691), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n740), .B(new_n738), .C1(new_n669), .C2(new_n671), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT106), .B(G119), .Z(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G21));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n375), .A2(new_n449), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n641), .B2(new_n651), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n629), .A2(new_n632), .ZN(new_n766));
  INV_X1    g580(.A(new_n569), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n549), .B1(new_n577), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n768), .B2(new_n577), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n551), .A2(new_n559), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n766), .A2(new_n772), .A3(new_n454), .A4(new_n638), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n743), .A2(new_n763), .A3(new_n765), .A4(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n753), .A2(new_n754), .A3(new_n773), .A4(new_n765), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT108), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G122), .ZN(G24));
  NOR3_X1   g592(.A1(new_n690), .A2(new_n772), .A3(new_n638), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n724), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT109), .B1(new_n759), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n751), .A2(new_n752), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n723), .A2(new_n690), .A3(new_n772), .A4(new_n638), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n652), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G125), .ZN(G27));
  INV_X1    g601(.A(new_n519), .ZN(new_n788));
  OAI211_X1 g602(.A(G469), .B(new_n500), .C1(new_n509), .C2(new_n461), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n736), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n456), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n647), .A2(new_n187), .A3(new_n648), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(KEYINPUT42), .A3(new_n724), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n588), .A2(new_n633), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT110), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n724), .A2(KEYINPUT42), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n798));
  INV_X1    g612(.A(new_n795), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .A4(new_n793), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n791), .A2(new_n766), .A3(new_n792), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n590), .A2(new_n801), .A3(new_n591), .A4(new_n724), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n796), .B(new_n800), .C1(new_n802), .C2(KEYINPUT42), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G131), .ZN(G33));
  NAND4_X1  g618(.A1(new_n801), .A2(new_n590), .A3(new_n591), .A4(new_n702), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n497), .A2(new_n807), .A3(new_n501), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n502), .A2(new_n510), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n518), .B(new_n808), .C1(new_n809), .C2(new_n807), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n519), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  OR3_X1    g626(.A1(new_n811), .A2(new_n812), .A3(KEYINPUT46), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n812), .B1(new_n811), .B2(KEYINPUT46), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n517), .B1(new_n811), .B2(KEYINPUT46), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n792), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n639), .A2(new_n690), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n425), .B1(new_n681), .B2(new_n446), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n658), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT43), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT43), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n658), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n817), .B1(new_n825), .B2(KEYINPUT44), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(KEYINPUT44), .B2(new_n825), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n816), .A2(new_n827), .A3(new_n456), .A4(new_n707), .ZN(new_n828));
  XNOR2_X1  g642(.A(KEYINPUT112), .B(G137), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(G39));
  NAND2_X1  g644(.A1(new_n590), .A2(new_n591), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n633), .A2(new_n723), .A3(new_n792), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n816), .A2(KEYINPUT47), .A3(new_n456), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT47), .B1(new_n816), .B2(new_n456), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G140), .ZN(G42));
  NOR3_X1   g650(.A1(new_n751), .A2(new_n752), .A3(new_n792), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n821), .A2(new_n451), .A3(new_n823), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n795), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT48), .Z(new_n841));
  NOR3_X1   g655(.A1(new_n766), .A2(new_n638), .A3(new_n772), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n759), .ZN(new_n844));
  INV_X1    g658(.A(G952), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n844), .A2(new_n845), .A3(G953), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n711), .A2(new_n717), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n837), .A2(new_n633), .A3(new_n451), .A4(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n841), .B(new_n846), .C1(new_n659), .C2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n843), .A2(new_n792), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n833), .A2(new_n834), .ZN(new_n853));
  INV_X1    g667(.A(new_n750), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n456), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT118), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n852), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n706), .A2(new_n782), .A3(new_n670), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n858), .A2(new_n843), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n449), .A2(new_n658), .ZN(new_n868));
  INV_X1    g682(.A(new_n779), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n849), .A2(new_n868), .B1(new_n839), .B2(new_n869), .ZN(new_n870));
  OR4_X1    g684(.A1(new_n857), .A2(new_n865), .A3(new_n867), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n855), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n852), .B1(new_n853), .B2(new_n872), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n863), .A2(new_n870), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n850), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n722), .A2(new_n725), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n791), .A2(new_n697), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n765), .A2(new_n718), .A3(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n786), .A2(new_n704), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT52), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n659), .B1(new_n449), .B2(new_n374), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n187), .A3(new_n649), .A4(new_n678), .ZN(new_n883));
  OAI221_X1 g697(.A(new_n692), .B1(new_n883), .B2(new_n640), .C1(new_n634), .C2(new_n522), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n783), .A2(new_n793), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n805), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n425), .A2(new_n697), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n374), .A2(new_n682), .A3(new_n679), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n817), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n374), .A2(new_n682), .A3(new_n679), .A4(new_n887), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT114), .B1(new_n891), .B2(new_n792), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n722), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT115), .B1(new_n886), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n890), .A2(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n695), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT115), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n805), .A4(new_n885), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n884), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n729), .A2(new_n754), .A3(new_n753), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n664), .B2(new_n662), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n760), .A2(new_n755), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n900), .A2(new_n904), .A3(new_n777), .A4(new_n803), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT53), .B1(new_n881), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n895), .A2(new_n899), .ZN(new_n907));
  INV_X1    g721(.A(new_n884), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n760), .A2(new_n755), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n777), .A2(new_n910), .A3(new_n744), .A4(new_n803), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT52), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(KEYINPUT116), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n880), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT102), .B1(new_n672), .B2(new_n699), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n652), .A2(new_n701), .A3(new_n702), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n726), .B1(new_n918), .B2(new_n695), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n786), .A3(new_n879), .A4(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT53), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n912), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n906), .A2(new_n924), .A3(KEYINPUT54), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n923), .B1(new_n881), .B2(new_n905), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT117), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n904), .A2(new_n927), .A3(new_n777), .A4(new_n803), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n911), .A2(KEYINPUT117), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n923), .B(new_n884), .C1(new_n895), .C2(new_n899), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n922), .A2(new_n928), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n876), .A2(new_n925), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(G952), .B2(G953), .ZN(new_n935));
  NOR4_X1   g749(.A1(new_n766), .A2(new_n820), .A3(new_n457), .A4(new_n670), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT49), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n750), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT113), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n847), .B1(new_n937), .B2(new_n750), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n706), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n935), .A2(new_n941), .ZN(G75));
  NOR2_X1   g756(.A1(new_n379), .A2(G952), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n328), .B1(new_n926), .B2(new_n931), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT56), .B1(new_n945), .B2(G210), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n314), .A2(new_n320), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n318), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT55), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n944), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n946), .B2(new_n949), .ZN(G51));
  XNOR2_X1  g765(.A(new_n932), .B(KEYINPUT54), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n519), .B(KEYINPUT57), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n735), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n945), .A2(new_n810), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n943), .B1(new_n955), .B2(new_n956), .ZN(G54));
  NAND3_X1  g771(.A1(new_n945), .A2(KEYINPUT58), .A3(G475), .ZN(new_n958));
  INV_X1    g772(.A(new_n443), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n960), .A2(new_n961), .A3(new_n943), .ZN(G60));
  NAND2_X1  g776(.A1(new_n653), .A2(new_n654), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n656), .B(KEYINPUT59), .Z(new_n964));
  AND3_X1   g778(.A1(new_n952), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n933), .A2(new_n925), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n963), .B1(new_n966), .B2(new_n964), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n965), .A2(new_n967), .A3(new_n943), .ZN(G63));
  NAND2_X1  g782(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AND4_X1   g786(.A1(new_n922), .A2(new_n928), .A3(new_n929), .A4(new_n930), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n880), .B(new_n913), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT53), .B1(new_n912), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n972), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n630), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n969), .B1(new_n978), .B2(KEYINPUT124), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT122), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n980), .A2(new_n932), .A3(new_n689), .A4(new_n972), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n971), .B1(new_n926), .B2(new_n931), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n982), .B2(new_n689), .ZN(new_n983));
  OAI221_X1 g797(.A(new_n979), .B1(KEYINPUT124), .B2(new_n978), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n944), .B1(new_n982), .B2(new_n630), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n932), .A2(new_n689), .A3(new_n972), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT122), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n982), .A2(new_n980), .A3(new_n689), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g803(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n989), .A2(KEYINPUT123), .A3(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT123), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n943), .B1(new_n976), .B2(new_n977), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n981), .B2(new_n983), .ZN(new_n994));
  INV_X1    g808(.A(new_n990), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n984), .B1(new_n991), .B2(new_n996), .ZN(G66));
  INV_X1    g811(.A(new_n453), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n379), .B1(new_n998), .B2(G224), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n904), .A2(new_n777), .A3(new_n908), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(new_n379), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n947), .B1(G898), .B2(new_n379), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1001), .B(new_n1002), .Z(G69));
  NAND2_X1  g817(.A1(G227), .A2(G900), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n379), .A2(G900), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n672), .A2(new_n764), .A3(new_n795), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n816), .A2(new_n456), .A3(new_n707), .A4(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT125), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n919), .A2(new_n786), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n828), .A2(new_n803), .A3(new_n805), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1008), .A2(new_n835), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1005), .B1(new_n1011), .B2(new_n379), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT126), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n554), .A2(new_n556), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n428), .A2(new_n430), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  OAI211_X1 g832(.A(G953), .B(new_n1004), .C1(new_n1014), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1011), .A2(new_n379), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1005), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1013), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g836(.A(KEYINPUT126), .B(new_n1005), .C1(new_n1011), .C2(new_n379), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1017), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1004), .A2(G953), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1009), .A2(new_n720), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1028));
  INV_X1    g842(.A(new_n708), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n729), .A2(new_n1029), .A3(new_n817), .A4(new_n882), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n828), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1027), .A2(new_n835), .A3(new_n1028), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1018), .B1(new_n1033), .B2(G953), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1024), .A2(new_n1025), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1019), .A2(new_n1035), .ZN(G72));
  NAND2_X1  g850(.A1(G472), .A2(G902), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT63), .Z(new_n1038));
  OAI21_X1  g852(.A(new_n1038), .B1(new_n1011), .B2(new_n1000), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n544), .A2(new_n714), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT127), .Z(new_n1041));
  AOI21_X1  g855(.A(new_n943), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1038), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n712), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n906), .A2(new_n924), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1038), .B1(new_n1032), .B2(new_n1000), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n712), .ZN(new_n1047));
  AND3_X1   g861(.A1(new_n1042), .A2(new_n1045), .A3(new_n1047), .ZN(G57));
endmodule


