//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G101), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT3), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT75), .A2(G107), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT75), .A2(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n189), .B1(new_n194), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT4), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT75), .A2(G107), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT75), .A2(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n205), .A2(new_n191), .B1(new_n198), .B2(new_n197), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT76), .B1(new_n206), .B2(new_n189), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n194), .A2(new_n199), .A3(KEYINPUT76), .A4(new_n189), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n202), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT77), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G116), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n201), .A2(new_n200), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n210), .A2(new_n211), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n211), .B1(new_n210), .B2(new_n220), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n192), .A2(new_n193), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n190), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n189), .B1(new_n224), .B2(new_n198), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n194), .A2(new_n199), .A3(new_n189), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT76), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n225), .B1(new_n228), .B2(new_n208), .ZN(new_n229));
  INV_X1    g043(.A(G113), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n214), .A2(G119), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT5), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT5), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n233), .A2(KEYINPUT78), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT78), .B1(new_n233), .B2(new_n234), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n216), .A2(new_n217), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT79), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n229), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n239), .B1(new_n229), .B2(new_n238), .ZN(new_n241));
  OAI22_X1  g055(.A1(new_n221), .A2(new_n222), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G110), .B(G122), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT4), .B1(new_n206), .B2(new_n189), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n228), .B2(new_n208), .ZN(new_n247));
  INV_X1    g061(.A(new_n220), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT77), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n210), .A2(new_n211), .A3(new_n220), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n238), .ZN(new_n252));
  INV_X1    g066(.A(new_n225), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n207), .B2(new_n209), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT79), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n229), .A2(new_n238), .A3(new_n239), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n251), .A2(new_n257), .A3(new_n243), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n245), .A2(KEYINPUT6), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n242), .A2(new_n260), .A3(new_n244), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT64), .A2(G143), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(G146), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT65), .B1(new_n263), .B2(G146), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n264), .A2(new_n270), .A3(G146), .A4(new_n265), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n273), .ZN(new_n277));
  INV_X1    g091(.A(G146), .ZN(new_n278));
  AND2_X1   g092(.A1(KEYINPUT64), .A2(G143), .ZN(new_n279));
  NOR2_X1   g093(.A1(KEYINPUT64), .A2(G143), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n263), .A2(G146), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n277), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n275), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT80), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(G125), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n283), .B1(new_n272), .B2(new_n274), .ZN(new_n288));
  INV_X1    g102(.A(G125), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT80), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT1), .B1(new_n263), .B2(G146), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n281), .A2(new_n282), .B1(G128), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G128), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(KEYINPUT1), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n272), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n289), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n287), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G224), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(G953), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n297), .B(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n259), .A2(new_n261), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n297), .B1(new_n302), .B2(new_n299), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n299), .A2(new_n302), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n287), .A2(new_n290), .A3(new_n296), .A4(new_n304), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n233), .A2(new_n234), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n229), .B1(new_n237), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n243), .B(KEYINPUT8), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n307), .B(new_n308), .C1(new_n229), .C2(new_n252), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n303), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(G902), .B1(new_n310), .B2(new_n258), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n301), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G210), .B1(G237), .B2(G902), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n301), .A2(new_n311), .A3(new_n313), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n188), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(KEYINPUT18), .A2(G131), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  INV_X1    g134(.A(G953), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G214), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n322), .A2(new_n264), .A3(new_n323), .A4(new_n265), .ZN(new_n324));
  INV_X1    g138(.A(G214), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n325), .A2(G237), .A3(G953), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G143), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n279), .A2(new_n280), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n323), .B1(new_n329), .B2(new_n322), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n319), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n289), .A2(G140), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT70), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n289), .A2(KEYINPUT70), .A3(G140), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(G146), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n333), .A2(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n278), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT64), .B(G143), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT81), .B1(new_n341), .B2(new_n326), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n342), .A2(new_n318), .A3(new_n327), .A4(new_n324), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n331), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT82), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n331), .A2(KEYINPUT82), .A3(new_n340), .A4(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G113), .B(G122), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(new_n190), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT16), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT16), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n333), .A2(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n351), .A2(new_n278), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n278), .B1(new_n351), .B2(new_n353), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G131), .B1(new_n328), .B2(new_n330), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT17), .ZN(new_n358));
  INV_X1    g172(.A(G131), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n342), .A2(new_n359), .A3(new_n327), .A4(new_n324), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(KEYINPUT17), .B(G131), .C1(new_n328), .C2(new_n330), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n356), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n348), .A2(new_n350), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n350), .B1(new_n348), .B2(new_n363), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT85), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n343), .A2(new_n340), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT82), .B1(new_n367), .B2(new_n331), .ZN(new_n368));
  INV_X1    g182(.A(new_n347), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n350), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(KEYINPUT85), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G902), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT86), .B1(new_n366), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n371), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n348), .A2(new_n350), .A3(new_n363), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(G902), .B1(new_n365), .B2(KEYINPUT85), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(G475), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n384));
  NOR2_X1   g198(.A1(G475), .A2(G902), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n357), .A2(new_n360), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT83), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n357), .A2(new_n388), .A3(new_n360), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n333), .A2(new_n334), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT19), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n335), .A2(new_n336), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n392), .B1(new_n393), .B2(new_n391), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n355), .B1(new_n394), .B2(new_n278), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n387), .A2(new_n389), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n350), .B1(new_n348), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n384), .B(new_n385), .C1(new_n364), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT84), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n351), .A2(new_n353), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G146), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n391), .B1(new_n335), .B2(new_n336), .ZN(new_n402));
  INV_X1    g216(.A(new_n392), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n278), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(KEYINPUT83), .B2(new_n386), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n406), .A2(new_n389), .B1(new_n346), .B2(new_n347), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n378), .B1(new_n407), .B2(new_n350), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n384), .A4(new_n385), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n385), .B1(new_n364), .B2(new_n397), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT20), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n399), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n264), .A2(G128), .A3(new_n265), .ZN(new_n414));
  INV_X1    g228(.A(G134), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n263), .A2(G128), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G122), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT88), .B1(new_n420), .B2(G116), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT88), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n214), .A3(G122), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(KEYINPUT87), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G122), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n214), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n223), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n427), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G116), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n423), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n205), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n419), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT13), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n414), .B1(new_n435), .B2(new_n416), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n279), .A2(new_n280), .A3(new_n293), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT13), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT89), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G134), .B1(new_n436), .B2(new_n439), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n434), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n415), .B1(new_n414), .B2(new_n417), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n419), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G134), .B1(new_n437), .B2(new_n416), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n418), .A3(KEYINPUT90), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n433), .A2(KEYINPUT91), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT91), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n431), .A2(new_n450), .A3(new_n205), .A4(new_n432), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT14), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n421), .B2(new_n423), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n452), .A2(new_n454), .A3(new_n428), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n449), .B(new_n451), .C1(new_n455), .C2(new_n196), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n442), .B1(new_n448), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT9), .B(G234), .ZN(new_n458));
  INV_X1    g272(.A(G217), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n458), .A2(new_n459), .A3(G953), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n442), .B(new_n460), .C1(new_n448), .C2(new_n456), .ZN(new_n463));
  AOI21_X1  g277(.A(G902), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G478), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(KEYINPUT15), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n464), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(G234), .A2(G237), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n468), .A2(G952), .A3(new_n321), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(G902), .A3(G953), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT92), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(G898), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AND4_X1   g288(.A1(new_n383), .A2(new_n413), .A3(new_n467), .A4(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G221), .B1(new_n458), .B2(G902), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G469), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(new_n373), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n200), .A2(new_n201), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n275), .A2(new_n284), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT10), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n267), .B1(new_n329), .B2(G146), .ZN(new_n483));
  INV_X1    g297(.A(new_n271), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n294), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n292), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n481), .A2(new_n210), .B1(new_n487), .B2(new_n229), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n293), .B1(new_n281), .B2(KEYINPUT1), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n485), .B1(new_n272), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n229), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n482), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n415), .A2(G137), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT11), .ZN(new_n494));
  INV_X1    g308(.A(G137), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(G134), .B2(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n415), .A2(KEYINPUT11), .A3(G137), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G131), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n359), .B(new_n493), .C1(new_n496), .C2(new_n497), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n488), .A2(new_n492), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G110), .B(G140), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT73), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n321), .A2(G227), .ZN(new_n506));
  XOR2_X1   g320(.A(new_n505), .B(new_n506), .Z(new_n507));
  NAND2_X1  g321(.A1(new_n254), .A2(new_n295), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n502), .B1(new_n508), .B2(new_n491), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT12), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT12), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n511), .B(new_n502), .C1(new_n508), .C2(new_n491), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n503), .B(new_n507), .C1(new_n510), .C2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n507), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n288), .A2(new_n480), .ZN(new_n515));
  INV_X1    g329(.A(new_n294), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n269), .B2(new_n271), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT10), .B1(new_n517), .B2(new_n292), .ZN(new_n518));
  OAI22_X1  g332(.A1(new_n247), .A2(new_n515), .B1(new_n254), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT10), .B1(new_n490), .B2(new_n229), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n519), .A2(new_n501), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n502), .B1(new_n488), .B2(new_n492), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n514), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(G902), .B1(new_n513), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n479), .B1(new_n524), .B2(new_n478), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n521), .A2(new_n514), .ZN(new_n526));
  INV_X1    g340(.A(new_n522), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n509), .A2(KEYINPUT12), .ZN(new_n529));
  INV_X1    g343(.A(new_n512), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n507), .B(KEYINPUT74), .Z(new_n532));
  OAI211_X1 g346(.A(new_n528), .B(G469), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n477), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n317), .A2(new_n475), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n459), .B1(G234), .B2(new_n373), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n212), .A2(G128), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n293), .A2(G119), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n538), .B2(new_n539), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT24), .B(G110), .ZN(new_n543));
  OR3_X1    g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n293), .A2(KEYINPUT23), .A3(G119), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n212), .A2(G128), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n538), .B(new_n545), .C1(new_n546), .C2(KEYINPUT23), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G110), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n544), .B(new_n548), .C1(new_n354), .C2(new_n355), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n543), .B1(new_n541), .B2(new_n542), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(G110), .B2(new_n547), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n401), .A3(new_n339), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n321), .A2(G221), .A3(G234), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT71), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT22), .B(G137), .Z(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n553), .B1(new_n549), .B2(new_n552), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n549), .A2(new_n552), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n562), .A2(new_n553), .A3(new_n558), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n373), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT25), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n560), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n554), .A3(new_n558), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n559), .A2(new_n560), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT25), .B1(new_n570), .B2(new_n373), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n537), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n537), .A2(G902), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n320), .A2(new_n321), .A3(G210), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n577), .B(KEYINPUT27), .Z(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT26), .B(G101), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT28), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT67), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT66), .B1(new_n495), .B2(G134), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT66), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n415), .A3(G137), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n495), .A2(G134), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G131), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n500), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n582), .B1(new_n295), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n501), .A2(new_n275), .A3(new_n284), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n588), .A2(new_n500), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n592), .B(KEYINPUT67), .C1(new_n517), .C2(new_n292), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n218), .A2(new_n219), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n589), .B1(new_n485), .B2(new_n486), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n501), .B2(new_n288), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT68), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n218), .A2(KEYINPUT68), .A3(new_n219), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n581), .B1(new_n596), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n500), .B(new_n588), .C1(new_n517), .C2(new_n292), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n591), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n602), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(KEYINPUT28), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n580), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT30), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n593), .A2(new_n591), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n597), .A2(KEYINPUT67), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n591), .A2(new_n605), .A3(KEYINPUT30), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n616), .A3(new_n595), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT31), .ZN(new_n618));
  INV_X1    g432(.A(new_n580), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n603), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n615), .B1(new_n611), .B2(new_n594), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n608), .B1(new_n622), .B2(new_n595), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n618), .B1(new_n623), .B2(new_n619), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n576), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT32), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT32), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n627), .B(new_n576), .C1(new_n621), .C2(new_n624), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n623), .A2(new_n580), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n619), .B1(new_n604), .B2(new_n609), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT29), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n602), .B1(new_n591), .B2(new_n605), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT28), .B1(new_n608), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n603), .A2(new_n581), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT29), .A4(new_n619), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n373), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n632), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n575), .B1(new_n629), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n536), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G101), .ZN(G3));
  OAI21_X1  g455(.A(new_n373), .B1(new_n621), .B2(new_n624), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n617), .A2(new_n603), .A3(new_n619), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT31), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n620), .A3(new_n610), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n642), .A2(G472), .B1(new_n576), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n572), .A2(new_n574), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n534), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n301), .A2(new_n311), .A3(new_n313), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n313), .B1(new_n301), .B2(new_n311), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n187), .B(new_n474), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n383), .A2(new_n413), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n465), .A2(G902), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT93), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n463), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n463), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n445), .A2(new_n447), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n431), .B1(new_n424), .B2(new_n453), .ZN(new_n660));
  OAI21_X1  g474(.A(G107), .B1(new_n660), .B2(new_n452), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n659), .A2(new_n661), .A3(new_n449), .A4(new_n451), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n460), .B1(new_n662), .B2(new_n442), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n657), .B(KEYINPUT33), .C1(new_n658), .C2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT33), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n462), .B(new_n463), .C1(new_n656), .C2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n655), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT94), .B1(new_n464), .B2(G478), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI211_X1 g483(.A(KEYINPUT94), .B(new_n655), .C1(new_n664), .C2(new_n666), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n653), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n652), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n649), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT34), .B(G104), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT95), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n674), .B(new_n676), .ZN(G6));
  INV_X1    g491(.A(new_n466), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n464), .B(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n398), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n384), .B1(new_n408), .B2(new_n385), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n383), .B(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(KEYINPUT96), .B1(new_n652), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT96), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n379), .A2(new_n381), .A3(new_n380), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n381), .B1(new_n379), .B2(new_n380), .ZN(new_n687));
  INV_X1    g501(.A(G475), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n317), .A2(new_n684), .A3(new_n474), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n649), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT35), .B(G107), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G9));
  OAI21_X1  g509(.A(new_n187), .B1(new_n650), .B2(new_n651), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n513), .A2(new_n523), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n478), .A3(new_n373), .ZN(new_n698));
  INV_X1    g512(.A(new_n479), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n533), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n476), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n645), .A2(new_n576), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n564), .A2(new_n565), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n570), .A2(KEYINPUT25), .A3(new_n373), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OR3_X1    g520(.A1(new_n558), .A2(KEYINPUT97), .A3(KEYINPUT36), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT97), .B1(new_n558), .B2(KEYINPUT36), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n562), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n706), .A2(new_n537), .B1(new_n573), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(G472), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n645), .B2(new_n373), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n703), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n702), .A2(new_n714), .A3(new_n475), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT37), .B(G110), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT98), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n715), .B(new_n717), .ZN(G12));
  AOI21_X1  g532(.A(new_n711), .B1(new_n629), .B2(new_n638), .ZN(new_n719));
  INV_X1    g533(.A(G900), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n469), .B1(new_n471), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n682), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n702), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G128), .ZN(G30));
  AND3_X1   g538(.A1(new_n399), .A2(new_n412), .A3(new_n410), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n679), .B1(new_n689), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n710), .A2(new_n573), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n572), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n726), .A2(new_n188), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT99), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n315), .A2(new_n316), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT38), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n623), .A2(new_n580), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n608), .A2(new_n633), .ZN(new_n735));
  AOI21_X1  g549(.A(G902), .B1(new_n735), .B2(new_n580), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G472), .ZN(new_n738));
  INV_X1    g552(.A(new_n628), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n627), .B1(new_n645), .B2(new_n576), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(new_n721), .B(KEYINPUT39), .Z(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  OR3_X1    g557(.A1(new_n701), .A2(KEYINPUT40), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT40), .B1(new_n701), .B2(new_n743), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n732), .A2(new_n741), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n730), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n329), .ZN(G45));
  NAND2_X1  g562(.A1(new_n664), .A2(new_n666), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT94), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n654), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n667), .B2(new_n668), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n383), .B2(new_n413), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT100), .ZN(new_n754));
  INV_X1    g568(.A(new_n721), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n753), .A2(new_n317), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n653), .A2(new_n671), .A3(new_n755), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT100), .B1(new_n757), .B2(new_n696), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n756), .A2(new_n758), .A3(new_n719), .A4(new_n534), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G146), .ZN(G48));
  OAI21_X1  g574(.A(new_n638), .B1(new_n739), .B2(new_n740), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n524), .A2(new_n478), .ZN(new_n762));
  AOI211_X1 g576(.A(G469), .B(G902), .C1(new_n513), .C2(new_n523), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n762), .A2(new_n763), .A3(new_n477), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n761), .A2(new_n647), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n673), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT41), .B(G113), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT101), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n766), .B(new_n768), .ZN(G15));
  NAND2_X1  g583(.A1(new_n692), .A2(new_n765), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G116), .ZN(G18));
  INV_X1    g585(.A(KEYINPUT102), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n524), .A2(new_n478), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n476), .A3(new_n698), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n772), .B1(new_n696), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n317), .A2(KEYINPUT102), .A3(new_n764), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n761), .A2(new_n475), .A3(new_n728), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT103), .B(G119), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(G21));
  AOI21_X1  g595(.A(KEYINPUT106), .B1(new_n653), .B2(new_n679), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n783), .B(new_n467), .C1(new_n383), .C2(new_n413), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n696), .A2(new_n774), .A3(new_n473), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n576), .B(KEYINPUT104), .Z(new_n787));
  INV_X1    g601(.A(new_n620), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n619), .B1(new_n634), .B2(new_n635), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(KEYINPUT31), .B2(new_n643), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT105), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT105), .B1(new_n624), .B2(new_n789), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n787), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n575), .A3(new_n713), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n785), .A2(new_n786), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G122), .ZN(G24));
  NOR4_X1   g611(.A1(new_n757), .A2(new_n794), .A3(new_n713), .A4(new_n711), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n777), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G125), .ZN(G27));
  INV_X1    g614(.A(KEYINPUT42), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n650), .A2(new_n651), .A3(new_n188), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n761), .A2(new_n647), .A3(new_n534), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n801), .B1(new_n803), .B2(new_n757), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n653), .A2(new_n671), .A3(new_n755), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n315), .A2(new_n187), .A3(new_n316), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n701), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n639), .A2(KEYINPUT42), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G131), .ZN(G33));
  INV_X1    g624(.A(new_n803), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n722), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G134), .ZN(G36));
  OAI21_X1  g627(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n478), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(KEYINPUT46), .A3(new_n699), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT107), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n817), .A2(KEYINPUT107), .A3(KEYINPUT46), .A4(new_n699), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(KEYINPUT108), .A3(new_n698), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT46), .ZN(new_n823));
  INV_X1    g637(.A(new_n817), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n823), .B1(new_n824), .B2(new_n479), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n821), .A2(new_n698), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT108), .B1(new_n827), .B2(new_n820), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n476), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n743), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n653), .A2(new_n752), .A3(KEYINPUT43), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT43), .B1(new_n653), .B2(new_n752), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n646), .A2(new_n711), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(KEYINPUT44), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT44), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n806), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n830), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G137), .ZN(G39));
  NOR4_X1   g654(.A1(new_n761), .A2(new_n757), .A3(new_n806), .A4(new_n647), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT47), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n829), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT108), .ZN(new_n844));
  INV_X1    g658(.A(new_n820), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n821), .A2(new_n698), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n825), .A3(new_n822), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT47), .B1(new_n848), .B2(new_n476), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n841), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(G140), .ZN(G42));
  AND3_X1   g665(.A1(new_n831), .A2(new_n469), .A3(new_n832), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n806), .A2(new_n774), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n639), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT48), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n852), .A2(new_n795), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n777), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n321), .A2(G952), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n626), .A2(new_n628), .B1(G472), .B2(new_n737), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n647), .A2(new_n853), .A3(new_n469), .A4(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n858), .B1(new_n860), .B2(new_n753), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n857), .A2(KEYINPUT117), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT117), .B1(new_n857), .B2(new_n861), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n855), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT118), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n855), .B(new_n866), .C1(new_n862), .C2(new_n863), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n794), .A2(new_n713), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n852), .A2(new_n728), .A3(new_n868), .A4(new_n853), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n860), .A2(new_n383), .A3(new_n413), .A4(new_n752), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n764), .A2(new_n188), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT115), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n732), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n856), .A2(new_n873), .A3(KEYINPUT50), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT50), .B1(new_n856), .B2(new_n873), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n869), .B(new_n870), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n829), .A2(new_n842), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n848), .A2(KEYINPUT47), .A3(new_n476), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n762), .A2(new_n763), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n477), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n856), .A2(new_n802), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT114), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n876), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n865), .B(new_n867), .C1(new_n884), .C2(KEYINPUT51), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(KEYINPUT51), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT116), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n884), .A2(new_n888), .A3(KEYINPUT51), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n885), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT110), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n726), .A2(new_n783), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n653), .A2(KEYINPUT106), .A3(new_n679), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n317), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n728), .A2(new_n721), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n741), .A2(new_n534), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n892), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n711), .A2(new_n700), .A3(new_n476), .A4(new_n755), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n859), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n785), .A3(KEYINPUT110), .A4(new_n317), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n799), .A2(new_n759), .A3(new_n723), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n891), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n759), .A2(new_n723), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n898), .A2(new_n901), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n905), .A2(KEYINPUT52), .A3(new_n906), .A4(new_n799), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n868), .A2(new_n728), .A3(new_n805), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n467), .B(new_n755), .C1(new_n680), .C2(new_n681), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n689), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n761), .A2(new_n911), .A3(new_n728), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n807), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n809), .A2(new_n812), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n646), .A2(new_n728), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n383), .A2(new_n413), .A3(new_n679), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(new_n731), .A3(new_n187), .A4(new_n474), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n535), .A2(new_n916), .B1(new_n918), .B2(new_n648), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT109), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n917), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n652), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n649), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n715), .A3(KEYINPUT109), .ZN(new_n925));
  AOI22_X1  g739(.A1(new_n536), .A2(new_n639), .B1(new_n649), .B2(new_n673), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n921), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n770), .A2(new_n779), .A3(new_n766), .A4(new_n796), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n915), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n908), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT53), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n904), .A2(new_n907), .A3(KEYINPUT111), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT53), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT111), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n934), .B(new_n891), .C1(new_n902), .C2(new_n903), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n932), .A2(new_n933), .A3(new_n929), .A4(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n931), .A2(KEYINPUT54), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT112), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n931), .A2(new_n936), .A3(KEYINPUT112), .A4(KEYINPUT54), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n928), .A2(KEYINPUT113), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT113), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n317), .A2(new_n474), .A3(new_n764), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n943), .A2(new_n782), .A3(new_n784), .ZN(new_n944));
  AOI22_X1  g758(.A1(new_n944), .A2(new_n795), .B1(new_n765), .B2(new_n673), .ZN(new_n945));
  AOI22_X1  g759(.A1(new_n692), .A2(new_n765), .B1(new_n777), .B2(new_n778), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n921), .A2(new_n925), .A3(KEYINPUT53), .A4(new_n926), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n941), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n915), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(new_n950), .A3(new_n932), .A4(new_n935), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n930), .A2(new_n933), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT54), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n940), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n890), .A2(new_n939), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(G952), .B2(G953), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n879), .B(KEYINPUT49), .Z(new_n958));
  NOR4_X1   g772(.A1(new_n958), .A2(new_n575), .A3(new_n188), .A4(new_n477), .ZN(new_n959));
  INV_X1    g773(.A(new_n732), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n653), .A2(new_n752), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n959), .A2(new_n859), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n957), .A2(new_n962), .ZN(G75));
  NAND2_X1  g777(.A1(new_n951), .A2(new_n952), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(G902), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT56), .B1(new_n966), .B2(G210), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n259), .A2(new_n261), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(new_n300), .Z(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n321), .A2(G952), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n967), .B2(new_n971), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n972), .A2(new_n975), .ZN(G51));
  NAND2_X1  g790(.A1(new_n964), .A2(KEYINPUT54), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n954), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n479), .B(KEYINPUT57), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n697), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n966), .A2(new_n824), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n973), .B1(new_n981), .B2(new_n982), .ZN(G54));
  NAND3_X1  g797(.A1(new_n966), .A2(KEYINPUT58), .A3(G475), .ZN(new_n984));
  INV_X1    g798(.A(new_n408), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n986), .A2(new_n987), .A3(new_n973), .ZN(G60));
  INV_X1    g802(.A(KEYINPUT120), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n939), .A2(new_n954), .A3(new_n940), .ZN(new_n990));
  NAND2_X1  g804(.A1(G478), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT59), .Z(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n749), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n992), .B1(new_n664), .B2(new_n666), .ZN(new_n995));
  INV_X1    g809(.A(new_n954), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n953), .B1(new_n951), .B2(new_n952), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n974), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n989), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n973), .B1(new_n978), .B2(new_n995), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n992), .B1(new_n955), .B2(new_n939), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n1001), .B(KEYINPUT120), .C1(new_n1002), .C2(new_n749), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1000), .A2(new_n1003), .ZN(G63));
  NAND2_X1  g818(.A1(G217), .A2(G902), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT121), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT60), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n964), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n570), .B(KEYINPUT123), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n973), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT122), .ZN(new_n1011));
  AOI21_X1  g825(.A(KEYINPUT61), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n964), .A2(new_n710), .A3(new_n1007), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1010), .B(new_n1013), .C1(new_n1011), .C2(KEYINPUT61), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(G66));
  OR2_X1    g831(.A1(new_n927), .A2(new_n928), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n321), .ZN(new_n1019));
  OAI21_X1  g833(.A(G953), .B1(new_n472), .B2(new_n298), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n968), .B1(G898), .B2(new_n321), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1021), .B(new_n1022), .ZN(G69));
  XOR2_X1   g837(.A(new_n622), .B(new_n394), .Z(new_n1024));
  AOI21_X1  g838(.A(new_n1024), .B1(G900), .B2(G953), .ZN(new_n1025));
  INV_X1    g839(.A(new_n639), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1026), .A2(new_n895), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n903), .B1(new_n830), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n809), .A2(new_n812), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT124), .Z(new_n1030));
  NAND4_X1  g844(.A1(new_n850), .A2(new_n1028), .A3(new_n1030), .A4(new_n839), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1025), .B1(new_n1031), .B2(G953), .ZN(new_n1032));
  OAI21_X1  g846(.A(KEYINPUT62), .B1(new_n747), .B2(new_n903), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n747), .A2(new_n903), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT62), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n743), .B1(new_n922), .B2(new_n672), .ZN(new_n1036));
  AOI22_X1  g850(.A1(new_n1034), .A2(new_n1035), .B1(new_n811), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n850), .A2(new_n839), .A3(new_n1033), .A4(new_n1037), .ZN(new_n1038));
  AND2_X1   g852(.A1(new_n1038), .A2(new_n321), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1024), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1032), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n321), .B1(G227), .B2(G900), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n1041), .B(new_n1042), .ZN(G72));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT63), .Z(new_n1045));
  OAI21_X1  g859(.A(new_n1045), .B1(new_n1038), .B2(new_n1018), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(KEYINPUT125), .ZN(new_n1047));
  INV_X1    g861(.A(KEYINPUT125), .ZN(new_n1048));
  OAI211_X1 g862(.A(new_n1048), .B(new_n1045), .C1(new_n1038), .C2(new_n1018), .ZN(new_n1049));
  AND3_X1   g863(.A1(new_n1047), .A2(new_n733), .A3(new_n1049), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1045), .B1(new_n1031), .B2(new_n1018), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1051), .A2(new_n623), .A3(new_n580), .ZN(new_n1052));
  AND2_X1   g866(.A1(new_n931), .A2(new_n936), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n734), .A2(new_n630), .A3(new_n1045), .ZN(new_n1054));
  XNOR2_X1  g868(.A(new_n1054), .B(KEYINPUT126), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n973), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g871(.A(KEYINPUT127), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n1047), .A2(new_n733), .A3(new_n1049), .ZN(new_n1059));
  INV_X1    g873(.A(KEYINPUT127), .ZN(new_n1060));
  NAND4_X1  g874(.A1(new_n1059), .A2(new_n1060), .A3(new_n1052), .A4(new_n1056), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1058), .A2(new_n1061), .ZN(G57));
endmodule


