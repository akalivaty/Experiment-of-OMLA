

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586;

  INV_X1 U320 ( .A(KEYINPUT48), .ZN(n371) );
  XNOR2_X1 U321 ( .A(n371), .B(KEYINPUT64), .ZN(n372) );
  XNOR2_X1 U322 ( .A(n373), .B(n372), .ZN(n526) );
  XNOR2_X1 U323 ( .A(n356), .B(n355), .ZN(n357) );
  INV_X1 U324 ( .A(KEYINPUT121), .ZN(n452) );
  XNOR2_X1 U325 ( .A(n358), .B(n357), .ZN(n361) );
  XNOR2_X1 U326 ( .A(n453), .B(n452), .ZN(n583) );
  XNOR2_X1 U327 ( .A(n336), .B(n335), .ZN(n573) );
  XNOR2_X1 U328 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U329 ( .A(n457), .B(n456), .ZN(G1353GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n289) );
  XNOR2_X1 U331 ( .A(KEYINPUT15), .B(KEYINPUT76), .ZN(n288) );
  XNOR2_X1 U332 ( .A(n289), .B(n288), .ZN(n305) );
  XOR2_X1 U333 ( .A(KEYINPUT77), .B(G78GAT), .Z(n291) );
  XNOR2_X1 U334 ( .A(G71GAT), .B(G155GAT), .ZN(n290) );
  XNOR2_X1 U335 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U336 ( .A(G57GAT), .B(KEYINPUT13), .Z(n359) );
  XOR2_X1 U337 ( .A(n292), .B(n359), .Z(n294) );
  XNOR2_X1 U338 ( .A(G127GAT), .B(G211GAT), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U340 ( .A(KEYINPUT14), .B(G64GAT), .Z(n296) );
  NAND2_X1 U341 ( .A1(G231GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U343 ( .A(n298), .B(n297), .Z(n303) );
  XOR2_X1 U344 ( .A(G15GAT), .B(G22GAT), .Z(n300) );
  XNOR2_X1 U345 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U347 ( .A(G1GAT), .B(n301), .Z(n327) );
  XOR2_X1 U348 ( .A(G8GAT), .B(G183GAT), .Z(n374) );
  XNOR2_X1 U349 ( .A(n327), .B(n374), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U351 ( .A(n305), .B(n304), .Z(n563) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(KEYINPUT70), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n306), .B(G29GAT), .ZN(n307) );
  XOR2_X1 U354 ( .A(n307), .B(KEYINPUT7), .Z(n309) );
  XNOR2_X1 U355 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n328) );
  XOR2_X1 U357 ( .A(G99GAT), .B(G85GAT), .Z(n344) );
  XOR2_X1 U358 ( .A(G36GAT), .B(G190GAT), .Z(n388) );
  XNOR2_X1 U359 ( .A(n344), .B(n388), .ZN(n311) );
  AND2_X1 U360 ( .A1(G232GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U362 ( .A(G92GAT), .B(KEYINPUT11), .Z(n313) );
  XNOR2_X1 U363 ( .A(G134GAT), .B(G106GAT), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U365 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U366 ( .A(G50GAT), .B(G162GAT), .Z(n437) );
  XOR2_X1 U367 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n317) );
  XNOR2_X1 U368 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n437), .B(n318), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n328), .B(n321), .ZN(n567) );
  XNOR2_X1 U373 ( .A(KEYINPUT36), .B(n567), .ZN(n584) );
  NOR2_X1 U374 ( .A1(n563), .A2(n584), .ZN(n322) );
  XNOR2_X1 U375 ( .A(KEYINPUT45), .B(n322), .ZN(n337) );
  XOR2_X1 U376 ( .A(G113GAT), .B(G197GAT), .Z(n324) );
  XNOR2_X1 U377 ( .A(G169GAT), .B(G141GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n326) );
  XOR2_X1 U379 ( .A(G50GAT), .B(G36GAT), .Z(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n334) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U382 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n330) );
  XNOR2_X1 U383 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n336) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n335) );
  NAND2_X1 U388 ( .A1(n337), .A2(n573), .ZN(n362) );
  INV_X1 U389 ( .A(G92GAT), .ZN(n338) );
  NAND2_X1 U390 ( .A1(G64GAT), .A2(n338), .ZN(n341) );
  INV_X1 U391 ( .A(G64GAT), .ZN(n339) );
  NAND2_X1 U392 ( .A1(n339), .A2(G92GAT), .ZN(n340) );
  NAND2_X1 U393 ( .A1(n341), .A2(n340), .ZN(n343) );
  XNOR2_X1 U394 ( .A(G176GAT), .B(G204GAT), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n376) );
  XNOR2_X1 U396 ( .A(n376), .B(n344), .ZN(n346) );
  AND2_X1 U397 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n349) );
  INV_X1 U399 ( .A(n349), .ZN(n347) );
  NAND2_X1 U400 ( .A1(n347), .A2(KEYINPUT32), .ZN(n351) );
  INV_X1 U401 ( .A(KEYINPUT32), .ZN(n348) );
  NAND2_X1 U402 ( .A1(n349), .A2(n348), .ZN(n350) );
  NAND2_X1 U403 ( .A1(n351), .A2(n350), .ZN(n358) );
  XNOR2_X1 U404 ( .A(G106GAT), .B(G78GAT), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n352), .B(G148GAT), .ZN(n436) );
  XNOR2_X1 U406 ( .A(n436), .B(KEYINPUT31), .ZN(n356) );
  XOR2_X1 U407 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n354) );
  XNOR2_X1 U408 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n353) );
  XOR2_X1 U409 ( .A(n354), .B(n353), .Z(n355) );
  XOR2_X1 U410 ( .A(G120GAT), .B(G71GAT), .Z(n425) );
  XNOR2_X1 U411 ( .A(n425), .B(n359), .ZN(n360) );
  XNOR2_X1 U412 ( .A(n361), .B(n360), .ZN(n458) );
  NOR2_X1 U413 ( .A1(n362), .A2(n458), .ZN(n363) );
  XNOR2_X1 U414 ( .A(KEYINPUT111), .B(n363), .ZN(n370) );
  INV_X1 U415 ( .A(n563), .ZN(n579) );
  XNOR2_X1 U416 ( .A(n458), .B(KEYINPUT41), .ZN(n546) );
  NOR2_X1 U417 ( .A1(n546), .A2(n573), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n364), .B(KEYINPUT46), .ZN(n365) );
  NOR2_X1 U419 ( .A1(n579), .A2(n365), .ZN(n366) );
  NAND2_X1 U420 ( .A1(n366), .A2(n567), .ZN(n368) );
  XOR2_X1 U421 ( .A(KEYINPUT110), .B(KEYINPUT47), .Z(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n369) );
  NAND2_X1 U423 ( .A1(n370), .A2(n369), .ZN(n373) );
  XNOR2_X1 U424 ( .A(n374), .B(KEYINPUT95), .ZN(n375) );
  XNOR2_X1 U425 ( .A(n375), .B(KEYINPUT96), .ZN(n377) );
  XOR2_X1 U426 ( .A(n377), .B(n376), .Z(n386) );
  XOR2_X1 U427 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n379) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n378) );
  XNOR2_X1 U429 ( .A(n379), .B(n378), .ZN(n429) );
  XOR2_X1 U430 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n381) );
  XNOR2_X1 U431 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n380) );
  XNOR2_X1 U432 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U433 ( .A(n382), .B(KEYINPUT86), .Z(n384) );
  XNOR2_X1 U434 ( .A(G197GAT), .B(G211GAT), .ZN(n383) );
  XNOR2_X1 U435 ( .A(n384), .B(n383), .ZN(n448) );
  XNOR2_X1 U436 ( .A(n429), .B(n448), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U438 ( .A(n388), .B(n387), .Z(n390) );
  NAND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U440 ( .A(n390), .B(n389), .ZN(n504) );
  XNOR2_X1 U441 ( .A(n504), .B(KEYINPUT117), .ZN(n391) );
  NOR2_X1 U442 ( .A1(n526), .A2(n391), .ZN(n392) );
  XNOR2_X1 U443 ( .A(n392), .B(KEYINPUT54), .ZN(n418) );
  XOR2_X1 U444 ( .A(KEYINPUT5), .B(G57GAT), .Z(n394) );
  XNOR2_X1 U445 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U447 ( .A(G148GAT), .B(G162GAT), .Z(n396) );
  XNOR2_X1 U448 ( .A(G1GAT), .B(G120GAT), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n398), .B(n397), .ZN(n410) );
  XOR2_X1 U451 ( .A(KEYINPUT89), .B(KEYINPUT92), .Z(n400) );
  XNOR2_X1 U452 ( .A(KEYINPUT91), .B(KEYINPUT93), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U454 ( .A(KEYINPUT1), .B(KEYINPUT88), .Z(n402) );
  XNOR2_X1 U455 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U458 ( .A(KEYINPUT0), .B(G134GAT), .Z(n406) );
  XNOR2_X1 U459 ( .A(KEYINPUT79), .B(G127GAT), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U461 ( .A(G113GAT), .B(n407), .ZN(n434) );
  XNOR2_X1 U462 ( .A(n408), .B(n434), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(n411), .ZN(n417) );
  XOR2_X1 U465 ( .A(G155GAT), .B(KEYINPUT2), .Z(n413) );
  XNOR2_X1 U466 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n440) );
  XOR2_X1 U468 ( .A(G85GAT), .B(n440), .Z(n415) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n513) );
  NAND2_X1 U472 ( .A1(n418), .A2(n513), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n419), .B(KEYINPUT65), .ZN(n552) );
  XOR2_X1 U474 ( .A(KEYINPUT80), .B(G183GAT), .Z(n421) );
  XNOR2_X1 U475 ( .A(G15GAT), .B(G176GAT), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n433) );
  XOR2_X1 U477 ( .A(KEYINPUT82), .B(G190GAT), .Z(n423) );
  XNOR2_X1 U478 ( .A(G43GAT), .B(G99GAT), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U480 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U481 ( .A1(G227GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U483 ( .A(n428), .B(KEYINPUT81), .Z(n431) );
  XNOR2_X1 U484 ( .A(n429), .B(KEYINPUT20), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n555) );
  XOR2_X1 U488 ( .A(G204GAT), .B(KEYINPUT23), .Z(n439) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n444) );
  XOR2_X1 U491 ( .A(n440), .B(KEYINPUT22), .Z(n442) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U494 ( .A(n444), .B(n443), .Z(n450) );
  XOR2_X1 U495 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n446) );
  XNOR2_X1 U496 ( .A(G22GAT), .B(KEYINPUT83), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U499 ( .A(n450), .B(n449), .ZN(n553) );
  NOR2_X1 U500 ( .A1(n555), .A2(n553), .ZN(n451) );
  XNOR2_X1 U501 ( .A(n451), .B(KEYINPUT26), .ZN(n540) );
  NAND2_X1 U502 ( .A1(n552), .A2(n540), .ZN(n453) );
  INV_X1 U503 ( .A(n583), .ZN(n578) );
  NAND2_X1 U504 ( .A1(n578), .A2(n458), .ZN(n457) );
  XOR2_X1 U505 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n455) );
  INV_X1 U506 ( .A(G204GAT), .ZN(n454) );
  XOR2_X1 U507 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n474) );
  INV_X1 U508 ( .A(n513), .ZN(n487) );
  NOR2_X1 U509 ( .A1(n573), .A2(n458), .ZN(n485) );
  NAND2_X1 U510 ( .A1(n504), .A2(n555), .ZN(n459) );
  NAND2_X1 U511 ( .A1(n553), .A2(n459), .ZN(n460) );
  XOR2_X1 U512 ( .A(KEYINPUT25), .B(n460), .Z(n462) );
  XNOR2_X1 U513 ( .A(n504), .B(KEYINPUT27), .ZN(n464) );
  NAND2_X1 U514 ( .A1(n540), .A2(n464), .ZN(n461) );
  NAND2_X1 U515 ( .A1(n462), .A2(n461), .ZN(n463) );
  NAND2_X1 U516 ( .A1(n463), .A2(n513), .ZN(n468) );
  NAND2_X1 U517 ( .A1(n487), .A2(n464), .ZN(n525) );
  NOR2_X1 U518 ( .A1(n555), .A2(n525), .ZN(n466) );
  XOR2_X1 U519 ( .A(n553), .B(KEYINPUT67), .Z(n465) );
  XNOR2_X1 U520 ( .A(KEYINPUT28), .B(n465), .ZN(n528) );
  NAND2_X1 U521 ( .A1(n466), .A2(n528), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n468), .A2(n467), .ZN(n482) );
  NAND2_X1 U523 ( .A1(n567), .A2(n579), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT16), .B(n469), .Z(n470) );
  NAND2_X1 U525 ( .A1(n482), .A2(n470), .ZN(n471) );
  XNOR2_X1 U526 ( .A(n471), .B(KEYINPUT97), .ZN(n500) );
  NAND2_X1 U527 ( .A1(n485), .A2(n500), .ZN(n472) );
  XOR2_X1 U528 ( .A(KEYINPUT98), .B(n472), .Z(n479) );
  NAND2_X1 U529 ( .A1(n487), .A2(n479), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U532 ( .A1(n479), .A2(n504), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U535 ( .A1(n479), .A2(n555), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  XNOR2_X1 U537 ( .A(G22GAT), .B(KEYINPUT100), .ZN(n481) );
  INV_X1 U538 ( .A(n528), .ZN(n496) );
  NAND2_X1 U539 ( .A1(n496), .A2(n479), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(G1327GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n489) );
  NAND2_X1 U542 ( .A1(n563), .A2(n482), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n584), .A2(n483), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT37), .B(n484), .Z(n512) );
  NAND2_X1 U545 ( .A1(n512), .A2(n485), .ZN(n486) );
  XOR2_X1 U546 ( .A(KEYINPUT38), .B(n486), .Z(n495) );
  NAND2_X1 U547 ( .A1(n487), .A2(n495), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U549 ( .A(G29GAT), .B(n490), .Z(G1328GAT) );
  NAND2_X1 U550 ( .A1(n495), .A2(n504), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n491), .B(KEYINPUT102), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  NAND2_X1 U553 ( .A1(n495), .A2(n555), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  XOR2_X1 U556 ( .A(G50GAT), .B(KEYINPUT103), .Z(n498) );
  NAND2_X1 U557 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  INV_X1 U559 ( .A(n573), .ZN(n499) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(n546), .Z(n558) );
  NOR2_X1 U561 ( .A1(n499), .A2(n558), .ZN(n511) );
  NAND2_X1 U562 ( .A1(n500), .A2(n511), .ZN(n508) );
  NOR2_X1 U563 ( .A1(n513), .A2(n508), .ZN(n502) );
  XNOR2_X1 U564 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n503), .Z(G1332GAT) );
  INV_X1 U567 ( .A(n504), .ZN(n516) );
  NOR2_X1 U568 ( .A1(n516), .A2(n508), .ZN(n505) );
  XOR2_X1 U569 ( .A(KEYINPUT106), .B(n505), .Z(n506) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  INV_X1 U571 ( .A(n555), .ZN(n518) );
  NOR2_X1 U572 ( .A1(n518), .A2(n508), .ZN(n507) );
  XOR2_X1 U573 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U574 ( .A1(n528), .A2(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n522) );
  NOR2_X1 U578 ( .A1(n513), .A2(n522), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1336GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n522), .ZN(n517) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n517), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n522), .ZN(n519) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n521) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n524) );
  NOR2_X1 U588 ( .A1(n528), .A2(n522), .ZN(n523) );
  XOR2_X1 U589 ( .A(n524), .B(n523), .Z(G1339GAT) );
  NOR2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n539), .A2(n555), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT112), .B(n527), .Z(n529) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n536) );
  NOR2_X1 U594 ( .A1(n573), .A2(n536), .ZN(n530) );
  XOR2_X1 U595 ( .A(G113GAT), .B(n530), .Z(G1340GAT) );
  NOR2_X1 U596 ( .A1(n558), .A2(n536), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U599 ( .A1(n563), .A2(n536), .ZN(n534) );
  XNOR2_X1 U600 ( .A(KEYINPUT113), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  NOR2_X1 U603 ( .A1(n567), .A2(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n541), .B(KEYINPUT114), .ZN(n550) );
  NOR2_X1 U609 ( .A1(n573), .A2(n550), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n548) );
  NOR2_X1 U614 ( .A1(n550), .A2(n546), .ZN(n547) );
  XOR2_X1 U615 ( .A(n548), .B(n547), .Z(G1345GAT) );
  NOR2_X1 U616 ( .A1(n563), .A2(n550), .ZN(n549) );
  XOR2_X1 U617 ( .A(G155GAT), .B(n549), .Z(G1346GAT) );
  NOR2_X1 U618 ( .A1(n550), .A2(n567), .ZN(n551) );
  XOR2_X1 U619 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT55), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n566) );
  NOR2_X1 U623 ( .A1(n573), .A2(n566), .ZN(n557) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n557), .Z(G1348GAT) );
  XNOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT118), .ZN(n562) );
  NOR2_X1 U626 ( .A1(n566), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NOR2_X1 U630 ( .A1(n563), .A2(n566), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT119), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1350GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n569) );
  XNOR2_X1 U634 ( .A(KEYINPUT120), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(G190GAT), .B(n570), .Z(G1351GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n577) );
  NOR2_X1 U640 ( .A1(n573), .A2(n583), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n582) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n586) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(n586), .B(n585), .Z(G1355GAT) );
endmodule

