//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XOR2_X1   g0002(.A(new_n202), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0003(.A(G1), .ZN(new_n204));
  INV_X1    g0004(.A(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(G58), .A2(G68), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n215), .A2(G50), .A3(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT67), .Z(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT66), .Z(new_n224));
  OAI21_X1  g0024(.A(new_n207), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n210), .B1(new_n213), .B2(new_n217), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT68), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT69), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n232), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT70), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G58), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  XNOR2_X1  g0045(.A(KEYINPUT3), .B(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G222), .A2(G1698), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(G223), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n246), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n212), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n250), .B(new_n253), .C1(G77), .C2(new_n246), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT72), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(KEYINPUT72), .A2(G33), .A3(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(new_n212), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n204), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT71), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n204), .B(KEYINPUT71), .C1(G41), .C2(G45), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n258), .A2(new_n261), .A3(G274), .A4(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n258), .A2(G226), .A3(new_n259), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n254), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G169), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n211), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT8), .B(G58), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n205), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G150), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n270), .A2(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G50), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n205), .B1(new_n214), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n269), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n204), .A2(G13), .A3(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT73), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT73), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n281), .A2(new_n204), .A3(G13), .A4(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n276), .ZN(new_n285));
  INV_X1    g0085(.A(new_n269), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n204), .A2(G20), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n283), .A2(new_n286), .A3(G50), .A4(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n278), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n267), .B(new_n289), .C1(G179), .C2(new_n265), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT9), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n265), .A2(G200), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n278), .A2(new_n285), .A3(KEYINPUT9), .A4(new_n288), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n254), .A2(G190), .A3(new_n263), .A4(new_n264), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n294), .A2(new_n297), .A3(KEYINPUT10), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(new_n297), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n291), .A2(new_n289), .B1(new_n265), .B2(G200), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n290), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n246), .A2(G238), .A3(G1698), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n246), .A2(G232), .A3(new_n248), .ZN(new_n305));
  INV_X1    g0105(.A(G107), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n246), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n253), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n258), .A2(G244), .A3(new_n259), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n263), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(G169), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n310), .B1(new_n253), .B2(new_n307), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n270), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n273), .A2(KEYINPUT75), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n273), .A2(KEYINPUT75), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G20), .A2(G77), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(KEYINPUT76), .A3(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n271), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT76), .B1(new_n319), .B2(new_n320), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n269), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n284), .A2(new_n269), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n204), .B2(G20), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n326), .A2(new_n328), .B1(new_n327), .B2(new_n284), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n315), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n308), .A2(new_n311), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G200), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n333), .A2(KEYINPUT74), .B1(new_n314), .B2(G190), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n308), .A2(new_n311), .A3(KEYINPUT74), .A4(G190), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n325), .A2(new_n335), .A3(new_n329), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n331), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT77), .B1(new_n303), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n333), .A2(KEYINPUT74), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n314), .A2(G190), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n325), .A2(new_n335), .A3(new_n329), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n341), .A2(new_n342), .B1(new_n330), .B2(new_n315), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT10), .B1(new_n294), .B2(new_n297), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n300), .A2(new_n301), .A3(new_n299), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT77), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n343), .A2(new_n346), .A3(new_n347), .A4(new_n290), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n338), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n258), .A2(G238), .A3(new_n259), .ZN(new_n350));
  NOR2_X1   g0150(.A1(G226), .A2(G1698), .ZN(new_n351));
  INV_X1    g0151(.A(G232), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(G1698), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n246), .B1(G33), .B2(G97), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n263), .B(new_n350), .C1(new_n354), .C2(new_n252), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT13), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G97), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n352), .A2(G1698), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G226), .B2(G1698), .ZN(new_n359));
  INV_X1    g0159(.A(G33), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT3), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G33), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n357), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n253), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n350), .A4(new_n263), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n356), .A2(KEYINPUT78), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT78), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n355), .A2(new_n370), .A3(KEYINPUT13), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(G169), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT14), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n369), .A2(new_n374), .A3(G169), .A4(new_n371), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n356), .A2(G179), .A3(new_n368), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT80), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT80), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n356), .A2(new_n378), .A3(G179), .A4(new_n368), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n373), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT79), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n283), .A2(new_n286), .A3(G68), .A4(new_n287), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n273), .A2(G50), .ZN(new_n384));
  INV_X1    g0184(.A(G68), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G20), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n384), .B(new_n386), .C1(new_n327), .C2(new_n271), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n269), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(KEYINPUT11), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT11), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n387), .B2(new_n269), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n383), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n280), .A2(new_n385), .A3(new_n282), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n393), .B(KEYINPUT12), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n382), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n388), .B(KEYINPUT11), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n397), .A2(KEYINPUT79), .A3(new_n394), .A4(new_n383), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n381), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n369), .A2(G200), .A3(new_n371), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n356), .A2(G190), .A3(new_n368), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G58), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(new_n385), .ZN(new_n407));
  OAI21_X1  g0207(.A(G20), .B1(new_n407), .B2(new_n214), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n273), .A2(G159), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT81), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n362), .B2(G33), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n360), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n363), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT7), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(new_n205), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G68), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n415), .B2(new_n205), .ZN(new_n419));
  OAI211_X1 g0219(.A(KEYINPUT16), .B(new_n411), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT82), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n413), .A2(new_n363), .A3(new_n414), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT7), .B1(new_n422), .B2(G20), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(G68), .A3(new_n417), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT82), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT16), .A4(new_n411), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT83), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT7), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n416), .A2(KEYINPUT83), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n246), .B2(G20), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n364), .A2(new_n205), .A3(new_n430), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n410), .B1(new_n434), .B2(G68), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n269), .B1(new_n435), .B2(KEYINPUT16), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n427), .A2(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(G223), .A2(G1698), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(G226), .B2(new_n248), .ZN(new_n440));
  INV_X1    g0240(.A(G87), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n415), .A2(new_n440), .B1(new_n360), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n253), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n258), .A2(G232), .A3(new_n259), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n263), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G190), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n447), .B1(G200), .B2(new_n445), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n270), .B1(new_n204), .B2(G20), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n326), .A2(new_n449), .B1(new_n284), .B2(new_n270), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n438), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n445), .A2(G169), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n313), .B2(new_n445), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n436), .B1(new_n421), .B2(new_n426), .ZN(new_n456));
  INV_X1    g0256(.A(new_n450), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT18), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT18), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n455), .C1(new_n456), .C2(new_n457), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n427), .B2(new_n437), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(KEYINPUT17), .A3(new_n448), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n453), .A2(new_n459), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n349), .A2(new_n405), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n204), .A2(G45), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n466), .A2(G250), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n258), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT85), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT85), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n258), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G274), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n211), .B1(new_n255), .B2(new_n251), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(new_n257), .ZN(new_n475));
  INV_X1    g0275(.A(new_n466), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n414), .A2(new_n363), .ZN(new_n480));
  INV_X1    g0280(.A(G238), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G1698), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n480), .A2(KEYINPUT86), .A3(new_n413), .A4(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n413), .A2(new_n414), .A3(new_n482), .A4(new_n363), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT86), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G116), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n413), .A2(new_n414), .A3(G244), .A4(new_n363), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n248), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT87), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n253), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n487), .B2(new_n491), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n313), .B(new_n479), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT88), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n479), .B1(new_n494), .B2(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n266), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n487), .A2(new_n491), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT87), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(new_n253), .A3(new_n493), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(KEYINPUT88), .A3(new_n313), .A4(new_n479), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n422), .A2(new_n205), .A3(G68), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n360), .A2(G20), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT19), .B1(new_n506), .B2(G97), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT19), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n205), .B1(new_n357), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G97), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n441), .A2(new_n510), .A3(new_n306), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n269), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n284), .A2(new_n322), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n360), .A2(G1), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n516), .B(new_n269), .C1(new_n280), .C2(new_n282), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n514), .B(new_n515), .C1(new_n322), .C2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n498), .A2(new_n500), .A3(new_n504), .A4(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G190), .B(new_n479), .C1(new_n494), .C2(new_n495), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(G87), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n514), .A2(new_n522), .A3(new_n515), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n490), .B1(new_n486), .B2(new_n483), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n252), .B1(new_n524), .B2(new_n492), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n478), .B1(new_n525), .B2(new_n502), .ZN(new_n526));
  INV_X1    g0326(.A(G200), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n521), .B(new_n523), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n306), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  XOR2_X1   g0330(.A(G97), .B(G107), .Z(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G20), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n327), .B2(new_n274), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n434), .A2(G107), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n269), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n284), .A2(new_n510), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n517), .A2(G97), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n246), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n246), .A2(G250), .A3(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT4), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n489), .B2(G1698), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n252), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G41), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n204), .B(G45), .C1(new_n548), .C2(KEYINPUT5), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT84), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(KEYINPUT5), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n549), .B2(KEYINPUT84), .ZN(new_n553));
  OAI211_X1 g0353(.A(G257), .B(new_n258), .C1(new_n551), .C2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT84), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n476), .B(new_n555), .C1(KEYINPUT5), .C2(new_n548), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n475), .A2(new_n556), .A3(new_n550), .A4(new_n552), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n313), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n266), .B1(new_n547), .B2(new_n558), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n540), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n539), .A2(new_n538), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n535), .B(new_n533), .C1(new_n327), .C2(new_n274), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(new_n269), .ZN(new_n565));
  OAI21_X1  g0365(.A(G200), .B1(new_n547), .B2(new_n558), .ZN(new_n566));
  INV_X1    g0366(.A(new_n558), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n544), .A2(new_n546), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n568), .B2(new_n252), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n565), .B(new_n566), .C1(new_n569), .C2(new_n446), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n306), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT25), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n283), .B2(G107), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n571), .A2(new_n573), .B1(new_n517), .B2(G107), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT91), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n205), .A2(G87), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n364), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n205), .B2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n306), .A2(KEYINPUT23), .A3(G20), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n580), .A2(new_n581), .B1(new_n506), .B2(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n576), .A2(new_n441), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n415), .A2(G20), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT24), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n422), .A2(new_n205), .A3(new_n584), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT24), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(new_n578), .A4(new_n582), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n575), .B1(new_n591), .B2(new_n269), .ZN(new_n592));
  AOI211_X1 g0392(.A(KEYINPUT91), .B(new_n286), .C1(new_n587), .C2(new_n590), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n574), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(G264), .B(new_n258), .C1(new_n551), .C2(new_n553), .ZN(new_n595));
  OR2_X1    g0395(.A1(G250), .A2(G1698), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G257), .B2(new_n248), .ZN(new_n597));
  INV_X1    g0397(.A(G294), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n415), .A2(new_n597), .B1(new_n360), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n253), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n595), .B(new_n557), .C1(new_n600), .C2(KEYINPUT92), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n600), .A2(KEYINPUT92), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n595), .A3(new_n557), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n603), .A2(new_n446), .B1(new_n527), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n562), .B(new_n570), .C1(new_n594), .C2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n516), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n283), .A2(new_n286), .A3(G116), .A4(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n280), .A2(new_n610), .A3(new_n282), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(G20), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n269), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT89), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n269), .A2(KEYINPUT89), .A3(new_n614), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n543), .B(new_n205), .C1(G33), .C2(new_n510), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT20), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n269), .A2(KEYINPUT89), .A3(new_n614), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT89), .B1(new_n269), .B2(new_n614), .ZN(new_n623));
  OAI211_X1 g0423(.A(KEYINPUT20), .B(new_n620), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n613), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  OR2_X1    g0426(.A1(G257), .A2(G1698), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(G264), .B2(new_n248), .ZN(new_n628));
  INV_X1    g0428(.A(G303), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n415), .A2(new_n628), .B1(new_n629), .B2(new_n246), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n253), .ZN(new_n631));
  OAI211_X1 g0431(.A(G270), .B(new_n258), .C1(new_n551), .C2(new_n553), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n632), .A3(new_n557), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n626), .A2(KEYINPUT21), .A3(G169), .A4(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(G169), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT20), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n612), .B1(new_n639), .B2(new_n624), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n635), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n633), .A2(new_n313), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n626), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n634), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n603), .A2(new_n266), .B1(new_n313), .B2(new_n604), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n594), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n633), .A2(G200), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n640), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT90), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n648), .A2(new_n640), .A3(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n650), .B(new_n652), .C1(new_n446), .C2(new_n633), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n645), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n465), .A2(new_n529), .A3(new_n607), .A4(new_n654), .ZN(G372));
  INV_X1    g0455(.A(new_n562), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n520), .A2(KEYINPUT26), .A3(new_n528), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n521), .A2(new_n523), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT93), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n526), .B2(new_n527), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n499), .A2(KEYINPUT93), .A3(G200), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n496), .B(new_n519), .C1(new_n526), .C2(G169), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n662), .A2(new_n664), .A3(new_n562), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n657), .B1(new_n665), .B2(KEYINPUT26), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n644), .B1(new_n594), .B2(new_n646), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n606), .ZN(new_n668));
  INV_X1    g0468(.A(new_n658), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n526), .A2(new_n659), .A3(new_n527), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT93), .B1(new_n499), .B2(G200), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n664), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n465), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT94), .ZN(new_n677));
  INV_X1    g0477(.A(new_n290), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n459), .A2(new_n461), .ZN(new_n679));
  INV_X1    g0479(.A(new_n331), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n381), .A2(new_n400), .B1(new_n680), .B2(new_n404), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n453), .A2(new_n463), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n678), .B1(new_n683), .B2(new_n346), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n677), .A2(new_n684), .ZN(G369));
  NAND3_X1  g0485(.A1(new_n204), .A2(new_n205), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n626), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n645), .A2(new_n653), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n645), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n594), .A2(new_n691), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n647), .B(new_n697), .C1(new_n594), .C2(new_n605), .ZN(new_n698));
  INV_X1    g0498(.A(new_n691), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n647), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n594), .A2(new_n646), .A3(new_n699), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n644), .A2(new_n699), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n208), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n511), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n217), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n529), .A2(new_n654), .A3(new_n607), .A4(new_n699), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n633), .A2(new_n313), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT96), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n569), .B2(new_n604), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n715), .B(new_n604), .C1(new_n547), .C2(new_n558), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n499), .B(new_n714), .C1(new_n716), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n559), .A2(new_n642), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n600), .A2(new_n595), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n479), .B(new_n721), .C1(new_n494), .C2(new_n495), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT95), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n503), .A2(KEYINPUT95), .A3(new_n479), .A4(new_n721), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n720), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n719), .B1(new_n726), .B2(KEYINPUT30), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  AOI211_X1 g0528(.A(new_n728), .B(new_n720), .C1(new_n724), .C2(new_n725), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n691), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n713), .A2(new_n730), .A3(KEYINPUT31), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n691), .C1(new_n727), .C2(new_n729), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n520), .A2(new_n528), .A3(new_n656), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT26), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n672), .A2(KEYINPUT26), .A3(new_n656), .A4(new_n663), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n645), .A2(new_n647), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n607), .A2(new_n672), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n663), .ZN(new_n743));
  OAI211_X1 g0543(.A(KEYINPUT29), .B(new_n699), .C1(new_n740), .C2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n691), .B1(new_n666), .B2(new_n673), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(KEYINPUT29), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n735), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n712), .B1(new_n747), .B2(G1), .ZN(G364));
  INV_X1    g0548(.A(G13), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n204), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n707), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n696), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G330), .B2(new_n694), .ZN(new_n755));
  INV_X1    g0555(.A(new_n753), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n211), .B1(G20), .B2(new_n266), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n205), .A2(new_n313), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n760), .A2(new_n527), .A3(G190), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n760), .A2(new_n446), .A3(new_n527), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n762), .A2(new_n385), .B1(new_n764), .B2(new_n276), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G190), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n765), .B1(G77), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n205), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n446), .A3(G200), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT97), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G107), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n446), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n205), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n510), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n770), .A2(new_n766), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n777), .A2(KEYINPUT32), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n441), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n776), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT32), .ZN(new_n783));
  INV_X1    g0583(.A(new_n777), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(new_n784), .B2(G159), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n760), .A2(new_n446), .A3(G200), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n364), .B(new_n785), .C1(G58), .C2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n769), .A2(new_n773), .A3(new_n782), .A4(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n364), .B1(new_n767), .B2(new_n789), .C1(new_n775), .C2(new_n598), .ZN(new_n790));
  INV_X1    g0590(.A(new_n780), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(G303), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n772), .A2(G283), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G326), .A2(new_n763), .B1(new_n761), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n786), .A2(G322), .B1(G329), .B2(new_n784), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n792), .A2(new_n793), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n758), .B1(new_n788), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n757), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n706), .A2(new_n364), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n803), .A2(G355), .B1(new_n610), .B2(new_n706), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n706), .A2(new_n422), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(G45), .B2(new_n217), .ZN(new_n806));
  INV_X1    g0606(.A(G45), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n244), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n804), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n756), .B(new_n798), .C1(new_n802), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n801), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n694), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n755), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  AOI22_X1  g0614(.A1(new_n341), .A2(new_n342), .B1(new_n330), .B2(new_n691), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(new_n680), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n680), .A2(new_n699), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n691), .B(new_n818), .C1(new_n666), .C2(new_n673), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(KEYINPUT99), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n818), .B1(new_n674), .B2(new_n691), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n820), .B(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n753), .B1(new_n822), .B2(new_n735), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n735), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n757), .A2(new_n799), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n753), .B1(G77), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  INV_X1    g0628(.A(new_n786), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n828), .A2(new_n762), .B1(new_n829), .B2(new_n598), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n764), .A2(new_n629), .B1(new_n777), .B2(new_n789), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n246), .B(new_n776), .C1(G116), .C2(new_n768), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n772), .A2(G87), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n791), .A2(G107), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n786), .A2(G143), .B1(new_n763), .B2(G137), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n272), .B2(new_n762), .C1(new_n778), .C2(new_n767), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT34), .Z(new_n839));
  NAND2_X1  g0639(.A1(new_n772), .A2(G68), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n415), .B1(new_n784), .B2(G132), .ZN(new_n841));
  INV_X1    g0641(.A(new_n775), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n842), .A2(G58), .B1(new_n791), .B2(G50), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n836), .B1(new_n839), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n827), .B1(new_n845), .B2(new_n757), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT98), .Z(new_n847));
  INV_X1    g0647(.A(new_n818), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(new_n800), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n824), .A2(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n750), .A2(new_n204), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n689), .B(KEYINPUT102), .Z(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n456), .B2(new_n457), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n464), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n451), .A2(new_n458), .A3(new_n854), .ZN(new_n857));
  XOR2_X1   g0657(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n451), .A2(new_n458), .A3(new_n854), .A4(new_n858), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n852), .B1(new_n856), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n424), .A2(new_n411), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT16), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n286), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n427), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n450), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n455), .ZN(new_n869));
  INV_X1    g0669(.A(new_n689), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n871), .A3(new_n451), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n861), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n464), .A2(new_n870), .A3(new_n868), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n863), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n381), .A2(new_n400), .A3(new_n699), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT104), .Z(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n464), .A2(new_n870), .A3(new_n868), .ZN(new_n883));
  INV_X1    g0683(.A(new_n861), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(KEYINPUT37), .B2(new_n872), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n852), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(KEYINPUT39), .A3(new_n876), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n879), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n876), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n404), .A2(new_n373), .A3(new_n375), .A4(new_n380), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n399), .A2(new_n699), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT101), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n401), .B(new_n404), .C1(new_n399), .C2(new_n699), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n890), .B2(new_n891), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n817), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n889), .B(new_n896), .C1(new_n819), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n679), .A2(new_n853), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n888), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT105), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n888), .A2(new_n898), .A3(new_n903), .A4(new_n900), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n744), .B(new_n465), .C1(KEYINPUT29), .C2(new_n745), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n684), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n905), .B(new_n907), .Z(new_n908));
  INV_X1    g0708(.A(G330), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n875), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n874), .B2(new_n875), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n731), .A2(new_n896), .A3(new_n733), .A4(new_n848), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n896), .A2(new_n848), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n734), .A2(new_n877), .A3(new_n916), .A4(KEYINPUT40), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n734), .A2(new_n465), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n909), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n918), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n851), .B1(new_n908), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n921), .B2(new_n908), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n610), .B(new_n213), .C1(new_n532), .C2(KEYINPUT35), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(KEYINPUT35), .B2(new_n532), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT36), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n217), .A2(new_n327), .A3(new_n407), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n276), .B2(G68), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n749), .A2(G1), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT100), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n923), .A2(new_n931), .ZN(G367));
  INV_X1    g0732(.A(new_n805), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n236), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n802), .B1(new_n208), .B2(new_n322), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n753), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n764), .A2(new_n789), .B1(new_n767), .B2(new_n828), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(G294), .B2(new_n761), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n791), .A2(G116), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT46), .ZN(new_n940));
  INV_X1    g0740(.A(G317), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n777), .A2(new_n941), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n422), .B(new_n942), .C1(new_n786), .C2(G303), .ZN(new_n943));
  INV_X1    g0743(.A(new_n771), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n842), .A2(G107), .B1(new_n944), .B2(G97), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n938), .A2(new_n940), .A3(new_n943), .A4(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(G143), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n762), .A2(new_n778), .B1(new_n764), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(KEYINPUT110), .B(G137), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n948), .B1(new_n784), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n246), .B1(new_n767), .B2(new_n276), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(G58), .B2(new_n791), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n951), .B(new_n953), .C1(new_n327), .C2(new_n771), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n775), .A2(new_n385), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G150), .B2(new_n786), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT109), .Z(new_n957));
  OAI21_X1  g0757(.A(new_n946), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT47), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n936), .B1(new_n959), .B2(new_n757), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n672), .B(new_n663), .C1(new_n523), .C2(new_n699), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n663), .A2(new_n523), .A3(new_n699), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n960), .B1(new_n963), .B2(new_n811), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n704), .A2(new_n702), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n656), .A2(new_n691), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n562), .B(new_n570), .C1(new_n565), .C2(new_n699), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n969));
  OR3_X1    g0769(.A1(new_n965), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n965), .B2(new_n968), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT108), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT44), .B1(new_n965), .B2(new_n968), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n970), .A2(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n972), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n965), .A2(KEYINPUT44), .A3(new_n968), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(new_n701), .ZN(new_n979));
  INV_X1    g0779(.A(new_n703), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n704), .B1(new_n700), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(new_n695), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n747), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n747), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n707), .B(KEYINPUT41), .Z(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n752), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n704), .A2(new_n968), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT42), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n562), .B1(new_n967), .B2(new_n647), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n699), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT43), .B1(new_n963), .B2(KEYINPUT106), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(KEYINPUT106), .B2(new_n963), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n995), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n997), .B2(new_n995), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n701), .A2(new_n968), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1000), .B(new_n1001), .Z(new_n1002));
  OAI21_X1  g0802(.A(new_n964), .B1(new_n990), .B2(new_n1002), .ZN(G387));
  NAND2_X1  g0803(.A1(new_n232), .A2(G45), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n807), .B1(new_n385), .B2(new_n327), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n709), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT111), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n316), .A2(KEYINPUT50), .A3(new_n276), .ZN(new_n1009));
  AOI21_X1  g0809(.A(KEYINPUT50), .B1(new_n316), .B2(new_n276), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1008), .B1(new_n1007), .B2(new_n1006), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1004), .A2(new_n805), .A3(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n803), .A2(new_n1006), .B1(new_n306), .B2(new_n706), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n801), .B(new_n757), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n422), .B1(G326), .B2(new_n784), .ZN(new_n1015));
  INV_X1    g0815(.A(G322), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n829), .A2(new_n941), .B1(new_n764), .B2(new_n1016), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n762), .A2(new_n789), .B1(new_n767), .B2(new_n629), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n842), .A2(G283), .B1(new_n791), .B2(G294), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1019), .A2(KEYINPUT48), .B1(KEYINPUT113), .B2(new_n1020), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1020), .A2(KEYINPUT113), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(KEYINPUT48), .C2(new_n1019), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT49), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1015), .B1(new_n610), .B2(new_n771), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n780), .A2(new_n327), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n415), .B(new_n1027), .C1(G150), .C2(new_n784), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n772), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n510), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT112), .Z(new_n1031));
  AOI22_X1  g0831(.A1(new_n316), .A2(new_n761), .B1(new_n786), .B2(G50), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n763), .A2(G159), .B1(G68), .B2(new_n768), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n322), .C2(new_n775), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n1025), .A2(new_n1026), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT114), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n758), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n756), .B(new_n1014), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n700), .A2(new_n811), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n983), .A2(new_n752), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n984), .A2(KEYINPUT115), .A3(new_n707), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n747), .B2(new_n983), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT115), .B1(new_n984), .B2(new_n707), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(G393));
  AOI21_X1  g0845(.A(new_n708), .B1(new_n979), .B2(new_n985), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n985), .B2(new_n979), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n979), .A2(new_n752), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n802), .B1(new_n510), .B2(new_n208), .C1(new_n241), .C2(new_n933), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT116), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n756), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n761), .A2(G303), .B1(G294), .B2(new_n768), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n610), .B2(new_n775), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT118), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n786), .A2(G311), .B1(new_n763), .B2(G317), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  OAI21_X1  g0857(.A(new_n364), .B1(new_n777), .B2(new_n1016), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G283), .B2(new_n791), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1055), .A2(new_n773), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n786), .A2(G159), .B1(new_n763), .B2(G150), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT51), .Z(new_n1062));
  NOR2_X1   g0862(.A1(new_n775), .A2(new_n327), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n422), .B1(new_n947), .B2(new_n777), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(G68), .C2(new_n791), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n761), .A2(G50), .B1(new_n316), .B2(new_n768), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT117), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1062), .A2(new_n834), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n758), .B1(new_n1060), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1052), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n968), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n811), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1047), .A2(new_n1048), .A3(new_n1072), .ZN(G390));
  NAND2_X1  g0873(.A1(new_n879), .A2(new_n887), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n799), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n306), .A2(new_n762), .B1(new_n829), .B2(new_n610), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n764), .A2(new_n828), .B1(new_n777), .B2(new_n598), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1063), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n246), .B(new_n781), .C1(G97), .C2(new_n768), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1078), .A2(new_n840), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n780), .A2(new_n272), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT53), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(KEYINPUT54), .B(G143), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n364), .B1(new_n768), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n762), .A2(new_n949), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G125), .B2(new_n784), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n842), .A2(G159), .B1(new_n944), .B2(G50), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1083), .A2(new_n1086), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n786), .A2(G132), .B1(new_n763), .B2(G128), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT121), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1081), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT122), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n758), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n756), .B1(new_n270), .B2(new_n825), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1075), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n731), .A2(G330), .A3(new_n733), .A4(new_n848), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n896), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n896), .B1(new_n819), .B2(new_n897), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1102), .A2(new_n881), .B1(new_n879), .B2(new_n887), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n877), .A2(new_n881), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n738), .A2(new_n739), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n691), .B1(new_n673), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n897), .B1(new_n1106), .B2(new_n816), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1104), .B1(new_n1108), .B2(new_n896), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1101), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n745), .A2(new_n848), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1100), .B1(new_n1111), .B2(new_n817), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1074), .B1(new_n1112), .B2(new_n882), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n877), .B(new_n881), .C1(new_n1107), .C2(new_n1100), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1098), .B1(new_n1117), .B2(new_n751), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1119), .A2(new_n1101), .B1(new_n897), .B2(new_n819), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1114), .A2(new_n1107), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NOR4_X1   g0923(.A1(new_n349), .A2(new_n405), .A3(new_n464), .A4(new_n909), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1124), .A2(new_n731), .A3(new_n733), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT119), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT120), .B1(new_n1127), .B2(new_n907), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n734), .A2(new_n1126), .A3(new_n1124), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1125), .A2(KEYINPUT119), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT120), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1131), .A2(new_n1132), .A3(new_n684), .A4(new_n906), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1123), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n708), .B1(new_n1117), .B2(new_n1134), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1118), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(G378));
  AND2_X1   g0940(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1117), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n915), .A2(G330), .A3(new_n917), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n303), .B(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n289), .A2(new_n870), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT123), .Z(new_n1148));
  XNOR2_X1  g0948(.A(new_n1146), .B(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1144), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n915), .A2(G330), .A3(new_n917), .A4(new_n1149), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n902), .A2(new_n1151), .A3(new_n904), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n905), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1143), .A2(KEYINPUT57), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n707), .ZN(new_n1157));
  AND4_X1   g0957(.A1(new_n904), .A2(new_n902), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n904), .A2(new_n902), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT57), .B1(new_n1160), .B2(new_n1143), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1155), .A2(new_n752), .A3(new_n1153), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n756), .B1(new_n276), .B2(new_n825), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n761), .A2(G132), .B1(new_n763), .B2(G125), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n786), .A2(G128), .B1(G137), .B2(new_n768), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n842), .A2(G150), .B1(new_n791), .B2(new_n1085), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n944), .A2(G159), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n784), .C2(G124), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n829), .A2(new_n306), .B1(new_n777), .B2(new_n828), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n771), .A2(new_n406), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(new_n1174), .A2(new_n955), .A3(new_n1027), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n761), .A2(G97), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n322), .B2(new_n767), .C1(new_n764), .C2(new_n610), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n548), .A3(new_n415), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1183));
  AOI21_X1  g0983(.A(G50), .B1(new_n360), .B2(new_n548), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n422), .B2(G41), .ZN(new_n1185));
  AND4_X1   g0985(.A1(new_n1173), .A2(new_n1182), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1164), .B1(new_n758), .B2(new_n1186), .C1(new_n1149), .C2(new_n800), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1163), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1162), .A2(new_n1189), .ZN(G375));
  OAI22_X1  g0990(.A1(new_n610), .A2(new_n762), .B1(new_n829), .B2(new_n828), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n764), .A2(new_n598), .B1(new_n777), .B2(new_n629), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n775), .A2(new_n322), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n246), .B(new_n1194), .C1(G107), .C2(new_n768), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n772), .A2(G77), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n791), .A2(G97), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n775), .A2(new_n276), .B1(new_n767), .B2(new_n272), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT124), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n415), .B(new_n1175), .C1(G159), .C2(new_n791), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1085), .A2(new_n761), .B1(new_n763), .B2(G132), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n786), .A2(new_n950), .B1(new_n784), .B2(G128), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1198), .B1(new_n1200), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n758), .B1(new_n1205), .B2(KEYINPUT125), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(KEYINPUT125), .B2(new_n1205), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1207), .B(new_n753), .C1(G68), .C2(new_n826), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1100), .B2(new_n799), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1123), .B2(new_n752), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1134), .A2(new_n989), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1123), .B1(new_n1133), .B2(new_n1128), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(G381));
  OR2_X1    g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  OR4_X1    g1014(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1214), .ZN(new_n1215));
  OR4_X1    g1015(.A1(G378), .A2(new_n1215), .A3(G375), .A4(G381), .ZN(G407));
  AND2_X1   g1016(.A1(new_n690), .A2(G213), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1139), .A2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(G407), .B(G213), .C1(G375), .C2(new_n1218), .ZN(G409));
  NAND2_X1  g1019(.A1(new_n1217), .A2(G2897), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT60), .B1(new_n1221), .B2(new_n1142), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT126), .B1(new_n1222), .B2(new_n1135), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT126), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1224), .B(new_n1134), .C1(new_n1212), .C2(KEYINPUT60), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n708), .B1(new_n1212), .B2(KEYINPUT60), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1210), .ZN(new_n1228));
  INV_X1    g1028(.A(G384), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(G384), .A3(new_n1210), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1220), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G378), .B(new_n1189), .C1(new_n1157), .C2(new_n1161), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1160), .A2(new_n989), .A3(new_n1143), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1139), .B1(new_n1234), .B2(new_n1188), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1217), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1232), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT127), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1227), .A2(G384), .A3(new_n1210), .ZN(new_n1239));
  AOI21_X1  g1039(.A(G384), .B1(new_n1227), .B2(new_n1210), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1230), .A2(KEYINPUT127), .A3(new_n1231), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n1220), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1237), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1236), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(KEYINPUT62), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT62), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1236), .A2(new_n1241), .A3(new_n1242), .A4(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1244), .A2(new_n1246), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n990), .A2(new_n1002), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G390), .B1(new_n1251), .B2(new_n964), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G393), .A2(G396), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n964), .A3(G390), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n1214), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1214), .A2(new_n1254), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1255), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n1252), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1250), .A2(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1237), .B2(new_n1243), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1245), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1236), .A2(new_n1241), .A3(new_n1242), .A4(KEYINPUT63), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1262), .A2(new_n1263), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1261), .A2(new_n1267), .ZN(G405));
  NAND2_X1  g1068(.A1(G375), .A2(new_n1139), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1233), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(new_n1242), .A3(new_n1241), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1269), .B(new_n1233), .C1(new_n1240), .C2(new_n1239), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1271), .A2(new_n1260), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1260), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(G402));
endmodule


