

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  NOR2_X1 U323 ( .A1(n526), .A2(n475), .ZN(n566) );
  XNOR2_X1 U324 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U325 ( .A(n364), .B(n363), .ZN(n518) );
  XOR2_X1 U326 ( .A(n449), .B(n448), .Z(n291) );
  INV_X1 U327 ( .A(KEYINPUT47), .ZN(n462) );
  INV_X1 U328 ( .A(KEYINPUT100), .ZN(n353) );
  XNOR2_X1 U329 ( .A(n354), .B(n353), .ZN(n355) );
  INV_X1 U330 ( .A(n575), .ZN(n451) );
  NOR2_X1 U331 ( .A1(n542), .A2(n492), .ZN(n528) );
  INV_X1 U332 ( .A(KEYINPUT106), .ZN(n452) );
  XNOR2_X1 U333 ( .A(n450), .B(n291), .ZN(n575) );
  XNOR2_X1 U334 ( .A(n575), .B(KEYINPUT41), .ZN(n549) );
  XNOR2_X1 U335 ( .A(n452), .B(KEYINPUT38), .ZN(n453) );
  INV_X1 U336 ( .A(G190GAT), .ZN(n476) );
  XNOR2_X1 U337 ( .A(n454), .B(n453), .ZN(n498) );
  XNOR2_X1 U338 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U339 ( .A(n455), .B(G43GAT), .ZN(n456) );
  XNOR2_X1 U340 ( .A(n479), .B(n478), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n457), .B(n456), .ZN(G1330GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT90), .B(G127GAT), .Z(n293) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(G183GAT), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n311) );
  XOR2_X1 U345 ( .A(KEYINPUT94), .B(G99GAT), .Z(n295) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U348 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n297) );
  XNOR2_X1 U349 ( .A(G15GAT), .B(G71GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U351 ( .A(n299), .B(n298), .Z(n309) );
  XNOR2_X1 U352 ( .A(KEYINPUT93), .B(KEYINPUT19), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n300), .B(KEYINPUT17), .ZN(n301) );
  XOR2_X1 U354 ( .A(n301), .B(KEYINPUT92), .Z(n303) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n364) );
  XNOR2_X1 U357 ( .A(G134GAT), .B(G120GAT), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n304), .B(KEYINPUT0), .ZN(n338) );
  XOR2_X1 U359 ( .A(n338), .B(G176GAT), .Z(n306) );
  NAND2_X1 U360 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n364), .B(n307), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n526) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n312), .B(G36GAT), .ZN(n313) );
  XOR2_X1 U367 ( .A(n313), .B(KEYINPUT7), .Z(n315) );
  XNOR2_X1 U368 ( .A(G50GAT), .B(KEYINPUT68), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n426) );
  XOR2_X1 U370 ( .A(KEYINPUT82), .B(KEYINPUT10), .Z(n317) );
  XNOR2_X1 U371 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n322) );
  XNOR2_X1 U373 ( .A(G190GAT), .B(G92GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n318), .B(KEYINPUT83), .ZN(n356) );
  XOR2_X1 U375 ( .A(n356), .B(G134GAT), .Z(n320) );
  NAND2_X1 U376 ( .A1(G232GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U378 ( .A(n322), .B(n321), .Z(n329) );
  XOR2_X1 U379 ( .A(KEYINPUT77), .B(G85GAT), .Z(n324) );
  XNOR2_X1 U380 ( .A(G99GAT), .B(G106GAT), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n433) );
  XOR2_X1 U382 ( .A(KEYINPUT81), .B(KEYINPUT11), .Z(n326) );
  XNOR2_X1 U383 ( .A(G29GAT), .B(G162GAT), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n433), .B(n327), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n426), .B(n330), .ZN(n557) );
  XNOR2_X1 U388 ( .A(KEYINPUT36), .B(n557), .ZN(n584) );
  XOR2_X1 U389 ( .A(G127GAT), .B(G57GAT), .Z(n402) );
  XOR2_X1 U390 ( .A(KEYINPUT5), .B(G85GAT), .Z(n332) );
  XNOR2_X1 U391 ( .A(G155GAT), .B(G148GAT), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n402), .B(n333), .ZN(n335) );
  AND2_X1 U394 ( .A1(G225GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n337) );
  INV_X1 U396 ( .A(KEYINPUT98), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n338), .B(KEYINPUT1), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U400 ( .A(KEYINPUT4), .B(KEYINPUT97), .Z(n342) );
  XNOR2_X1 U401 ( .A(KEYINPUT6), .B(KEYINPUT96), .ZN(n341) );
  XOR2_X1 U402 ( .A(n342), .B(n341), .Z(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n349) );
  XOR2_X1 U404 ( .A(G1GAT), .B(G141GAT), .Z(n346) );
  XNOR2_X1 U405 ( .A(G29GAT), .B(G113GAT), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n425) );
  XNOR2_X1 U407 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n347), .B(KEYINPUT3), .ZN(n370) );
  XNOR2_X1 U409 ( .A(n425), .B(n370), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n391) );
  XNOR2_X1 U411 ( .A(KEYINPUT99), .B(n391), .ZN(n516) );
  XOR2_X1 U412 ( .A(KEYINPUT95), .B(G218GAT), .Z(n351) );
  XNOR2_X1 U413 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U415 ( .A(G197GAT), .B(n352), .Z(n378) );
  NAND2_X1 U416 ( .A1(G226GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n378), .B(n357), .ZN(n362) );
  XOR2_X1 U418 ( .A(G8GAT), .B(G183GAT), .Z(n396) );
  XNOR2_X1 U419 ( .A(G176GAT), .B(G64GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n358), .B(KEYINPUT78), .ZN(n435) );
  XOR2_X1 U421 ( .A(n396), .B(n435), .Z(n360) );
  XNOR2_X1 U422 ( .A(G36GAT), .B(G204GAT), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U425 ( .A(KEYINPUT27), .B(n518), .ZN(n387) );
  NOR2_X1 U426 ( .A1(n516), .A2(n387), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n365), .B(KEYINPUT101), .ZN(n542) );
  XOR2_X1 U428 ( .A(G148GAT), .B(G204GAT), .Z(n367) );
  XNOR2_X1 U429 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n436) );
  XOR2_X1 U431 ( .A(G155GAT), .B(G78GAT), .Z(n403) );
  XOR2_X1 U432 ( .A(n436), .B(n403), .Z(n369) );
  XNOR2_X1 U433 ( .A(G50GAT), .B(G106GAT), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n374) );
  XOR2_X1 U435 ( .A(G141GAT), .B(n370), .Z(n372) );
  NAND2_X1 U436 ( .A1(G228GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U438 ( .A(n374), .B(n373), .Z(n380) );
  XOR2_X1 U439 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n376) );
  XNOR2_X1 U440 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U442 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n473) );
  XNOR2_X1 U444 ( .A(n473), .B(KEYINPUT28), .ZN(n492) );
  XNOR2_X1 U445 ( .A(KEYINPUT102), .B(n528), .ZN(n381) );
  NAND2_X1 U446 ( .A1(n381), .A2(n526), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n382), .B(KEYINPUT103), .ZN(n393) );
  NOR2_X1 U448 ( .A1(n526), .A2(n518), .ZN(n383) );
  NOR2_X1 U449 ( .A1(n473), .A2(n383), .ZN(n384) );
  XOR2_X1 U450 ( .A(n384), .B(KEYINPUT25), .Z(n385) );
  XNOR2_X1 U451 ( .A(KEYINPUT104), .B(n385), .ZN(n389) );
  NAND2_X1 U452 ( .A1(n526), .A2(n473), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n386), .B(KEYINPUT26), .ZN(n570) );
  NOR2_X1 U454 ( .A1(n570), .A2(n387), .ZN(n388) );
  NOR2_X1 U455 ( .A1(n389), .A2(n388), .ZN(n390) );
  NOR2_X1 U456 ( .A1(n391), .A2(n390), .ZN(n392) );
  NOR2_X1 U457 ( .A1(n393), .A2(n392), .ZN(n481) );
  NOR2_X1 U458 ( .A1(n584), .A2(n481), .ZN(n415) );
  XOR2_X1 U459 ( .A(KEYINPUT12), .B(KEYINPUT86), .Z(n395) );
  XNOR2_X1 U460 ( .A(G64GAT), .B(KEYINPUT88), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n397) );
  XOR2_X1 U462 ( .A(n397), .B(n396), .Z(n399) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(G211GAT), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n401) );
  XNOR2_X1 U465 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n400), .B(KEYINPUT72), .ZN(n434) );
  XOR2_X1 U467 ( .A(n401), .B(n434), .Z(n405) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n414) );
  XOR2_X1 U470 ( .A(KEYINPUT15), .B(KEYINPUT84), .Z(n407) );
  XNOR2_X1 U471 ( .A(KEYINPUT14), .B(KEYINPUT85), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n412) );
  XNOR2_X1 U473 ( .A(G15GAT), .B(G22GAT), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n408), .B(KEYINPUT69), .ZN(n423) );
  XOR2_X1 U475 ( .A(n423), .B(KEYINPUT87), .Z(n410) );
  NAND2_X1 U476 ( .A1(G231GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U478 ( .A(n412), .B(n411), .Z(n413) );
  XNOR2_X1 U479 ( .A(n414), .B(n413), .ZN(n554) );
  NAND2_X1 U480 ( .A1(n415), .A2(n554), .ZN(n416) );
  XOR2_X1 U481 ( .A(KEYINPUT37), .B(n416), .Z(n514) );
  XOR2_X1 U482 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n418) );
  XNOR2_X1 U483 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U485 ( .A(G169GAT), .B(G197GAT), .Z(n419) );
  XNOR2_X1 U486 ( .A(n420), .B(n419), .ZN(n430) );
  XOR2_X1 U487 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n422) );
  XNOR2_X1 U488 ( .A(KEYINPUT70), .B(KEYINPUT64), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n422), .B(n421), .ZN(n424) );
  XOR2_X1 U490 ( .A(n424), .B(n423), .Z(n428) );
  XNOR2_X1 U491 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n432) );
  NAND2_X1 U494 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n571) );
  XOR2_X1 U496 ( .A(n571), .B(KEYINPUT71), .Z(n559) );
  XOR2_X1 U497 ( .A(n434), .B(n433), .Z(n438) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n450) );
  XOR2_X1 U500 ( .A(G92GAT), .B(G57GAT), .Z(n440) );
  XNOR2_X1 U501 ( .A(G120GAT), .B(G78GAT), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U503 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n442) );
  XNOR2_X1 U504 ( .A(KEYINPUT79), .B(KEYINPUT31), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U506 ( .A(n444), .B(n443), .Z(n449) );
  XOR2_X1 U507 ( .A(KEYINPUT80), .B(KEYINPUT74), .Z(n446) );
  NAND2_X1 U508 ( .A1(G230GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U509 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U510 ( .A(KEYINPUT73), .B(n447), .ZN(n448) );
  NAND2_X1 U511 ( .A1(n559), .A2(n451), .ZN(n480) );
  NOR2_X1 U512 ( .A1(n514), .A2(n480), .ZN(n454) );
  NOR2_X1 U513 ( .A1(n526), .A2(n498), .ZN(n457) );
  XNOR2_X1 U514 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n455) );
  INV_X1 U515 ( .A(n557), .ZN(n537) );
  INV_X1 U516 ( .A(n554), .ZN(n580) );
  XNOR2_X1 U517 ( .A(n580), .B(KEYINPUT114), .ZN(n565) );
  INV_X1 U518 ( .A(n549), .ZN(n561) );
  NAND2_X1 U519 ( .A1(n571), .A2(n561), .ZN(n458) );
  XOR2_X1 U520 ( .A(KEYINPUT46), .B(n458), .Z(n459) );
  NOR2_X1 U521 ( .A1(n565), .A2(n459), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n460), .B(KEYINPUT115), .ZN(n461) );
  NOR2_X1 U523 ( .A1(n537), .A2(n461), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(n462), .ZN(n469) );
  NOR2_X1 U525 ( .A1(n584), .A2(n554), .ZN(n464) );
  XOR2_X1 U526 ( .A(KEYINPUT45), .B(n464), .Z(n465) );
  NOR2_X1 U527 ( .A1(n575), .A2(n465), .ZN(n466) );
  XOR2_X1 U528 ( .A(KEYINPUT116), .B(n466), .Z(n467) );
  NOR2_X1 U529 ( .A1(n559), .A2(n467), .ZN(n468) );
  NOR2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U531 ( .A(KEYINPUT48), .B(n470), .ZN(n541) );
  NOR2_X1 U532 ( .A1(n518), .A2(n541), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n471), .B(KEYINPUT54), .ZN(n472) );
  NAND2_X1 U534 ( .A1(n472), .A2(n516), .ZN(n569) );
  NOR2_X1 U535 ( .A1(n473), .A2(n569), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n474), .B(KEYINPUT55), .ZN(n475) );
  NAND2_X1 U537 ( .A1(n566), .A2(n537), .ZN(n479) );
  XOR2_X1 U538 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n477) );
  INV_X1 U539 ( .A(n480), .ZN(n485) );
  XOR2_X1 U540 ( .A(KEYINPUT89), .B(KEYINPUT16), .Z(n483) );
  NAND2_X1 U541 ( .A1(n580), .A2(n557), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  NOR2_X1 U543 ( .A1(n481), .A2(n484), .ZN(n502) );
  NAND2_X1 U544 ( .A1(n485), .A2(n502), .ZN(n493) );
  NOR2_X1 U545 ( .A1(n516), .A2(n493), .ZN(n486) );
  XOR2_X1 U546 ( .A(KEYINPUT34), .B(n486), .Z(n487) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NOR2_X1 U548 ( .A1(n518), .A2(n493), .ZN(n488) );
  XOR2_X1 U549 ( .A(G8GAT), .B(n488), .Z(G1325GAT) );
  NOR2_X1 U550 ( .A1(n526), .A2(n493), .ZN(n490) );
  XNOR2_X1 U551 ( .A(KEYINPUT105), .B(KEYINPUT35), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U553 ( .A(G15GAT), .B(n491), .Z(G1326GAT) );
  INV_X1 U554 ( .A(n492), .ZN(n523) );
  NOR2_X1 U555 ( .A1(n523), .A2(n493), .ZN(n494) );
  XOR2_X1 U556 ( .A(G22GAT), .B(n494), .Z(G1327GAT) );
  NOR2_X1 U557 ( .A1(n516), .A2(n498), .ZN(n496) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NOR2_X1 U560 ( .A1(n518), .A2(n498), .ZN(n497) );
  XOR2_X1 U561 ( .A(G36GAT), .B(n497), .Z(G1329GAT) );
  NOR2_X1 U562 ( .A1(n523), .A2(n498), .ZN(n499) );
  XOR2_X1 U563 ( .A(G50GAT), .B(n499), .Z(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n501) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(n505) );
  INV_X1 U567 ( .A(n571), .ZN(n545) );
  NAND2_X1 U568 ( .A1(n561), .A2(n545), .ZN(n513) );
  INV_X1 U569 ( .A(n513), .ZN(n503) );
  NAND2_X1 U570 ( .A1(n503), .A2(n502), .ZN(n510) );
  NOR2_X1 U571 ( .A1(n516), .A2(n510), .ZN(n504) );
  XOR2_X1 U572 ( .A(n505), .B(n504), .Z(G1332GAT) );
  NOR2_X1 U573 ( .A1(n518), .A2(n510), .ZN(n506) );
  XOR2_X1 U574 ( .A(KEYINPUT110), .B(n506), .Z(n507) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  NOR2_X1 U576 ( .A1(n526), .A2(n510), .ZN(n509) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n508) );
  XNOR2_X1 U578 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  NOR2_X1 U579 ( .A1(n523), .A2(n510), .ZN(n512) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U581 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n514), .A2(n513), .ZN(n515) );
  XOR2_X1 U583 ( .A(KEYINPUT112), .B(n515), .Z(n522) );
  NOR2_X1 U584 ( .A1(n522), .A2(n516), .ZN(n517) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(KEYINPUT113), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1337GAT) );
  NOR2_X1 U589 ( .A1(n522), .A2(n526), .ZN(n521) );
  XOR2_X1 U590 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U591 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U592 ( .A(KEYINPUT44), .B(n524), .Z(n525) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n541), .ZN(n527) );
  NAND2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(KEYINPUT117), .B(n529), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n538), .A2(n559), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n530), .B(KEYINPUT118), .ZN(n531) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U601 ( .A1(n538), .A2(n561), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  NAND2_X1 U604 ( .A1(n565), .A2(n538), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U608 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  INV_X1 U610 ( .A(n541), .ZN(n544) );
  NOR2_X1 U611 ( .A1(n570), .A2(n542), .ZN(n543) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n556) );
  NOR2_X1 U613 ( .A1(n545), .A2(n556), .ZN(n546) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n548) );
  XNOR2_X1 U616 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n549), .A2(n556), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n554), .A2(n556), .ZN(n555) );
  XOR2_X1 U623 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  NAND2_X1 U626 ( .A1(n559), .A2(n566), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(n560), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n563) );
  NAND2_X1 U629 ( .A1(n566), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(n564), .ZN(G1349GAT) );
  XOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT123), .Z(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n573) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n582) );
  NAND2_X1 U637 ( .A1(n582), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n577) );
  NAND2_X1 U641 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n579) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT125), .Z(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n582), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U647 ( .A(n582), .ZN(n583) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

