//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n208), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n211), .B1(new_n214), .B2(new_n215), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n229), .B(new_n232), .Z(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G33), .ZN(new_n241));
  INV_X1    g0041(.A(G41), .ZN(new_n242));
  OAI211_X1 g0042(.A(G1), .B(G13), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G77), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n243), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G222), .A2(G1698), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT66), .B(G223), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n250), .B1(new_n251), .B2(G1698), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n249), .B1(new_n252), .B2(new_n247), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n243), .A2(new_n254), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n256), .B1(new_n257), .B2(G226), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G190), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT70), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n262), .A2(KEYINPUT67), .A3(new_n212), .ZN(new_n263));
  AOI21_X1  g0063(.A(KEYINPUT67), .B1(new_n262), .B2(new_n212), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G13), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n267), .A2(new_n206), .A3(G1), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n269), .B(G50), .C1(G1), .C2(new_n206), .ZN(new_n270));
  OAI21_X1  g0070(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n271));
  INV_X1    g0071(.A(G150), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n206), .A2(G33), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n271), .B1(new_n272), .B2(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G50), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n277), .A2(new_n266), .B1(new_n278), .B2(new_n268), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n270), .A2(new_n279), .A3(KEYINPUT9), .ZN(new_n280));
  INV_X1    g0080(.A(G200), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n259), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n270), .A2(new_n279), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT9), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n261), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  OR2_X1    g0086(.A1(new_n282), .A2(KEYINPUT71), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n287), .A2(KEYINPUT10), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n286), .B(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n283), .B1(new_n259), .B2(G169), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n290), .A2(KEYINPUT68), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n259), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n290), .B2(KEYINPUT68), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G68), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n273), .A2(G50), .B1(G20), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n248), .B2(new_n276), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n266), .A2(KEYINPUT11), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n268), .A2(new_n298), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT12), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n262), .A2(new_n212), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n205), .B2(G20), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G68), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT11), .B1(new_n266), .B2(new_n300), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT14), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT13), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT3), .B(G33), .ZN(new_n313));
  INV_X1    g0113(.A(G1698), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(G226), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT72), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT72), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n313), .A2(new_n317), .A3(G226), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n247), .A2(new_n226), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g0122(.A1(G33), .A2(G41), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n212), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n256), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT73), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n257), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n243), .A2(new_n254), .ZN(new_n329));
  OAI21_X1  g0129(.A(G238), .B1(new_n329), .B2(KEYINPUT73), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n326), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n312), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n243), .B1(new_n319), .B2(new_n321), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n334), .A2(new_n331), .A3(KEYINPUT13), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n311), .B(G169), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n325), .A2(new_n312), .A3(new_n332), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT13), .B1(new_n334), .B2(new_n331), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G179), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(new_n338), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n311), .B1(new_n341), .B2(G169), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n310), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(G200), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n344), .B(new_n309), .C1(new_n345), .C2(new_n341), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n313), .A2(G238), .A3(G1698), .ZN(new_n348));
  INV_X1    g0148(.A(G107), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n313), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n247), .A2(new_n226), .A3(G1698), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n324), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n256), .B1(new_n257), .B2(G244), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(G179), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT69), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G20), .A2(G77), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n357), .B1(new_n275), .B2(new_n274), .C1(new_n276), .C2(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n359), .A2(new_n304), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n305), .A2(G77), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n267), .A2(G1), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G20), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(G77), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n354), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n356), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n365), .ZN(new_n369));
  INV_X1    g0169(.A(new_n354), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(G190), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n354), .A2(G200), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n297), .A2(new_n347), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G58), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n298), .ZN(new_n377));
  OAI21_X1  g0177(.A(G20), .B1(new_n377), .B2(new_n201), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n273), .A2(G159), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT74), .B1(new_n241), .B2(KEYINPUT3), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT74), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n244), .A3(G33), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n383), .A3(new_n246), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT75), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n385), .B1(new_n313), .B2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n380), .B1(new_n392), .B2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT76), .B1(new_n393), .B2(KEYINPUT16), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n390), .A2(new_n391), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n389), .B1(new_n384), .B2(new_n386), .ZN(new_n396));
  OAI21_X1  g0196(.A(G68), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n380), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n247), .A2(new_n386), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT7), .B1(new_n247), .B2(new_n206), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n398), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n304), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n394), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n275), .B1(new_n205), .B2(G20), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n269), .A2(new_n410), .B1(new_n268), .B2(new_n275), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n326), .B1(new_n329), .B2(new_n226), .ZN(new_n414));
  MUX2_X1   g0214(.A(G223), .B(G226), .S(G1698), .Z(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n313), .ZN(new_n416));
  INV_X1    g0216(.A(G87), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n241), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n414), .B1(new_n418), .B2(new_n324), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(new_n366), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(G179), .B2(new_n419), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n412), .A2(new_n413), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n345), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(G200), .B2(new_n419), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n402), .A2(new_n408), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT16), .B1(new_n397), .B2(new_n398), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(new_n400), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n411), .B(new_n425), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n411), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n407), .B1(new_n427), .B2(new_n400), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n394), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT18), .B1(new_n434), .B2(new_n421), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(KEYINPUT17), .A3(new_n425), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n423), .A2(new_n431), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n375), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n304), .ZN(new_n440));
  OAI21_X1  g0240(.A(G107), .B1(new_n395), .B2(new_n396), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT6), .ZN(new_n442));
  INV_X1    g0242(.A(G97), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n442), .A2(new_n443), .A3(G107), .ZN(new_n444));
  XNOR2_X1  g0244(.A(G97), .B(G107), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n444), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n446), .A2(new_n206), .B1(new_n248), .B2(new_n274), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n440), .B1(new_n441), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT5), .B(G41), .ZN(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n450), .A2(new_n243), .A3(G274), .A4(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  NOR2_X1   g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n243), .ZN(new_n457));
  INV_X1    g0257(.A(G257), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n453), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n245), .A2(new_n246), .A3(G244), .A4(new_n314), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT77), .A2(KEYINPUT4), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n461), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n313), .A2(G244), .A3(new_n314), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n313), .A2(G250), .A3(G1698), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n462), .A2(new_n464), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n459), .B1(new_n467), .B2(new_n324), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n281), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n268), .A2(new_n443), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n241), .A2(G1), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n265), .A2(new_n363), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n470), .B1(new_n473), .B2(new_n443), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n449), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n467), .A2(new_n324), .ZN(new_n476));
  INV_X1    g0276(.A(new_n459), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT78), .B1(new_n478), .B2(new_n345), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT78), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n468), .A2(new_n480), .A3(G190), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n473), .A2(new_n443), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n447), .B1(new_n392), .B2(G107), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n470), .C1(new_n484), .C2(new_n440), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n476), .A2(new_n292), .A3(new_n477), .ZN(new_n486));
  AOI21_X1  g0286(.A(G169), .B1(new_n476), .B2(new_n477), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n475), .A2(new_n482), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n245), .A2(new_n246), .A3(new_n206), .A4(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT22), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT22), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n313), .A2(new_n492), .A3(new_n206), .A4(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT81), .B(KEYINPUT24), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G116), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(G20), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT23), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n206), .B2(G107), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n349), .A2(KEYINPUT23), .A3(G20), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n494), .A2(new_n495), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n495), .B1(new_n494), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n304), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n268), .A2(new_n349), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT25), .ZN(new_n506));
  INV_X1    g0306(.A(new_n473), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G107), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n245), .A2(new_n246), .A3(G257), .A4(G1698), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n245), .A2(new_n246), .A3(G250), .A4(new_n314), .ZN(new_n511));
  INV_X1    g0311(.A(G294), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n510), .B(new_n511), .C1(new_n241), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n324), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n324), .B1(new_n452), .B2(new_n450), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G264), .ZN(new_n516));
  AND4_X1   g0316(.A1(new_n345), .A2(new_n514), .A3(new_n453), .A4(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n513), .A2(new_n324), .B1(new_n515), .B2(G264), .ZN(new_n518));
  AOI21_X1  g0318(.A(G200), .B1(new_n518), .B2(new_n453), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT83), .B1(new_n509), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n514), .A2(new_n453), .A3(new_n516), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n281), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(G190), .B2(new_n522), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT83), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n524), .A2(new_n525), .A3(new_n504), .A4(new_n508), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n522), .A2(G169), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n518), .A2(G179), .A3(new_n453), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(KEYINPUT82), .B1(new_n504), .B2(new_n508), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT82), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n521), .A2(new_n526), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n362), .ZN(new_n534));
  INV_X1    g0334(.A(G116), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G20), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n268), .A2(new_n535), .A3(new_n471), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n440), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n466), .B(new_n206), .C1(G33), .C2(new_n443), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n304), .A3(new_n536), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT20), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n245), .A2(new_n246), .A3(G264), .A4(G1698), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT80), .B(G303), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n313), .B2(new_n547), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n247), .A2(new_n458), .A3(G1698), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n324), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n324), .A2(new_n255), .ZN(new_n551));
  INV_X1    g0351(.A(new_n456), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n515), .A2(G270), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n545), .B1(new_n554), .B2(G200), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n345), .B2(new_n554), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n545), .A3(G169), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT21), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n550), .A2(new_n553), .A3(G179), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n557), .A2(new_n558), .B1(new_n559), .B2(new_n545), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n554), .A2(new_n545), .A3(KEYINPUT21), .A4(G169), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n245), .A2(new_n246), .A3(G238), .A4(new_n314), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n245), .A2(new_n246), .A3(G244), .A4(G1698), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n496), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n324), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n205), .A2(G45), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n567), .B(G250), .C1(new_n323), .C2(new_n212), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n452), .A2(G274), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n566), .A2(new_n292), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT79), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n566), .A2(new_n571), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n366), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n570), .B1(new_n565), .B2(new_n324), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT79), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n577), .A3(new_n292), .ZN(new_n578));
  XOR2_X1   g0378(.A(KEYINPUT15), .B(G87), .Z(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n363), .ZN(new_n580));
  NAND3_X1  g0380(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n206), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n417), .A2(new_n443), .A3(new_n349), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n245), .A2(new_n246), .A3(new_n206), .A4(G68), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n276), .B2(new_n443), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n580), .B1(new_n588), .B2(new_n304), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n265), .A2(new_n363), .A3(new_n579), .A4(new_n472), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n573), .A2(new_n575), .A3(new_n578), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n574), .A2(G200), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n576), .A2(G190), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n265), .A2(G87), .A3(new_n363), .A4(new_n472), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n589), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n562), .A2(new_n597), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n439), .A2(new_n489), .A3(new_n533), .A4(new_n598), .ZN(G372));
  NAND2_X1  g0399(.A1(new_n423), .A2(new_n435), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n343), .ZN(new_n602));
  INV_X1    g0402(.A(new_n368), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n602), .B1(new_n346), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n431), .A2(new_n436), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n295), .B1(new_n606), .B2(new_n289), .ZN(new_n607));
  INV_X1    g0407(.A(new_n439), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n345), .B(new_n570), .C1(new_n565), .C2(new_n324), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n589), .A2(new_n595), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT84), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n568), .B2(new_n569), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n568), .A2(new_n612), .A3(new_n569), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n566), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G200), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n589), .A2(new_n590), .B1(new_n576), .B2(new_n292), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n366), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n611), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n485), .A4(new_n488), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n591), .A2(new_n572), .ZN(new_n623));
  INV_X1    g0423(.A(new_n613), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n614), .ZN(new_n625));
  AOI21_X1  g0425(.A(G169), .B1(new_n625), .B2(new_n566), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n592), .A2(new_n596), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n441), .A2(new_n448), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n474), .B1(new_n631), .B2(new_n304), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n476), .A2(new_n477), .A3(new_n292), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(G169), .B2(new_n468), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n621), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT86), .B1(new_n629), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n478), .A2(new_n366), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n638), .B(new_n633), .C1(new_n449), .C2(new_n474), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT26), .B1(new_n639), .B2(new_n597), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT86), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n628), .A4(new_n622), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n521), .A2(new_n526), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n489), .A2(new_n643), .A3(new_n620), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n557), .A2(new_n558), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n559), .A2(new_n545), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n561), .A3(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n504), .A2(new_n508), .B1(new_n527), .B2(new_n528), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT85), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n509), .A2(new_n529), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT85), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(new_n561), .A4(new_n560), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n637), .A2(new_n642), .B1(new_n644), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n607), .B1(new_n608), .B2(new_n654), .ZN(G369));
  OAI21_X1  g0455(.A(KEYINPUT27), .B1(new_n534), .B2(G20), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n362), .A2(new_n657), .A3(new_n206), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT87), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(KEYINPUT88), .B(G343), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT89), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n659), .B(KEYINPUT87), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  INV_X1    g0465(.A(new_n662), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n509), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n533), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n530), .A2(new_n532), .A3(new_n668), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(new_n545), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n645), .A2(new_n561), .A3(new_n646), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n556), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n675), .B2(new_n674), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n675), .A2(new_n668), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n533), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n668), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n648), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n209), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n583), .A2(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n215), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT91), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n476), .A2(new_n518), .A3(new_n477), .A4(new_n576), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n550), .A2(new_n553), .A3(G179), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n518), .A2(new_n576), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n559), .A3(KEYINPUT30), .A4(new_n468), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n696), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n559), .A3(new_n468), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT91), .B1(new_n704), .B2(new_n697), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n554), .A2(new_n292), .A3(new_n616), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n514), .A2(new_n453), .A3(new_n516), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT90), .B1(new_n707), .B2(new_n468), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT90), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n478), .A2(new_n709), .A3(new_n522), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n706), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n703), .A2(new_n705), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n695), .B1(new_n712), .B2(new_n683), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n533), .A2(new_n598), .A3(new_n489), .A4(new_n683), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n700), .A2(new_n702), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT31), .B(new_n668), .C1(new_n715), .C2(new_n711), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n637), .A2(new_n642), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n594), .A2(new_n589), .A3(new_n595), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n281), .B1(new_n625), .B2(new_n566), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n721), .A2(new_n722), .B1(new_n623), .B2(new_n626), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n521), .B2(new_n526), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n489), .A3(new_n649), .A4(new_n652), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n668), .B1(new_n720), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT92), .B1(new_n654), .B2(new_n668), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n529), .A2(KEYINPUT82), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n509), .A3(new_n532), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n675), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n724), .A2(new_n489), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n630), .A2(new_n635), .A3(new_n621), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT26), .B1(new_n639), .B2(new_n723), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(new_n628), .A3(new_n738), .ZN(new_n739));
  OAI211_X1 g0539(.A(KEYINPUT29), .B(new_n683), .C1(new_n736), .C2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n719), .B1(new_n731), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n694), .B1(new_n741), .B2(G1), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT93), .ZN(G364));
  NOR2_X1   g0543(.A1(new_n267), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT94), .B1(new_n744), .B2(G45), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n205), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(KEYINPUT94), .A3(G45), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n689), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n677), .B2(G330), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G330), .B2(new_n677), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n209), .A2(new_n313), .ZN(new_n752));
  INV_X1    g0552(.A(G355), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n752), .A2(new_n753), .B1(G116), .B2(new_n209), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n688), .A2(new_n313), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n215), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n451), .B2(new_n757), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n236), .A2(new_n451), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n754), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n212), .B1(G20), .B2(new_n366), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n749), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n206), .A2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n281), .A2(G179), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(G20), .A3(G190), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n313), .B1(new_n770), .B2(new_n349), .C1(new_n417), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G179), .A2(G200), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n206), .B1(new_n773), .B2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G97), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n206), .A2(new_n292), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n345), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n778), .A2(G190), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n776), .B1(new_n780), .B2(new_n278), .C1(new_n298), .C2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n777), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n785));
  AOI21_X1  g0585(.A(G200), .B1(new_n784), .B2(KEYINPUT95), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n785), .A2(new_n345), .A3(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n772), .B(new_n783), .C1(G77), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n768), .A2(new_n773), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n790), .A2(KEYINPUT97), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(KEYINPUT97), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n785), .A2(G190), .A3(new_n786), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT96), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n789), .B(new_n796), .C1(new_n376), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G326), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n780), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(KEYINPUT33), .A2(G317), .ZN(new_n802));
  NAND2_X1  g0602(.A1(KEYINPUT33), .A2(G317), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n782), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n801), .B(new_n804), .C1(G294), .C2(new_n775), .ZN(new_n805));
  INV_X1    g0605(.A(new_n793), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G329), .ZN(new_n807));
  INV_X1    g0607(.A(G303), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n247), .B1(new_n771), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n770), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G283), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n805), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  INV_X1    g0613(.A(G322), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n813), .A2(new_n787), .B1(new_n797), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n799), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n767), .B1(new_n816), .B2(new_n764), .ZN(new_n817));
  INV_X1    g0617(.A(new_n763), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n677), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n751), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NOR2_X1   g0621(.A1(new_n368), .A2(new_n668), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n668), .A2(new_n369), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n373), .A2(new_n823), .B1(new_n356), .B2(new_n367), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n728), .B(new_n729), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n639), .A2(new_n723), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n627), .B1(new_n826), .B2(new_n621), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n641), .B1(new_n827), .B2(new_n640), .ZN(new_n828));
  INV_X1    g0628(.A(new_n642), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n725), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n822), .A2(new_n824), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n830), .A2(new_n683), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n719), .B1(new_n825), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n825), .A2(new_n719), .A3(new_n832), .ZN(new_n834));
  INV_X1    g0634(.A(new_n749), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n833), .B1(new_n836), .B2(KEYINPUT99), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(KEYINPUT99), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n764), .A2(new_n761), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n835), .B1(new_n248), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n771), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n313), .B1(new_n841), .B2(G107), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n842), .B1(new_n417), .B2(new_n770), .C1(new_n793), .C2(new_n813), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n776), .B1(new_n780), .B2(new_n808), .C1(new_n844), .C2(new_n782), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n535), .A2(new_n787), .B1(new_n797), .B2(new_n512), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n793), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n247), .B1(new_n841), .B2(G50), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n810), .A2(G68), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n850), .B(new_n851), .C1(new_n376), .C2(new_n774), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n781), .A2(G150), .B1(new_n779), .B2(G137), .ZN(new_n853));
  INV_X1    g0653(.A(G143), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n794), .B2(new_n787), .C1(new_n798), .C2(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(KEYINPUT98), .B(KEYINPUT34), .Z(new_n856));
  AOI211_X1 g0656(.A(new_n849), .B(new_n852), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n847), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n764), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n840), .B1(new_n859), .B2(new_n860), .C1(new_n831), .C2(new_n762), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n838), .A2(new_n861), .ZN(G384));
  NOR2_X1   g0662(.A1(new_n744), .A2(new_n205), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n705), .A2(new_n711), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT31), .B(new_n668), .C1(new_n864), .C2(new_n703), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n713), .A2(new_n714), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n668), .A2(new_n310), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n343), .A2(new_n346), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n310), .B(new_n668), .C1(new_n340), .C2(new_n342), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n866), .A2(new_n870), .A3(new_n831), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n406), .A2(new_n266), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n405), .B2(new_n398), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n411), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n874), .A2(new_n664), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n437), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n412), .A2(new_n422), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n412), .A2(new_n664), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n429), .ZN(new_n880));
  INV_X1    g0680(.A(new_n429), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n421), .A2(new_n661), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n882), .A2(new_n874), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT37), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n429), .B1(new_n434), .B2(new_n421), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n434), .A2(new_n661), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n880), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n888), .B1(new_n600), .B2(new_n605), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n871), .B1(new_n886), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n876), .A2(new_n885), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  AND4_X1   g0699(.A1(new_n899), .A2(new_n866), .A3(new_n870), .A4(new_n831), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n893), .A2(KEYINPUT40), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n439), .A2(new_n866), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(G330), .A3(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT100), .Z(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n886), .B2(new_n892), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n896), .A2(KEYINPUT39), .A3(new_n897), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n602), .A2(new_n683), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n601), .A2(new_n664), .ZN(new_n914));
  INV_X1    g0714(.A(new_n870), .ZN(new_n915));
  INV_X1    g0715(.A(new_n822), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n832), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n914), .B1(new_n898), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n731), .A2(new_n439), .A3(new_n740), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n607), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n863), .B1(new_n907), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n907), .B2(new_n922), .ZN(new_n924));
  INV_X1    g0724(.A(new_n446), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n925), .A2(KEYINPUT35), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(KEYINPUT35), .ZN(new_n927));
  NOR4_X1   g0727(.A1(new_n926), .A2(new_n927), .A3(new_n535), .A4(new_n214), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT36), .Z(new_n929));
  OR3_X1    g0729(.A1(new_n215), .A2(new_n248), .A3(new_n377), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n278), .A2(G68), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(G1), .A3(new_n267), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n924), .A2(new_n929), .A3(new_n933), .ZN(G367));
  NOR2_X1   g0734(.A1(new_n774), .A2(new_n298), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n780), .A2(new_n854), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(G159), .C2(new_n781), .ZN(new_n937));
  INV_X1    g0737(.A(new_n797), .ZN(new_n938));
  AOI22_X1  g0738(.A1(G50), .A2(new_n788), .B1(new_n938), .B2(G150), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n770), .A2(new_n248), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n247), .B(new_n940), .C1(G58), .C2(new_n841), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n806), .A2(G137), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n937), .A2(new_n939), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT46), .B1(new_n841), .B2(G116), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT107), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(G283), .B2(new_n788), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n841), .A2(KEYINPUT46), .A3(G116), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n780), .B2(new_n813), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G294), .B2(new_n781), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n247), .B1(new_n774), .B2(new_n349), .C1(new_n443), .C2(new_n770), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n806), .B2(G317), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n946), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n798), .A2(new_n547), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n943), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT47), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n764), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n668), .A2(new_n610), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n620), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n628), .B2(new_n957), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(new_n818), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n765), .B1(new_n209), .B2(new_n358), .C1(new_n756), .C2(new_n232), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n961), .A2(KEYINPUT106), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(KEYINPUT106), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n962), .A2(new_n963), .A3(new_n835), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n956), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n668), .A2(new_n485), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n489), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n635), .A2(new_n668), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n680), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT42), .B1(new_n970), .B2(new_n682), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n639), .B1(new_n967), .B2(new_n733), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n683), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT42), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n969), .A2(new_n976), .A3(new_n533), .A4(new_n681), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n973), .A2(new_n975), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT101), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n973), .A2(new_n975), .A3(new_n977), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT103), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n959), .B(KEYINPUT43), .Z(new_n985));
  NAND3_X1  g0785(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n984), .B1(new_n983), .B2(new_n985), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n981), .B(new_n982), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(KEYINPUT102), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT102), .ZN(new_n991));
  INV_X1    g0791(.A(new_n988), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n986), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n979), .B(KEYINPUT101), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n972), .B1(new_n990), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n989), .A2(KEYINPUT102), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n993), .A2(new_n994), .A3(new_n991), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n971), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT104), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1001), .B(KEYINPUT44), .C1(new_n686), .C2(new_n969), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT44), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1001), .A2(KEYINPUT44), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n970), .A2(new_n685), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT45), .B1(new_n686), .B2(new_n969), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n685), .A2(new_n970), .A3(new_n1007), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1002), .B(new_n1005), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n679), .A2(KEYINPUT105), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n682), .B1(new_n672), .B2(new_n681), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(new_n678), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n741), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n689), .B(KEYINPUT41), .Z(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n748), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n965), .B1(new_n1000), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT108), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT108), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n965), .C1(new_n1000), .C2(new_n1017), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1019), .A2(new_n1021), .ZN(G387));
  INV_X1    g0822(.A(new_n1013), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n673), .A2(new_n763), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n752), .A2(new_n691), .B1(G107), .B2(new_n209), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n229), .A2(G45), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT109), .Z(new_n1027));
  NOR3_X1   g0827(.A1(new_n275), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT50), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n275), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1029), .B1(new_n1030), .B2(new_n278), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n691), .B(new_n451), .C1(new_n298), .C2(new_n248), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1028), .B(new_n1031), .C1(new_n1033), .C2(KEYINPUT110), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n756), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1025), .B1(new_n1027), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n749), .B1(new_n1037), .B2(new_n766), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n775), .A2(new_n579), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n780), .B2(new_n794), .C1(new_n275), .C2(new_n782), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n793), .A2(new_n272), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n313), .B1(new_n770), .B2(new_n443), .C1(new_n248), .C2(new_n771), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n278), .B2(new_n797), .C1(new_n298), .C2(new_n787), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n313), .B1(new_n810), .B2(G116), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n771), .A2(new_n512), .B1(new_n774), .B2(new_n844), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n781), .A2(G311), .B1(new_n779), .B2(G322), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n547), .B2(new_n787), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n798), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1048), .B1(new_n1049), .B2(G317), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1046), .B1(new_n1050), .B2(KEYINPUT48), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(KEYINPUT48), .B2(new_n1050), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1045), .B1(new_n800), .B2(new_n793), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1044), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1038), .B1(new_n1056), .B2(new_n764), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1023), .A2(new_n748), .B1(new_n1024), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n741), .A2(new_n1023), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n689), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n741), .A2(new_n1023), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1058), .B1(new_n1060), .B2(new_n1061), .ZN(G393));
  OAI21_X1  g0862(.A(new_n689), .B1(new_n1011), .B2(new_n1059), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1009), .B(new_n679), .ZN(new_n1064));
  AOI21_X1  g0864(.A(KEYINPUT111), .B1(new_n1064), .B2(new_n1059), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1059), .A3(KEYINPUT111), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n748), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n970), .A2(new_n763), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n765), .B1(new_n443), .B2(new_n209), .C1(new_n756), .C2(new_n239), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n749), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n774), .A2(new_n248), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n313), .B1(new_n770), .B2(new_n417), .C1(new_n298), .C2(new_n771), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(G50), .C2(new_n781), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n854), .B2(new_n793), .C1(new_n275), .C2(new_n787), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n797), .A2(new_n794), .B1(new_n272), .B2(new_n780), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT51), .Z(new_n1079));
  AOI22_X1  g0879(.A1(new_n938), .A2(G311), .B1(G317), .B2(new_n779), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT52), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n782), .A2(new_n547), .B1(new_n535), .B2(new_n774), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n247), .B1(new_n770), .B2(new_n349), .C1(new_n844), .C2(new_n771), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n512), .B2(new_n787), .C1(new_n814), .C2(new_n793), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1077), .A2(new_n1079), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1073), .B1(new_n1086), .B2(new_n764), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1070), .B1(new_n1071), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1068), .A2(new_n1088), .ZN(G390));
  NAND3_X1  g0889(.A1(new_n439), .A2(G330), .A3(new_n866), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n920), .A2(new_n1090), .A3(new_n607), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n737), .A2(new_n628), .A3(new_n738), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n668), .B(new_n824), .C1(new_n1092), .C2(new_n735), .ZN(new_n1093));
  OAI21_X1  g0893(.A(KEYINPUT112), .B1(new_n1093), .B2(new_n822), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n824), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n683), .B(new_n1095), .C1(new_n736), .C2(new_n739), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT112), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n916), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n717), .A2(new_n831), .A3(G330), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1094), .A2(new_n1098), .B1(new_n1099), .B2(new_n870), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n866), .A2(G330), .A3(new_n831), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n915), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n866), .A2(new_n870), .A3(G330), .A4(new_n831), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n1099), .B2(new_n870), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n822), .B1(new_n726), .B2(new_n831), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1100), .A2(new_n1102), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1091), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT113), .B1(new_n917), .B2(new_n912), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n909), .A2(new_n910), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT113), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n911), .C1(new_n1105), .C2(new_n915), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1110), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1099), .A2(new_n870), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1094), .A2(new_n870), .A3(new_n1098), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n880), .A2(new_n889), .B1(new_n437), .B2(new_n888), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n897), .B1(new_n1117), .B2(KEYINPUT38), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n1118), .A3(new_n911), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1114), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1103), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1109), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1114), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1094), .A2(new_n870), .A3(new_n1098), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1118), .A2(new_n911), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n911), .B1(new_n1105), .B2(new_n915), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1127), .A2(KEYINPUT113), .B1(new_n909), .B2(new_n910), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1126), .B1(new_n1128), .B2(new_n1113), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1123), .B(new_n1108), .C1(new_n1129), .C2(new_n1103), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1122), .A2(new_n689), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1111), .A2(new_n761), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n839), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n749), .B1(new_n1030), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n313), .B1(new_n770), .B2(new_n278), .ZN(new_n1135));
  INV_X1    g0935(.A(G137), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n782), .A2(new_n1136), .B1(new_n774), .B2(new_n794), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(G128), .C2(new_n779), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n806), .A2(G125), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n771), .A2(new_n272), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT53), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G132), .A2(new_n938), .B1(new_n788), .B2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .A4(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n313), .B(new_n1074), .C1(G87), .C2(new_n841), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n781), .A2(G107), .B1(new_n779), .B2(G283), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n443), .B2(new_n787), .C1(new_n535), .C2(new_n797), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n851), .B1(new_n793), .B2(new_n512), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT114), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1145), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1134), .B1(new_n1152), .B2(new_n764), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1132), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n748), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT115), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1131), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1131), .B2(new_n1156), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(G378));
  XOR2_X1   g0960(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1161));
  XOR2_X1   g0961(.A(new_n297), .B(new_n1161), .Z(new_n1162));
  NAND2_X1  g0962(.A1(new_n283), .A2(new_n664), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT118), .Z(new_n1164));
  OR2_X1    g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n761), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n787), .A2(new_n358), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n935), .B1(G58), .B2(new_n810), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n780), .B2(new_n535), .C1(new_n443), .C2(new_n782), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(G107), .C2(new_n938), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G41), .B(new_n313), .C1(new_n841), .C2(G77), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT116), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n806), .A2(G283), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1173), .A2(KEYINPUT116), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT58), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n242), .B1(new_n244), .B2(new_n241), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1177), .A2(new_n1178), .B1(new_n278), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n1178), .B2(new_n1177), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n806), .A2(G124), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G33), .B(G41), .C1(new_n810), .C2(G159), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n779), .A2(G125), .B1(new_n841), .B2(new_n1143), .ZN(new_n1184));
  INV_X1    g0984(.A(G128), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1184), .B1(new_n272), .B2(new_n774), .C1(new_n797), .C2(new_n1185), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n787), .A2(new_n1136), .B1(new_n848), .B2(new_n782), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT117), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(KEYINPUT117), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1186), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT59), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1182), .B(new_n1183), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1191), .B2(new_n1190), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n764), .B1(new_n1181), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n835), .B1(new_n278), .B2(new_n839), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1168), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(G330), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n893), .A2(KEYINPUT40), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n898), .A2(new_n900), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n919), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n913), .B(new_n918), .C1(new_n901), .C2(new_n1198), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT119), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1197), .B1(new_n1209), .B2(new_n748), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1091), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1130), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1209), .A2(new_n1212), .A3(KEYINPUT57), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n689), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1208), .A2(new_n1207), .B1(new_n1130), .B2(new_n1211), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT57), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1210), .B1(new_n1214), .B2(new_n1216), .ZN(G375));
  NAND2_X1  g1017(.A1(new_n1091), .A2(new_n1107), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1109), .A2(new_n1016), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1107), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n915), .A2(new_n761), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n749), .B1(G68), .B2(new_n1133), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1039), .B1(new_n780), .B2(new_n512), .C1(new_n535), .C2(new_n782), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G107), .A2(new_n788), .B1(new_n938), .B2(G283), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n806), .A2(G303), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n313), .B(new_n940), .C1(G97), .C2(new_n841), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n313), .B1(new_n770), .B2(new_n376), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n782), .A2(new_n1142), .B1(new_n278), .B2(new_n774), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(G159), .C2(new_n841), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n806), .A2(G128), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n779), .A2(G132), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT120), .Z(new_n1234));
  NAND2_X1  g1034(.A1(new_n788), .A2(G150), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1231), .A2(new_n1232), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n798), .A2(new_n1136), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1228), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT121), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n860), .B1(new_n1238), .B2(KEYINPUT121), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1222), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1220), .A2(new_n748), .B1(new_n1221), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1219), .A2(new_n1242), .ZN(G381));
  AND3_X1   g1043(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1205), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1196), .B1(new_n1246), .B2(new_n1069), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n690), .B1(new_n1215), .B2(KEYINPUT57), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT57), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1130), .A2(new_n1211), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1246), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1247), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1131), .A2(new_n1156), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  OR2_X1    g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1256), .ZN(new_n1257));
  OR3_X1    g1057(.A1(new_n1255), .A2(G387), .A3(new_n1257), .ZN(G407));
  NAND2_X1  g1058(.A1(new_n662), .A2(G213), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT122), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G407), .B(G213), .C1(new_n1255), .C2(new_n1261), .ZN(G409));
  INV_X1    g1062(.A(KEYINPUT127), .ZN(new_n1263));
  INV_X1    g1063(.A(G390), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1019), .A2(new_n1021), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n965), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n996), .A2(new_n999), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1017), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1269), .A2(G390), .B1(new_n1256), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1265), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1256), .A2(new_n1270), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1269), .A2(G390), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1018), .A2(KEYINPUT124), .A3(new_n1068), .A4(new_n1088), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT124), .B1(new_n1264), .B2(new_n1018), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1275), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1265), .A2(new_n1271), .A3(KEYINPUT125), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1274), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1251), .A2(new_n689), .A3(new_n1213), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1253), .A2(KEYINPUT115), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1131), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .A4(new_n1210), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1215), .A2(new_n1016), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1210), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1254), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1260), .B1(new_n1287), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT123), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1218), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT60), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1218), .A2(new_n1292), .A3(KEYINPUT60), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(new_n689), .A3(new_n1109), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1242), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n838), .A2(new_n861), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(G384), .A3(new_n1242), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1283), .B1(new_n1291), .B2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1253), .B1(new_n1288), .B2(new_n1210), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1252), .B2(G378), .ZN(new_n1307));
  NOR4_X1   g1107(.A1(new_n1307), .A2(KEYINPUT62), .A3(new_n1260), .A4(new_n1303), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1260), .A2(G2897), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1298), .A2(G384), .A3(new_n1242), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G384), .B1(new_n1298), .B2(new_n1242), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1312), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1301), .A2(new_n1302), .A3(new_n1311), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1290), .B1(G375), .B2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1317), .B1(new_n1261), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1310), .B1(new_n1320), .B2(KEYINPUT61), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1282), .B1(new_n1309), .B2(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1316), .B(new_n1315), .C1(new_n1307), .C2(new_n1260), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1274), .A2(new_n1280), .A3(new_n1310), .A4(new_n1281), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1323), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1319), .A2(new_n1261), .A3(new_n1304), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1291), .A2(KEYINPUT63), .A3(new_n1304), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1326), .B1(new_n1331), .B2(new_n1282), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1263), .B1(new_n1322), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1282), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1327), .A2(KEYINPUT62), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1291), .A2(new_n1283), .A3(new_n1304), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT126), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1334), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT63), .B1(new_n1291), .B2(new_n1304), .ZN(new_n1340));
  NOR4_X1   g1140(.A1(new_n1307), .A2(new_n1328), .A3(new_n1260), .A4(new_n1303), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1282), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1326), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1339), .A2(new_n1344), .A3(KEYINPUT127), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1333), .A2(new_n1345), .ZN(G405));
  OAI21_X1  g1146(.A(new_n1287), .B1(new_n1253), .B2(new_n1252), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1347), .B(new_n1303), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(new_n1348), .B(new_n1282), .ZN(G402));
endmodule


