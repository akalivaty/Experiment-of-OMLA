//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G128), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n188), .A3(G143), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT64), .B1(new_n190), .B2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n190), .A2(G146), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(G128), .B1(new_n199), .B2(new_n193), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT67), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n204), .A3(new_n201), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n195), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G134), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G137), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n208), .B1(KEYINPUT11), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(G134), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT66), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(KEYINPUT66), .B(new_n214), .C1(new_n209), .C2(G137), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n211), .B(new_n212), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n210), .B2(new_n208), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n206), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n218), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n210), .B2(KEYINPUT11), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n216), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n212), .B1(new_n225), .B2(new_n211), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT69), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n211), .B1(new_n215), .B2(new_n217), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(new_n218), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n200), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n200), .A2(KEYINPUT65), .A3(new_n236), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n239), .A2(new_n240), .B1(new_n234), .B2(new_n192), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n221), .B1(new_n232), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G116), .B(G119), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n244), .A2(KEYINPUT68), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT2), .B(G113), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n245), .B(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT28), .B1(new_n242), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n242), .B2(new_n248), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n229), .A2(new_n230), .A3(new_n218), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n230), .B1(new_n229), .B2(new_n218), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n241), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n205), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n204), .B1(new_n200), .B2(new_n201), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n194), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n220), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n248), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(KEYINPUT73), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n254), .A2(new_n259), .A3(new_n248), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n251), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n249), .B1(new_n264), .B2(KEYINPUT28), .ZN(new_n265));
  INV_X1    g079(.A(G237), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G210), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT27), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(G902), .B1(new_n265), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n240), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT65), .B1(new_n200), .B2(new_n236), .ZN(new_n277));
  INV_X1    g091(.A(new_n192), .ZN(new_n278));
  OAI22_X1  g092(.A1(new_n276), .A2(new_n277), .B1(new_n233), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n227), .B2(new_n231), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT30), .B1(new_n280), .B2(new_n221), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n229), .A2(new_n218), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n241), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n259), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n248), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n263), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n272), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n263), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n248), .B1(new_n283), .B2(new_n259), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n291), .B1(new_n242), .B2(new_n248), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n290), .B1(new_n292), .B2(new_n289), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n271), .B(KEYINPUT70), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n288), .B(new_n273), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n187), .B1(new_n275), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n283), .A2(new_n259), .A3(new_n284), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n260), .B2(KEYINPUT30), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n263), .B(new_n271), .C1(new_n299), .C2(new_n248), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n281), .A2(new_n285), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n287), .B1(new_n303), .B2(new_n261), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(KEYINPUT31), .A3(new_n271), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n283), .A2(new_n259), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n261), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n289), .B1(new_n263), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n294), .B1(new_n309), .B2(new_n249), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n293), .A2(KEYINPUT71), .A3(new_n294), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI211_X1 g128(.A(G472), .B(G902), .C1(new_n306), .C2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n297), .B1(new_n315), .B2(KEYINPUT72), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n310), .A2(new_n311), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT71), .B1(new_n293), .B2(new_n294), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT31), .B1(new_n304), .B2(new_n271), .ZN(new_n319));
  NOR4_X1   g133(.A1(new_n286), .A2(new_n287), .A3(new_n301), .A4(new_n272), .ZN(new_n320));
  OAI22_X1  g134(.A1(new_n317), .A2(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n187), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT32), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n296), .B1(new_n316), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT22), .B(G137), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT74), .B(G125), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT16), .ZN(new_n332));
  INV_X1    g146(.A(G140), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(G125), .A2(G140), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n331), .B2(G140), .ZN(new_n336));
  OAI211_X1 g150(.A(G146), .B(new_n334), .C1(new_n336), .C2(new_n332), .ZN(new_n337));
  XOR2_X1   g151(.A(G125), .B(G140), .Z(new_n338));
  OR2_X1    g152(.A1(new_n338), .A2(G146), .ZN(new_n339));
  INV_X1    g153(.A(G128), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G119), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G128), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT24), .B(G110), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n340), .A2(KEYINPUT23), .A3(G119), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n343), .A3(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT76), .B(G110), .Z(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n337), .B(new_n339), .C1(new_n346), .C2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n334), .B1(new_n336), .B2(new_n332), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n188), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n337), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n344), .A2(new_n345), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(G110), .B2(new_n350), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n356), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n353), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n330), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n363), .B2(new_n362), .ZN(new_n365));
  OR3_X1    g179(.A1(new_n362), .A2(new_n363), .A3(new_n329), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G217), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(G234), .B2(new_n322), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n367), .B2(new_n368), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n365), .A2(new_n366), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n371), .A2(G902), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n326), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(G214), .B1(G237), .B2(G902), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n380), .B(KEYINPUT85), .Z(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G210), .B1(G237), .B2(G902), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT81), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G104), .ZN(new_n388));
  AOI21_X1  g202(.A(G107), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT82), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT81), .B(G104), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n392), .B(KEYINPUT3), .C1(new_n393), .C2(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n386), .A2(new_n388), .A3(G107), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n390), .A2(new_n397), .A3(G104), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n384), .B1(new_n401), .B2(G101), .ZN(new_n402));
  INV_X1    g216(.A(G101), .ZN(new_n403));
  AND4_X1   g217(.A1(KEYINPUT83), .A2(new_n395), .A3(new_n403), .A4(new_n400), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n399), .B1(new_n391), .B2(new_n394), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT83), .B1(new_n405), .B2(new_n403), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n405), .A2(KEYINPUT4), .A3(new_n403), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n261), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n397), .A2(G104), .ZN(new_n411));
  OAI21_X1  g225(.A(G101), .B1(new_n389), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n342), .A3(G116), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G113), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(KEYINPUT5), .B2(new_n243), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n244), .A2(new_n246), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n412), .B(new_n418), .C1(new_n404), .C2(new_n406), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n395), .A2(new_n403), .A3(new_n400), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n405), .A2(KEYINPUT83), .A3(new_n403), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n426), .A2(KEYINPUT86), .A3(new_n412), .A4(new_n418), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n410), .A2(new_n421), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G110), .B(G122), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n410), .A2(new_n421), .A3(new_n429), .A4(new_n427), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(KEYINPUT6), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n279), .A2(new_n331), .ZN(new_n434));
  INV_X1    g248(.A(new_n331), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n194), .B(new_n435), .C1(new_n255), .C2(new_n256), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n434), .A2(KEYINPUT87), .A3(new_n436), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n267), .A2(G224), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n428), .A2(new_n444), .A3(new_n430), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n433), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT92), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(KEYINPUT7), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n437), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n448), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n434), .A2(KEYINPUT92), .A3(new_n436), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n436), .A2(KEYINPUT91), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT91), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n206), .A2(new_n453), .A3(new_n435), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n454), .A3(new_n434), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n449), .A2(new_n451), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n412), .B1(new_n404), .B2(new_n406), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n418), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n415), .A2(KEYINPUT88), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n414), .A2(new_n460), .A3(G113), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n459), .A2(new_n461), .B1(KEYINPUT5), .B2(new_n243), .ZN(new_n462));
  OR3_X1    g276(.A1(new_n462), .A2(KEYINPUT89), .A3(new_n417), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT89), .B1(new_n462), .B2(new_n417), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n426), .A2(new_n465), .A3(new_n412), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n429), .B(KEYINPUT8), .ZN(new_n467));
  AND4_X1   g281(.A1(KEYINPUT90), .A2(new_n458), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n467), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n457), .B2(new_n418), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT90), .B1(new_n470), .B2(new_n466), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n432), .B(new_n456), .C1(new_n468), .C2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT93), .B1(new_n472), .B2(new_n322), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n446), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n432), .A2(new_n456), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n458), .A2(new_n466), .A3(new_n467), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n470), .A2(KEYINPUT90), .A3(new_n466), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(G902), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT93), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n383), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n433), .A2(new_n443), .A3(new_n445), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n481), .B2(KEYINPUT93), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n472), .A2(new_n322), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT93), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n383), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n382), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G469), .ZN(new_n492));
  XOR2_X1   g306(.A(G110), .B(G140), .Z(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT80), .ZN(new_n494));
  INV_X1    g308(.A(G227), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(G953), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n494), .B(new_n496), .Z(new_n497));
  AOI21_X1  g311(.A(new_n408), .B1(new_n426), .B2(new_n402), .ZN(new_n498));
  INV_X1    g312(.A(new_n457), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT10), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n206), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n498), .A2(new_n241), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n278), .A2(new_n201), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n194), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n412), .B(new_n504), .C1(new_n404), .C2(new_n406), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT84), .B1(new_n505), .B2(new_n500), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n505), .A2(KEYINPUT84), .A3(new_n500), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n232), .ZN(new_n509));
  INV_X1    g323(.A(new_n232), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n502), .B(new_n510), .C1(new_n506), .C2(new_n507), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n497), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n457), .A2(new_n206), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n513), .A2(new_n505), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n282), .A2(KEYINPUT12), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n510), .B1(new_n513), .B2(new_n505), .ZN(new_n516));
  OAI22_X1  g330(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(KEYINPUT12), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n511), .A2(new_n517), .A3(new_n497), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n492), .B(new_n322), .C1(new_n512), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n511), .A2(new_n517), .ZN(new_n520));
  INV_X1    g334(.A(new_n497), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n509), .A2(new_n511), .A3(new_n497), .ZN(new_n523));
  AOI21_X1  g337(.A(G902), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n519), .B1(new_n524), .B2(new_n492), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT9), .B(G234), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n526), .B(KEYINPUT78), .Z(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G221), .B1(new_n528), .B2(G902), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n529), .B(KEYINPUT79), .Z(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(G116), .B(G122), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n533), .A2(new_n397), .ZN(new_n534));
  INV_X1    g348(.A(G116), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G122), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n536), .A2(KEYINPUT14), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n535), .A2(G122), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n538), .B2(KEYINPUT14), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n397), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n340), .A2(G143), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n190), .A2(G128), .ZN(new_n542));
  OR3_X1    g356(.A1(new_n541), .A2(new_n542), .A3(G134), .ZN(new_n543));
  OAI21_X1  g357(.A(G134), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  AOI211_X1 g358(.A(new_n534), .B(new_n540), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT96), .ZN(new_n546));
  INV_X1    g360(.A(new_n542), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n541), .B1(new_n547), .B2(KEYINPUT13), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n541), .A2(KEYINPUT13), .ZN(new_n549));
  OAI21_X1  g363(.A(G134), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n533), .A2(new_n397), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n550), .B(new_n543), .C1(new_n534), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n527), .A2(G217), .A3(new_n267), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n546), .B2(new_n552), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT97), .B1(new_n558), .B2(G902), .ZN(new_n559));
  INV_X1    g373(.A(G478), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT97), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n563), .B(new_n322), .C1(new_n555), .C2(new_n557), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n559), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n564), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OR3_X1    g381(.A1(new_n338), .A2(KEYINPUT94), .A3(KEYINPUT19), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT94), .B1(new_n338), .B2(KEYINPUT19), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(KEYINPUT19), .B2(new_n336), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n188), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n266), .A2(new_n267), .A3(G214), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G143), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(new_n212), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n337), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(G113), .B(G122), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(new_n385), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n574), .A2(new_n212), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT18), .ZN(new_n581));
  INV_X1    g395(.A(new_n336), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n339), .B1(new_n582), .B2(new_n188), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT18), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n574), .B1(new_n584), .B2(new_n212), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n576), .A2(new_n579), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n580), .A2(KEYINPUT17), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n575), .B2(KEYINPUT17), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n586), .B1(new_n589), .B2(new_n356), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n578), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT20), .ZN(new_n593));
  NOR2_X1   g407(.A1(G475), .A2(G902), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n587), .A2(new_n591), .ZN(new_n596));
  INV_X1    g410(.A(new_n594), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT20), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n578), .A2(KEYINPUT95), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n590), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n590), .A2(new_n600), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n322), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G475), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(G234), .A2(G237), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(G952), .A3(new_n267), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(G902), .A3(G953), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT21), .B(G898), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n567), .A2(new_n606), .A3(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n491), .A2(new_n532), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n379), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  NOR2_X1   g432(.A1(new_n532), .A2(new_n378), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n302), .A2(new_n305), .B1(new_n312), .B2(new_n313), .ZN(new_n620));
  OAI21_X1  g434(.A(G472), .B1(new_n620), .B2(G902), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(KEYINPUT98), .A3(new_n323), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n623), .B(G472), .C1(new_n620), .C2(G902), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT99), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n558), .A2(G478), .A3(G902), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n553), .B(new_n554), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(KEYINPUT33), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n558), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n322), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n628), .B1(new_n633), .B2(G478), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n605), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n489), .B1(new_n485), .B2(new_n488), .ZN(new_n637));
  INV_X1    g451(.A(new_n473), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n638), .A2(new_n482), .A3(new_n383), .A4(new_n484), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT100), .B1(new_n640), .B2(new_n382), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n642));
  AOI211_X1 g456(.A(new_n642), .B(new_n381), .C1(new_n637), .C2(new_n639), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n613), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n627), .A2(new_n636), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NOR2_X1   g462(.A1(new_n567), .A2(new_n605), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n627), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NOR2_X1   g466(.A1(new_n330), .A2(KEYINPUT36), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n362), .B(new_n653), .Z(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n369), .A2(new_n373), .B1(new_n376), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n625), .A2(KEYINPUT101), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT101), .B1(new_n625), .B2(new_n657), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n616), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  INV_X1    g476(.A(new_n296), .ZN(new_n663));
  INV_X1    g477(.A(new_n325), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT32), .B1(new_n323), .B2(new_n324), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n666), .B(new_n657), .C1(new_n641), .C2(new_n643), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n522), .A2(new_n523), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n322), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(G469), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n530), .B1(new_n670), .B2(new_n519), .ZN(new_n671));
  OR3_X1    g485(.A1(new_n610), .A2(KEYINPUT102), .A3(G900), .ZN(new_n672));
  OAI21_X1  g486(.A(KEYINPUT102), .B1(new_n610), .B2(G900), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n608), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n567), .A2(new_n605), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n667), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n340), .ZN(G30));
  NAND2_X1  g493(.A1(new_n316), .A2(new_n325), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n264), .A2(new_n294), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(G472), .A3(new_n300), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n187), .A2(new_n322), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT103), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n567), .A2(new_n606), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(new_n382), .A3(new_n656), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n640), .B(KEYINPUT38), .Z(new_n690));
  OR2_X1    g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(KEYINPUT104), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(KEYINPUT104), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n674), .B(KEYINPUT39), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n671), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT40), .Z(new_n696));
  NAND3_X1  g510(.A1(new_n692), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT105), .B(G143), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G45));
  INV_X1    g513(.A(new_n628), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n629), .A2(KEYINPUT33), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n558), .A2(new_n631), .ZN(new_n702));
  AOI21_X1  g516(.A(G902), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n700), .B1(new_n703), .B2(new_n560), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n704), .A2(new_n606), .A3(new_n675), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n671), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n667), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n188), .ZN(G48));
  OAI21_X1  g522(.A(new_n322), .B1(new_n512), .B2(new_n518), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n531), .A3(new_n519), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n326), .A2(new_n378), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n491), .A2(new_n642), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n381), .B1(new_n637), .B2(new_n639), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT100), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n712), .A2(new_n716), .A3(new_n614), .A4(new_n636), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  OAI211_X1 g533(.A(new_n614), .B(new_n649), .C1(new_n641), .C2(new_n643), .ZN(new_n720));
  AOI22_X1  g534(.A1(new_n369), .A2(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n721));
  INV_X1    g535(.A(new_n711), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n666), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n535), .ZN(G18));
  OR2_X1    g539(.A1(new_n326), .A2(new_n615), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n716), .B2(new_n722), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n728), .B(new_n722), .C1(new_n641), .C2(new_n643), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n657), .B(new_n727), .C1(new_n729), .C2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  INV_X1    g547(.A(new_n294), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n306), .B1(new_n734), .B2(new_n265), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n187), .A3(new_n322), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT107), .B(G472), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n620), .B2(G902), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n721), .A2(new_n736), .A3(new_n614), .A4(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n711), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(new_n688), .C1(new_n641), .C2(new_n643), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  INV_X1    g557(.A(new_n705), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n736), .A2(new_n739), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n657), .B(new_n746), .C1(new_n729), .C2(new_n731), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  AOI21_X1  g562(.A(new_n296), .B1(new_n323), .B2(new_n297), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n315), .A2(KEYINPUT32), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n378), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n637), .A2(new_n382), .A3(new_n639), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n671), .A3(new_n705), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT42), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n637), .A2(new_n382), .A3(new_n639), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n532), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n635), .A2(KEYINPUT42), .A3(new_n675), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n666), .A3(new_n757), .A4(new_n721), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  NAND4_X1  g574(.A1(new_n756), .A2(new_n666), .A3(new_n721), .A4(new_n676), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  XNOR2_X1  g576(.A(new_n605), .B(KEYINPUT108), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(KEYINPUT43), .A3(new_n634), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n763), .A2(new_n766), .A3(KEYINPUT43), .A4(new_n634), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n704), .A2(new_n605), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n765), .B(new_n767), .C1(KEYINPUT43), .C2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(new_n657), .ZN(new_n770));
  INV_X1    g584(.A(new_n625), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(KEYINPUT44), .A3(new_n771), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n775));
  OAI221_X1 g589(.A(new_n752), .B1(KEYINPUT44), .B2(new_n772), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n668), .B(KEYINPUT45), .Z(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n492), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(G469), .B2(G902), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT46), .ZN(new_n780));
  INV_X1    g594(.A(new_n519), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n779), .B2(KEYINPUT46), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n530), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n694), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n776), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n207), .ZN(G39));
  OR2_X1    g600(.A1(new_n783), .A2(KEYINPUT47), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n783), .A2(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n666), .A2(new_n744), .A3(new_n721), .A4(new_n755), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NOR2_X1   g606(.A1(new_n745), .A2(new_n656), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n711), .A2(new_n755), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n769), .A2(new_n609), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n687), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n721), .A2(new_n800), .A3(new_n794), .A4(new_n609), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n606), .A3(new_n704), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n769), .A2(new_n609), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n378), .A3(new_n745), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n381), .A3(new_n690), .A4(new_n722), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n799), .B(new_n802), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n710), .A2(new_n519), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n530), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n787), .A2(new_n788), .A3(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n804), .A2(new_n752), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n809), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n814), .B2(KEYINPUT116), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n815), .B(KEYINPUT51), .C1(new_n814), .C2(KEYINPUT116), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n804), .B1(new_n731), .B2(new_n729), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n801), .A2(new_n636), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(G952), .A3(new_n267), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n751), .B1(new_n797), .B2(new_n798), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT48), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT120), .Z(new_n825));
  NOR2_X1   g639(.A1(new_n823), .A2(KEYINPUT48), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT119), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n822), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n818), .A2(new_n819), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n667), .B1(new_n677), .B2(new_n706), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n644), .A2(new_n606), .A3(new_n567), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n532), .A2(new_n657), .A3(new_n675), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n687), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n747), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n722), .B1(new_n641), .B2(new_n643), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT106), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n656), .B1(new_n841), .B2(new_n730), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n830), .B1(new_n842), .B2(new_n746), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .A3(new_n834), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n837), .A2(new_n839), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n614), .B(new_n636), .C1(new_n641), .C2(new_n643), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n742), .B1(new_n847), .B2(new_n723), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n724), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n567), .B2(new_n605), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n606), .A2(new_n565), .A3(KEYINPUT111), .A4(new_n566), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n613), .B1(new_n853), .B2(new_n635), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n714), .A3(new_n619), .A4(new_n625), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n660), .A2(new_n617), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n732), .A2(new_n849), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n675), .B(new_n605), .C1(new_n566), .C2(new_n565), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n666), .A2(new_n657), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n756), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n326), .A2(new_n656), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(KEYINPUT112), .A3(new_n756), .A4(new_n859), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n756), .A2(new_n705), .A3(new_n793), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n759), .A3(new_n761), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n857), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n835), .A2(new_n838), .A3(new_n836), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n845), .A2(new_n846), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT52), .B1(new_n843), .B2(new_n834), .ZN(new_n871));
  AND4_X1   g685(.A1(KEYINPUT52), .A2(new_n747), .A3(new_n831), .A4(new_n834), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT53), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n874), .A3(KEYINPUT54), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n656), .B(new_n726), .C1(new_n841), .C2(new_n730), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n712), .A2(new_n716), .A3(new_n614), .A4(new_n649), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n717), .A2(new_n878), .A3(new_n742), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n876), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n732), .A2(new_n849), .A3(KEYINPUT115), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n862), .A2(new_n864), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n660), .A2(new_n617), .A3(KEYINPUT53), .A4(new_n855), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n754), .A2(new_n758), .A3(new_n761), .A4(new_n866), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n880), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n845), .A2(new_n886), .A3(new_n869), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n884), .B1(new_n862), .B2(new_n864), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n732), .A3(new_n856), .A4(new_n849), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n837), .B2(new_n844), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n890), .A2(KEYINPUT114), .A3(KEYINPUT53), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT114), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n873), .B2(new_n846), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n887), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n875), .B1(new_n894), .B2(KEYINPUT54), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n829), .A2(new_n895), .B1(G952), .B2(G953), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n810), .B(KEYINPUT49), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n530), .A2(new_n381), .ZN(new_n898));
  AND4_X1   g712(.A1(new_n721), .A2(new_n763), .A3(new_n634), .A4(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n897), .A2(new_n690), .A3(new_n800), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n896), .A2(new_n900), .ZN(G75));
  NOR2_X1   g715(.A1(new_n267), .A2(G952), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n845), .A2(new_n886), .A3(new_n869), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n873), .A2(new_n892), .A3(new_n846), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT114), .B1(new_n890), .B2(KEYINPUT53), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n322), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT56), .B1(new_n908), .B2(new_n489), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n433), .A2(new_n445), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n443), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n446), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n903), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n907), .B2(new_n322), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n894), .A2(KEYINPUT121), .A3(G902), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n489), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n914), .B1(new_n918), .B2(new_n920), .ZN(G51));
  AND3_X1   g735(.A1(new_n916), .A2(new_n778), .A3(new_n917), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n512), .A2(new_n518), .ZN(new_n923));
  NAND2_X1  g737(.A1(G469), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT57), .Z(new_n925));
  NOR2_X1   g739(.A1(new_n894), .A2(KEYINPUT54), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT54), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n906), .A2(new_n905), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n887), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n925), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n922), .A2(KEYINPUT122), .B1(new_n923), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n916), .A2(new_n778), .A3(new_n917), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n902), .B1(new_n931), .B2(new_n934), .ZN(G54));
  AND2_X1   g749(.A1(KEYINPUT58), .A2(G475), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n916), .A2(new_n917), .A3(new_n936), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n937), .A2(KEYINPUT123), .A3(new_n596), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT123), .B1(new_n937), .B2(new_n596), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n916), .A2(new_n917), .A3(new_n592), .A4(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n903), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(G60));
  NOR2_X1   g756(.A1(new_n630), .A2(new_n632), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT59), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n944), .B1(new_n895), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n926), .A2(new_n929), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n944), .A2(new_n946), .ZN(new_n949));
  AOI211_X1 g763(.A(new_n902), .B(new_n947), .C1(new_n948), .C2(new_n949), .ZN(G63));
  XOR2_X1   g764(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n951));
  OAI21_X1  g765(.A(KEYINPUT60), .B1(new_n370), .B2(new_n322), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n370), .A2(new_n322), .A3(KEYINPUT60), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n894), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n903), .B1(new_n954), .B2(new_n375), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n894), .A2(new_n952), .A3(new_n953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n654), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n951), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n957), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n366), .A3(new_n365), .ZN(new_n960));
  INV_X1    g774(.A(new_n951), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n959), .A2(new_n903), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n958), .A2(new_n962), .ZN(G66));
  NAND2_X1  g777(.A1(G224), .A2(G953), .ZN(new_n964));
  OAI22_X1  g778(.A1(new_n857), .A2(G953), .B1(new_n612), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(G898), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n910), .B1(new_n966), .B2(G953), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  INV_X1    g782(.A(new_n785), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n697), .A2(new_n843), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n695), .B1(new_n635), .B2(new_n853), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n379), .A3(new_n752), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n969), .A2(new_n972), .A3(new_n791), .A4(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(new_n267), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n303), .B(new_n571), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(G900), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n495), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT125), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n759), .A2(new_n761), .ZN(new_n984));
  AND4_X1   g798(.A1(new_n694), .A2(new_n783), .A3(new_n832), .A4(new_n751), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n785), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n791), .A3(new_n843), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n267), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n980), .A2(G953), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n977), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n979), .B(new_n983), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n988), .B2(new_n989), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n982), .B1(new_n993), .B2(new_n978), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(G72));
  XNOR2_X1  g809(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n684), .B(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n987), .B2(new_n857), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n286), .A2(new_n287), .A3(new_n271), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n997), .B1(new_n300), .B2(new_n288), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n870), .A2(new_n874), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1001), .A2(new_n903), .A3(new_n1003), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n975), .A2(new_n857), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(KEYINPUT127), .A3(new_n998), .ZN(new_n1006));
  AOI21_X1  g820(.A(KEYINPUT127), .B1(new_n1005), .B2(new_n998), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n271), .B1(new_n286), .B2(new_n287), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1004), .B1(new_n1006), .B2(new_n1009), .ZN(G57));
endmodule


