

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X2 U325 ( .A(n512), .B(KEYINPUT38), .ZN(n518) );
  INV_X1 U326 ( .A(n386), .ZN(n478) );
  NOR2_X1 U327 ( .A1(n586), .A2(n418), .ZN(n419) );
  XOR2_X1 U328 ( .A(G141GAT), .B(G22GAT), .Z(n428) );
  XOR2_X1 U329 ( .A(G162GAT), .B(G50GAT), .Z(n328) );
  XNOR2_X1 U330 ( .A(n395), .B(KEYINPUT99), .ZN(n496) );
  XNOR2_X1 U331 ( .A(n444), .B(n443), .ZN(n445) );
  NOR2_X1 U332 ( .A1(n385), .A2(n573), .ZN(n552) );
  XNOR2_X1 U333 ( .A(n473), .B(n472), .ZN(n551) );
  XNOR2_X1 U334 ( .A(n376), .B(n335), .ZN(n336) );
  XOR2_X1 U335 ( .A(n367), .B(n366), .Z(n554) );
  AND2_X1 U336 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U337 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n443) );
  INV_X1 U338 ( .A(n449), .ZN(n450) );
  XNOR2_X1 U339 ( .A(n363), .B(n293), .ZN(n335) );
  XNOR2_X1 U340 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U341 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n472) );
  XNOR2_X1 U342 ( .A(n453), .B(n452), .ZN(n455) );
  NOR2_X1 U343 ( .A1(n481), .A2(n541), .ZN(n570) );
  INV_X1 U344 ( .A(G106GAT), .ZN(n457) );
  XNOR2_X1 U345 ( .A(n347), .B(n346), .ZN(n541) );
  XNOR2_X1 U346 ( .A(n489), .B(G190GAT), .ZN(n490) );
  XNOR2_X1 U347 ( .A(n457), .B(KEYINPUT44), .ZN(n458) );
  XNOR2_X1 U348 ( .A(n491), .B(n490), .ZN(G1351GAT) );
  XOR2_X1 U349 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n295) );
  XNOR2_X1 U350 ( .A(G204GAT), .B(KEYINPUT22), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U352 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n297) );
  XNOR2_X1 U353 ( .A(n328), .B(n428), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U355 ( .A(n299), .B(n298), .Z(n301) );
  NAND2_X1 U356 ( .A1(G228GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U358 ( .A(n302), .B(KEYINPUT89), .Z(n305) );
  XNOR2_X1 U359 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n303), .B(KEYINPUT2), .ZN(n362) );
  XNOR2_X1 U361 ( .A(n362), .B(KEYINPUT90), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n315) );
  XOR2_X1 U363 ( .A(G197GAT), .B(KEYINPUT21), .Z(n307) );
  XNOR2_X1 U364 ( .A(G218GAT), .B(G211GAT), .ZN(n306) );
  XNOR2_X1 U365 ( .A(n307), .B(n306), .ZN(n373) );
  INV_X1 U366 ( .A(G78GAT), .ZN(n308) );
  NAND2_X1 U367 ( .A1(n308), .A2(KEYINPUT72), .ZN(n311) );
  INV_X1 U368 ( .A(KEYINPUT72), .ZN(n309) );
  NAND2_X1 U369 ( .A1(n309), .A2(G78GAT), .ZN(n310) );
  NAND2_X1 U370 ( .A1(n311), .A2(n310), .ZN(n313) );
  XNOR2_X1 U371 ( .A(G148GAT), .B(G106GAT), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n313), .B(n312), .ZN(n444) );
  XOR2_X1 U373 ( .A(n373), .B(n444), .Z(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n386) );
  XNOR2_X1 U375 ( .A(KEYINPUT28), .B(n386), .ZN(n530) );
  INV_X1 U376 ( .A(KEYINPUT37), .ZN(n420) );
  XOR2_X1 U377 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n317) );
  NAND2_X1 U378 ( .A1(G232GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U380 ( .A(n318), .B(KEYINPUT9), .Z(n323) );
  XOR2_X1 U381 ( .A(G43GAT), .B(KEYINPUT8), .Z(n320) );
  XNOR2_X1 U382 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n427) );
  XNOR2_X1 U384 ( .A(G36GAT), .B(KEYINPUT74), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n321), .B(G190GAT), .ZN(n379) );
  XNOR2_X1 U386 ( .A(n427), .B(n379), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U388 ( .A(G92GAT), .B(G106GAT), .Z(n325) );
  XNOR2_X1 U389 ( .A(G134GAT), .B(G218GAT), .ZN(n324) );
  XNOR2_X1 U390 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U391 ( .A(n327), .B(n326), .Z(n330) );
  XOR2_X1 U392 ( .A(G85GAT), .B(G99GAT), .Z(n449) );
  XNOR2_X1 U393 ( .A(n328), .B(n449), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n330), .B(n329), .ZN(n492) );
  XNOR2_X1 U395 ( .A(KEYINPUT36), .B(n492), .ZN(n586) );
  XOR2_X1 U396 ( .A(G120GAT), .B(G71GAT), .Z(n441) );
  XOR2_X1 U397 ( .A(G127GAT), .B(G15GAT), .Z(n407) );
  XOR2_X1 U398 ( .A(n441), .B(n407), .Z(n332) );
  XNOR2_X1 U399 ( .A(G43GAT), .B(G190GAT), .ZN(n331) );
  XNOR2_X1 U400 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U401 ( .A(G169GAT), .B(KEYINPUT19), .Z(n334) );
  XNOR2_X1 U402 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n333) );
  XNOR2_X1 U403 ( .A(n334), .B(n333), .ZN(n376) );
  XOR2_X1 U404 ( .A(G134GAT), .B(KEYINPUT0), .Z(n363) );
  XOR2_X1 U405 ( .A(n337), .B(n336), .Z(n339) );
  XNOR2_X1 U406 ( .A(G99GAT), .B(G183GAT), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n347) );
  XOR2_X1 U408 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n341) );
  XNOR2_X1 U409 ( .A(G176GAT), .B(KEYINPUT86), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U411 ( .A(KEYINPUT82), .B(KEYINPUT84), .Z(n343) );
  XNOR2_X1 U412 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n342) );
  XNOR2_X1 U413 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U414 ( .A(n345), .B(n344), .Z(n346) );
  XOR2_X1 U415 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n349) );
  XNOR2_X1 U416 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n348) );
  XNOR2_X1 U417 ( .A(n349), .B(n348), .ZN(n367) );
  XOR2_X1 U418 ( .A(G120GAT), .B(G85GAT), .Z(n351) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(G162GAT), .ZN(n350) );
  XNOR2_X1 U420 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U421 ( .A(G57GAT), .B(G148GAT), .Z(n353) );
  XNOR2_X1 U422 ( .A(G127GAT), .B(G141GAT), .ZN(n352) );
  XNOR2_X1 U423 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U424 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U425 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n357) );
  NAND2_X1 U426 ( .A1(G225GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U427 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U428 ( .A(KEYINPUT5), .B(n358), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U430 ( .A(G113GAT), .B(G1GAT), .Z(n424) );
  XOR2_X1 U431 ( .A(n361), .B(n424), .Z(n365) );
  XNOR2_X1 U432 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U434 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n369) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U437 ( .A(n370), .B(KEYINPUT95), .Z(n375) );
  XOR2_X1 U438 ( .A(G204GAT), .B(G176GAT), .Z(n372) );
  XNOR2_X1 U439 ( .A(G92GAT), .B(G64GAT), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n372), .B(n371), .ZN(n447) );
  XNOR2_X1 U441 ( .A(n373), .B(n447), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U443 ( .A(n377), .B(n376), .Z(n381) );
  XNOR2_X1 U444 ( .A(G183GAT), .B(G8GAT), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n378), .B(KEYINPUT75), .ZN(n408) );
  XNOR2_X1 U446 ( .A(n379), .B(n408), .ZN(n380) );
  XOR2_X1 U447 ( .A(n381), .B(n380), .Z(n535) );
  XNOR2_X1 U448 ( .A(n535), .B(KEYINPUT27), .ZN(n385) );
  INV_X1 U449 ( .A(n385), .ZN(n382) );
  NAND2_X1 U450 ( .A1(n530), .A2(n382), .ZN(n383) );
  NOR2_X1 U451 ( .A1(n554), .A2(n383), .ZN(n539) );
  NAND2_X1 U452 ( .A1(n541), .A2(n539), .ZN(n394) );
  NAND2_X1 U453 ( .A1(n541), .A2(n478), .ZN(n384) );
  XNOR2_X1 U454 ( .A(n384), .B(KEYINPUT26), .ZN(n573) );
  XNOR2_X1 U455 ( .A(n552), .B(KEYINPUT97), .ZN(n391) );
  XOR2_X1 U456 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n389) );
  OR2_X1 U457 ( .A1(n541), .A2(n535), .ZN(n387) );
  NAND2_X1 U458 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n389), .B(n388), .ZN(n390) );
  NAND2_X1 U460 ( .A1(n391), .A2(n390), .ZN(n392) );
  NAND2_X1 U461 ( .A1(n392), .A2(n554), .ZN(n393) );
  NAND2_X1 U462 ( .A1(n394), .A2(n393), .ZN(n395) );
  XOR2_X1 U463 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n397) );
  XNOR2_X1 U464 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n416) );
  XOR2_X1 U466 ( .A(G78GAT), .B(G211GAT), .Z(n399) );
  XNOR2_X1 U467 ( .A(G1GAT), .B(G22GAT), .ZN(n398) );
  XNOR2_X1 U468 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U469 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n401) );
  XNOR2_X1 U470 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n400) );
  XNOR2_X1 U471 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U472 ( .A(n403), .B(n402), .Z(n414) );
  XNOR2_X1 U473 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n404), .B(KEYINPUT13), .ZN(n448) );
  XOR2_X1 U475 ( .A(n448), .B(KEYINPUT79), .Z(n406) );
  NAND2_X1 U476 ( .A1(G231GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n406), .B(n405), .ZN(n412) );
  XOR2_X1 U478 ( .A(n408), .B(n407), .Z(n410) );
  XNOR2_X1 U479 ( .A(G155GAT), .B(G71GAT), .ZN(n409) );
  XNOR2_X1 U480 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U481 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U482 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n416), .B(n415), .ZN(n582) );
  NOR2_X1 U484 ( .A1(n496), .A2(n582), .ZN(n417) );
  XNOR2_X1 U485 ( .A(KEYINPUT105), .B(n417), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n420), .B(n419), .ZN(n510) );
  XOR2_X1 U487 ( .A(G197GAT), .B(G169GAT), .Z(n422) );
  XNOR2_X1 U488 ( .A(G15GAT), .B(G8GAT), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U490 ( .A(n423), .B(G36GAT), .Z(n426) );
  XNOR2_X1 U491 ( .A(n424), .B(G50GAT), .ZN(n425) );
  XNOR2_X1 U492 ( .A(n426), .B(n425), .ZN(n432) );
  XOR2_X1 U493 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U494 ( .A1(G229GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U495 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U496 ( .A(n432), .B(n431), .Z(n440) );
  XOR2_X1 U497 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n434) );
  XNOR2_X1 U498 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n433) );
  XNOR2_X1 U499 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U500 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n436) );
  XNOR2_X1 U501 ( .A(KEYINPUT65), .B(KEYINPUT66), .ZN(n435) );
  XNOR2_X1 U502 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U503 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n497) );
  INV_X1 U505 ( .A(n497), .ZN(n574) );
  XNOR2_X1 U506 ( .A(n441), .B(KEYINPUT32), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n442), .B(KEYINPUT73), .ZN(n446) );
  XOR2_X1 U508 ( .A(n446), .B(n445), .Z(n453) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n451) );
  NAND2_X1 U510 ( .A1(G230GAT), .A2(G233GAT), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n455), .B(n454), .ZN(n578) );
  XNOR2_X1 U512 ( .A(n578), .B(KEYINPUT41), .ZN(n485) );
  NOR2_X1 U513 ( .A1(n574), .A2(n485), .ZN(n523) );
  NAND2_X1 U514 ( .A1(n510), .A2(n523), .ZN(n456) );
  XNOR2_X1 U515 ( .A(KEYINPUT110), .B(n456), .ZN(n537) );
  NOR2_X1 U516 ( .A1(n530), .A2(n537), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(G1339GAT) );
  XOR2_X1 U518 ( .A(n535), .B(KEYINPUT120), .Z(n474) );
  NOR2_X1 U519 ( .A1(n497), .A2(n485), .ZN(n461) );
  XNOR2_X1 U520 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n461), .B(n460), .ZN(n463) );
  INV_X1 U522 ( .A(n492), .ZN(n566) );
  NOR2_X1 U523 ( .A1(n582), .A2(n566), .ZN(n462) );
  AND2_X1 U524 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U525 ( .A(n464), .B(KEYINPUT47), .ZN(n471) );
  INV_X1 U526 ( .A(n582), .ZN(n465) );
  NOR2_X1 U527 ( .A1(n465), .A2(n586), .ZN(n466) );
  XOR2_X1 U528 ( .A(KEYINPUT45), .B(n466), .Z(n467) );
  NOR2_X1 U529 ( .A1(n578), .A2(n467), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT112), .B(n468), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n469), .A2(n497), .ZN(n470) );
  NAND2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n474), .A2(n551), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT121), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(KEYINPUT54), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n477), .A2(n554), .ZN(n572) );
  NOR2_X1 U537 ( .A1(n478), .A2(n572), .ZN(n480) );
  XNOR2_X1 U538 ( .A(KEYINPUT122), .B(KEYINPUT55), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U540 ( .A1(n570), .A2(n574), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n482) );
  XNOR2_X1 U542 ( .A(n482), .B(G169GAT), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(G1348GAT) );
  INV_X1 U544 ( .A(n485), .ZN(n561) );
  NAND2_X1 U545 ( .A1(n570), .A2(n561), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n486) );
  XNOR2_X1 U547 ( .A(n486), .B(G176GAT), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1349GAT) );
  NAND2_X1 U549 ( .A1(n570), .A2(n566), .ZN(n491) );
  XOR2_X1 U550 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n500) );
  XOR2_X1 U552 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n494) );
  NAND2_X1 U553 ( .A1(n492), .A2(n582), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(n495) );
  NOR2_X1 U555 ( .A1(n496), .A2(n495), .ZN(n522) );
  NOR2_X1 U556 ( .A1(n497), .A2(n578), .ZN(n511) );
  NAND2_X1 U557 ( .A1(n522), .A2(n511), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(KEYINPUT100), .ZN(n508) );
  NOR2_X1 U559 ( .A1(n554), .A2(n508), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NOR2_X1 U562 ( .A1(n508), .A2(n535), .ZN(n502) );
  XOR2_X1 U563 ( .A(KEYINPUT102), .B(n502), .Z(n503) );
  XNOR2_X1 U564 ( .A(G8GAT), .B(n503), .ZN(G1325GAT) );
  NOR2_X1 U565 ( .A1(n541), .A2(n508), .ZN(n507) );
  XOR2_X1 U566 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n505) );
  XNOR2_X1 U567 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1326GAT) );
  NOR2_X1 U570 ( .A1(n530), .A2(n508), .ZN(n509) );
  XOR2_X1 U571 ( .A(G22GAT), .B(n509), .Z(G1327GAT) );
  NAND2_X1 U572 ( .A1(n511), .A2(n510), .ZN(n512) );
  NOR2_X1 U573 ( .A1(n518), .A2(n554), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n513), .B(KEYINPUT39), .ZN(n514) );
  XNOR2_X1 U575 ( .A(G29GAT), .B(n514), .ZN(G1328GAT) );
  NOR2_X1 U576 ( .A1(n518), .A2(n535), .ZN(n515) );
  XOR2_X1 U577 ( .A(G36GAT), .B(n515), .Z(G1329GAT) );
  NOR2_X1 U578 ( .A1(n518), .A2(n541), .ZN(n516) );
  XOR2_X1 U579 ( .A(KEYINPUT40), .B(n516), .Z(n517) );
  XNOR2_X1 U580 ( .A(G43GAT), .B(n517), .ZN(G1330GAT) );
  NOR2_X1 U581 ( .A1(n530), .A2(n518), .ZN(n519) );
  XOR2_X1 U582 ( .A(G50GAT), .B(n519), .Z(G1331GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n521) );
  XNOR2_X1 U584 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(n525) );
  NAND2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n529) );
  NOR2_X1 U587 ( .A1(n554), .A2(n529), .ZN(n524) );
  XOR2_X1 U588 ( .A(n525), .B(n524), .Z(G1332GAT) );
  NOR2_X1 U589 ( .A1(n535), .A2(n529), .ZN(n526) );
  XOR2_X1 U590 ( .A(KEYINPUT108), .B(n526), .Z(n527) );
  XNOR2_X1 U591 ( .A(G64GAT), .B(n527), .ZN(G1333GAT) );
  NOR2_X1 U592 ( .A1(n541), .A2(n529), .ZN(n528) );
  XOR2_X1 U593 ( .A(G71GAT), .B(n528), .Z(G1334GAT) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U595 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U597 ( .A(G78GAT), .B(n533), .Z(G1335GAT) );
  NOR2_X1 U598 ( .A1(n554), .A2(n537), .ZN(n534) );
  XOR2_X1 U599 ( .A(G85GAT), .B(n534), .Z(G1336GAT) );
  NOR2_X1 U600 ( .A1(n537), .A2(n535), .ZN(n536) );
  XOR2_X1 U601 ( .A(G92GAT), .B(n536), .Z(G1337GAT) );
  NOR2_X1 U602 ( .A1(n537), .A2(n541), .ZN(n538) );
  XOR2_X1 U603 ( .A(G99GAT), .B(n538), .Z(G1338GAT) );
  NAND2_X1 U604 ( .A1(n539), .A2(n551), .ZN(n540) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n574), .A2(n548), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n544) );
  NAND2_X1 U609 ( .A1(n548), .A2(n561), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(G120GAT), .B(n545), .Z(G1341GAT) );
  NAND2_X1 U612 ( .A1(n582), .A2(n548), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U616 ( .A1(n548), .A2(n566), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n556) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n567) );
  NAND2_X1 U621 ( .A1(n567), .A2(n574), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G141GAT), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n559) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT52), .B(n560), .Z(n563) );
  NAND2_X1 U628 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n582), .A2(n567), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT118), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G155GAT), .B(n565), .ZN(G1346GAT) );
  XOR2_X1 U633 ( .A(G162GAT), .B(KEYINPUT119), .Z(n569) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n582), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n584) );
  NAND2_X1 U640 ( .A1(n584), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n580) );
  NAND2_X1 U644 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n584), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U649 ( .A(n584), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

