

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808;

  OR2_X1 U381 ( .A1(n628), .A2(n758), .ZN(n617) );
  INV_X1 U382 ( .A(G902), .ZN(n507) );
  INV_X2 U383 ( .A(G953), .ZN(n796) );
  XNOR2_X2 U384 ( .A(n546), .B(n545), .ZN(n608) );
  NOR2_X2 U385 ( .A1(n568), .A2(n487), .ZN(n488) );
  XNOR2_X2 U386 ( .A(n459), .B(KEYINPUT0), .ZN(n568) );
  NOR2_X2 U387 ( .A1(n565), .A2(n610), .ZN(n554) );
  XNOR2_X1 U388 ( .A(n391), .B(n365), .ZN(n399) );
  INV_X1 U389 ( .A(KEYINPUT67), .ZN(n419) );
  XNOR2_X1 U390 ( .A(n606), .B(KEYINPUT45), .ZN(n657) );
  NOR2_X1 U391 ( .A1(n605), .A2(n604), .ZN(n606) );
  AND2_X1 U392 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U393 ( .A1(n399), .A2(n398), .ZN(n390) );
  BUF_X1 U394 ( .A(n565), .Z(n375) );
  XNOR2_X1 U395 ( .A(n482), .B(n481), .ZN(n571) );
  XNOR2_X1 U396 ( .A(n508), .B(G469), .ZN(n532) );
  XNOR2_X1 U397 ( .A(n480), .B(n392), .ZN(n771) );
  XNOR2_X1 U398 ( .A(n501), .B(n787), .ZN(n430) );
  XNOR2_X1 U399 ( .A(n410), .B(n409), .ZN(n509) );
  XNOR2_X1 U400 ( .A(n389), .B(KEYINPUT69), .ZN(n403) );
  XNOR2_X1 U401 ( .A(n417), .B(G146), .ZN(n466) );
  XOR2_X1 U402 ( .A(KEYINPUT67), .B(G101), .Z(n389) );
  XNOR2_X1 U403 ( .A(G116), .B(G113), .ZN(n401) );
  XNOR2_X1 U404 ( .A(G110), .B(G104), .ZN(n402) );
  XNOR2_X1 U405 ( .A(KEYINPUT15), .B(G902), .ZN(n544) );
  NAND2_X1 U406 ( .A1(n358), .A2(KEYINPUT2), .ZN(n668) );
  OR2_X2 U407 ( .A1(n657), .A2(n792), .ZN(n358) );
  NOR2_X1 U408 ( .A1(n568), .A2(n487), .ZN(n359) );
  OR2_X1 U409 ( .A1(n657), .A2(n792), .ZN(n360) );
  BUF_X1 U410 ( .A(n568), .Z(n569) );
  XNOR2_X1 U411 ( .A(n466), .B(n416), .ZN(n520) );
  INV_X1 U412 ( .A(KEYINPUT10), .ZN(n416) );
  OR2_X1 U413 ( .A1(n607), .A2(n552), .ZN(n487) );
  NOR2_X1 U414 ( .A1(n571), .A2(n581), .ZN(n397) );
  NOR2_X1 U415 ( .A1(G953), .A2(G237), .ZN(n492) );
  XNOR2_X1 U416 ( .A(KEYINPUT18), .B(KEYINPUT89), .ZN(n422) );
  XOR2_X1 U417 ( .A(G137), .B(G140), .Z(n519) );
  XNOR2_X1 U418 ( .A(n529), .B(KEYINPUT30), .ZN(n530) );
  INV_X1 U419 ( .A(KEYINPUT8), .ZN(n409) );
  NAND2_X1 U420 ( .A1(n796), .A2(G234), .ZN(n410) );
  XNOR2_X1 U421 ( .A(G107), .B(G116), .ZN(n476) );
  INV_X1 U422 ( .A(KEYINPUT9), .ZN(n394) );
  XNOR2_X1 U423 ( .A(G122), .B(KEYINPUT7), .ZN(n473) );
  XNOR2_X1 U424 ( .A(n470), .B(n471), .ZN(n689) );
  INV_X1 U425 ( .A(n519), .ZN(n503) );
  XNOR2_X1 U426 ( .A(n525), .B(n361), .ZN(n411) );
  NOR2_X1 U427 ( .A1(n771), .A2(G902), .ZN(n482) );
  INV_X1 U428 ( .A(G237), .ZN(n431) );
  AND2_X1 U429 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U430 ( .A(G104), .B(G113), .ZN(n463) );
  INV_X1 U431 ( .A(G131), .ZN(n462) );
  XNOR2_X1 U432 ( .A(G140), .B(G122), .ZN(n467) );
  XOR2_X1 U433 ( .A(KEYINPUT11), .B(G143), .Z(n468) );
  XOR2_X1 U434 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n461) );
  INV_X1 U435 ( .A(G125), .ZN(n417) );
  XNOR2_X1 U436 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n423) );
  XNOR2_X1 U437 ( .A(KEYINPUT76), .B(KEYINPUT91), .ZN(n512) );
  NAND2_X1 U438 ( .A1(G237), .A2(G234), .ZN(n456) );
  INV_X1 U439 ( .A(KEYINPUT112), .ZN(n408) );
  INV_X1 U440 ( .A(KEYINPUT109), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U442 ( .A(n472), .B(n414), .ZN(n413) );
  OR2_X1 U443 ( .A1(n689), .A2(G902), .ZN(n415) );
  INV_X1 U444 ( .A(G475), .ZN(n414) );
  XNOR2_X1 U445 ( .A(KEYINPUT95), .B(n533), .ZN(n587) );
  XNOR2_X1 U446 ( .A(n475), .B(n393), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U448 ( .A(n476), .B(n394), .ZN(n393) );
  XOR2_X1 U449 ( .A(KEYINPUT59), .B(n689), .Z(n690) );
  XNOR2_X1 U450 ( .A(n501), .B(n504), .ZN(n506) );
  XNOR2_X1 U451 ( .A(n503), .B(n502), .ZN(n504) );
  AND2_X1 U452 ( .A1(n678), .A2(G953), .ZN(n775) );
  NOR2_X1 U453 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U454 ( .A1(n591), .A2(n592), .ZN(n593) );
  XOR2_X1 U455 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n361) );
  OR2_X1 U456 ( .A1(n446), .A2(n445), .ZN(n362) );
  XOR2_X1 U457 ( .A(KEYINPUT4), .B(G131), .Z(n363) );
  XOR2_X1 U458 ( .A(KEYINPUT71), .B(KEYINPUT22), .Z(n364) );
  XOR2_X1 U459 ( .A(n563), .B(KEYINPUT32), .Z(n365) );
  XOR2_X1 U460 ( .A(KEYINPUT86), .B(KEYINPUT36), .Z(n366) );
  AND2_X1 U461 ( .A1(n574), .A2(KEYINPUT68), .ZN(n367) );
  XNOR2_X1 U462 ( .A(n521), .B(n794), .ZN(n695) );
  NAND2_X1 U463 ( .A1(n683), .A2(n507), .ZN(n368) );
  AND2_X1 U464 ( .A1(n561), .A2(n553), .ZN(n369) );
  XNOR2_X1 U465 ( .A(n584), .B(n551), .ZN(n565) );
  XNOR2_X1 U466 ( .A(n368), .B(n498), .ZN(n370) );
  XNOR2_X1 U467 ( .A(n499), .B(n498), .ZN(n584) );
  XNOR2_X1 U468 ( .A(n547), .B(KEYINPUT38), .ZN(n740) );
  OR2_X2 U469 ( .A1(n695), .A2(G902), .ZN(n412) );
  NOR2_X1 U470 ( .A1(n601), .A2(n373), .ZN(n371) );
  NOR2_X1 U471 ( .A1(n371), .A2(n372), .ZN(n384) );
  AND2_X1 U472 ( .A1(KEYINPUT44), .A2(n805), .ZN(n372) );
  OR2_X1 U473 ( .A1(KEYINPUT65), .A2(n574), .ZN(n373) );
  NOR2_X1 U474 ( .A1(n595), .A2(n594), .ZN(n374) );
  XNOR2_X1 U475 ( .A(n359), .B(n364), .ZN(n376) );
  XNOR2_X1 U476 ( .A(n488), .B(n364), .ZN(n560) );
  XNOR2_X1 U477 ( .A(KEYINPUT34), .B(n570), .ZN(n377) );
  XNOR2_X1 U478 ( .A(KEYINPUT42), .B(n617), .ZN(n378) );
  XNOR2_X1 U479 ( .A(KEYINPUT42), .B(n617), .ZN(n808) );
  AND2_X1 U480 ( .A1(n376), .A2(n375), .ZN(n591) );
  XNOR2_X1 U481 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X2 U482 ( .A(n624), .B(n623), .ZN(n806) );
  XNOR2_X1 U483 ( .A(n614), .B(n379), .ZN(n616) );
  XNOR2_X1 U484 ( .A(n396), .B(n573), .ZN(n380) );
  XNOR2_X1 U485 ( .A(n396), .B(n573), .ZN(n805) );
  XNOR2_X1 U486 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U487 ( .A1(n560), .A2(n381), .ZN(n391) );
  AND2_X1 U488 ( .A1(n375), .A2(n562), .ZN(n381) );
  NAND2_X1 U489 ( .A1(n600), .A2(n599), .ZN(n605) );
  XNOR2_X1 U490 ( .A(G143), .B(G128), .ZN(n382) );
  XNOR2_X1 U491 ( .A(n405), .B(n366), .ZN(n404) );
  NAND2_X1 U492 ( .A1(n407), .A2(n406), .ZN(n405) );
  NAND2_X1 U493 ( .A1(n603), .A2(n385), .ZN(n383) );
  NAND2_X1 U494 ( .A1(n383), .A2(n384), .ZN(n604) );
  AND2_X1 U495 ( .A1(n602), .A2(KEYINPUT44), .ZN(n385) );
  NOR2_X1 U496 ( .A1(n375), .A2(n583), .ZN(n567) );
  NOR2_X1 U497 ( .A1(n453), .A2(n362), .ZN(n386) );
  NAND2_X1 U498 ( .A1(n386), .A2(n447), .ZN(n638) );
  XNOR2_X1 U499 ( .A(n370), .B(n500), .ZN(n611) );
  BUF_X1 U500 ( .A(n370), .Z(n728) );
  BUF_X1 U501 ( .A(n399), .Z(n387) );
  XNOR2_X1 U502 ( .A(n419), .B(G101), .ZN(n388) );
  INV_X1 U503 ( .A(n577), .ZN(n398) );
  XNOR2_X1 U504 ( .A(n388), .B(G137), .ZN(n491) );
  XNOR2_X2 U505 ( .A(n390), .B(KEYINPUT85), .ZN(n601) );
  XNOR2_X2 U506 ( .A(n489), .B(n363), .ZN(n793) );
  XNOR2_X2 U507 ( .A(n477), .B(G134), .ZN(n489) );
  XNOR2_X2 U508 ( .A(G143), .B(G128), .ZN(n477) );
  NAND2_X1 U509 ( .A1(n395), .A2(n367), .ZN(n576) );
  INV_X1 U510 ( .A(n805), .ZN(n395) );
  NAND2_X1 U511 ( .A1(n377), .A2(n397), .ZN(n396) );
  XNOR2_X1 U512 ( .A(n637), .B(n408), .ZN(n407) );
  XNOR2_X2 U513 ( .A(G146), .B(n793), .ZN(n505) );
  XNOR2_X1 U514 ( .A(n387), .B(G119), .ZN(G21) );
  XNOR2_X2 U515 ( .A(n421), .B(n494), .ZN(n787) );
  XNOR2_X2 U516 ( .A(n401), .B(n400), .ZN(n494) );
  XNOR2_X2 U517 ( .A(KEYINPUT3), .B(G119), .ZN(n400) );
  XNOR2_X2 U518 ( .A(n403), .B(n784), .ZN(n501) );
  XNOR2_X2 U519 ( .A(n402), .B(G107), .ZN(n784) );
  NAND2_X1 U520 ( .A1(n404), .A2(n729), .ZN(n639) );
  INV_X1 U521 ( .A(n638), .ZN(n406) );
  XNOR2_X2 U522 ( .A(n412), .B(n411), .ZN(n561) );
  XNOR2_X2 U523 ( .A(n415), .B(n413), .ZN(n581) );
  XOR2_X1 U524 ( .A(n559), .B(KEYINPUT43), .Z(n418) );
  INV_X1 U525 ( .A(KEYINPUT5), .ZN(n490) );
  INV_X1 U526 ( .A(KEYINPUT108), .ZN(n529) );
  XNOR2_X1 U527 ( .A(n491), .B(n490), .ZN(n496) );
  XNOR2_X1 U528 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U529 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U530 ( .A(n465), .B(n464), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n517), .B(n518), .ZN(n521) );
  BUF_X1 U532 ( .A(n532), .Z(n615) );
  BUF_X1 U533 ( .A(n699), .Z(n770) );
  XNOR2_X1 U534 ( .A(KEYINPUT16), .B(G122), .ZN(n420) );
  XNOR2_X1 U535 ( .A(n420), .B(KEYINPUT72), .ZN(n421) );
  XNOR2_X1 U536 ( .A(n423), .B(n422), .ZN(n426) );
  NAND2_X1 U537 ( .A1(n796), .A2(G224), .ZN(n424) );
  XNOR2_X1 U538 ( .A(n424), .B(KEYINPUT88), .ZN(n425) );
  XNOR2_X1 U539 ( .A(n426), .B(n425), .ZN(n428) );
  XNOR2_X1 U540 ( .A(n382), .B(n466), .ZN(n427) );
  XNOR2_X1 U541 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X2 U542 ( .A(n430), .B(n429), .ZN(n675) );
  NAND2_X1 U543 ( .A1(n507), .A2(n431), .ZN(n433) );
  NAND2_X1 U544 ( .A1(n433), .A2(G214), .ZN(n432) );
  XNOR2_X1 U545 ( .A(n432), .B(KEYINPUT90), .ZN(n550) );
  NAND2_X1 U546 ( .A1(n550), .A2(n544), .ZN(n436) );
  NAND2_X1 U547 ( .A1(n433), .A2(G210), .ZN(n439) );
  XNOR2_X1 U548 ( .A(KEYINPUT79), .B(KEYINPUT87), .ZN(n434) );
  XNOR2_X1 U549 ( .A(n439), .B(n434), .ZN(n435) );
  NOR2_X1 U550 ( .A1(n436), .A2(n435), .ZN(n437) );
  NAND2_X1 U551 ( .A1(n675), .A2(n437), .ZN(n447) );
  INV_X1 U552 ( .A(KEYINPUT79), .ZN(n438) );
  XNOR2_X1 U553 ( .A(n439), .B(n438), .ZN(n545) );
  INV_X1 U554 ( .A(KEYINPUT87), .ZN(n443) );
  NAND2_X1 U555 ( .A1(n545), .A2(n443), .ZN(n450) );
  INV_X1 U556 ( .A(n450), .ZN(n440) );
  INV_X1 U557 ( .A(n544), .ZN(n669) );
  NAND2_X1 U558 ( .A1(n440), .A2(n669), .ZN(n442) );
  OR2_X1 U559 ( .A1(n550), .A2(KEYINPUT87), .ZN(n441) );
  NAND2_X1 U560 ( .A1(n442), .A2(n441), .ZN(n446) );
  NAND2_X1 U561 ( .A1(n550), .A2(n669), .ZN(n444) );
  OR2_X1 U562 ( .A1(n545), .A2(n443), .ZN(n448) );
  NOR2_X1 U563 ( .A1(n444), .A2(n448), .ZN(n445) );
  INV_X1 U564 ( .A(n448), .ZN(n449) );
  NAND2_X1 U565 ( .A1(n449), .A2(n550), .ZN(n451) );
  AND2_X1 U566 ( .A1(n451), .A2(n450), .ZN(n452) );
  NOR2_X1 U567 ( .A1(n675), .A2(n452), .ZN(n453) );
  XNOR2_X2 U568 ( .A(n638), .B(KEYINPUT19), .ZN(n626) );
  NOR2_X1 U569 ( .A1(G898), .A2(n796), .ZN(n789) );
  NAND2_X1 U570 ( .A1(n789), .A2(G902), .ZN(n454) );
  NAND2_X1 U571 ( .A1(n796), .A2(G952), .ZN(n539) );
  NAND2_X1 U572 ( .A1(n454), .A2(n539), .ZN(n457) );
  INV_X1 U573 ( .A(KEYINPUT14), .ZN(n455) );
  XNOR2_X1 U574 ( .A(n456), .B(n455), .ZN(n754) );
  INV_X1 U575 ( .A(n754), .ZN(n535) );
  AND2_X1 U576 ( .A1(n457), .A2(n535), .ZN(n458) );
  NAND2_X1 U577 ( .A1(n626), .A2(n458), .ZN(n459) );
  XNOR2_X1 U578 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n472) );
  NAND2_X1 U579 ( .A1(n492), .A2(G214), .ZN(n460) );
  XNOR2_X1 U580 ( .A(n461), .B(n460), .ZN(n465) );
  XNOR2_X1 U581 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U582 ( .A(n520), .B(n469), .ZN(n470) );
  XOR2_X1 U583 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n474) );
  XNOR2_X1 U584 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U585 ( .A1(G217), .A2(n509), .ZN(n479) );
  INV_X1 U586 ( .A(n489), .ZN(n478) );
  XNOR2_X1 U587 ( .A(KEYINPUT100), .B(G478), .ZN(n481) );
  NAND2_X1 U588 ( .A1(n581), .A2(n571), .ZN(n607) );
  NAND2_X1 U589 ( .A1(n544), .A2(G234), .ZN(n484) );
  XNOR2_X1 U590 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n483) );
  XNOR2_X1 U591 ( .A(n484), .B(n483), .ZN(n522) );
  NAND2_X1 U592 ( .A1(n522), .A2(G221), .ZN(n486) );
  INV_X1 U593 ( .A(KEYINPUT21), .ZN(n485) );
  XNOR2_X1 U594 ( .A(n486), .B(n485), .ZN(n725) );
  INV_X1 U595 ( .A(n725), .ZN(n552) );
  AND2_X1 U596 ( .A1(n492), .A2(G210), .ZN(n493) );
  XNOR2_X1 U597 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X2 U598 ( .A(n497), .B(n505), .ZN(n683) );
  NAND2_X1 U599 ( .A1(n683), .A2(n507), .ZN(n499) );
  INV_X1 U600 ( .A(G472), .ZN(n498) );
  INV_X1 U601 ( .A(KEYINPUT104), .ZN(n500) );
  NAND2_X1 U602 ( .A1(G227), .A2(n796), .ZN(n502) );
  XNOR2_X1 U603 ( .A(n506), .B(n505), .ZN(n701) );
  NAND2_X1 U604 ( .A1(n701), .A2(n507), .ZN(n508) );
  XNOR2_X1 U605 ( .A(n532), .B(KEYINPUT1), .ZN(n564) );
  INV_X1 U606 ( .A(n564), .ZN(n592) );
  INV_X1 U607 ( .A(n592), .ZN(n729) );
  NAND2_X1 U608 ( .A1(G221), .A2(n509), .ZN(n518) );
  XOR2_X1 U609 ( .A(KEYINPUT24), .B(G128), .Z(n511) );
  XNOR2_X1 U610 ( .A(G110), .B(G119), .ZN(n510) );
  XNOR2_X1 U611 ( .A(n511), .B(n510), .ZN(n516) );
  INV_X1 U612 ( .A(n512), .ZN(n514) );
  XNOR2_X1 U613 ( .A(KEYINPUT23), .B(KEYINPUT92), .ZN(n513) );
  XNOR2_X1 U614 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U615 ( .A(n520), .B(n519), .ZN(n794) );
  NAND2_X1 U616 ( .A1(n522), .A2(G217), .ZN(n524) );
  INV_X1 U617 ( .A(KEYINPUT75), .ZN(n523) );
  XNOR2_X1 U618 ( .A(n524), .B(n523), .ZN(n525) );
  INV_X1 U619 ( .A(n561), .ZN(n526) );
  OR2_X1 U620 ( .A1(n729), .A2(n526), .ZN(n527) );
  NOR2_X1 U621 ( .A1(n527), .A2(n611), .ZN(n528) );
  AND2_X1 U622 ( .A1(n376), .A2(n528), .ZN(n577) );
  XOR2_X1 U623 ( .A(G110), .B(n577), .Z(G12) );
  NAND2_X1 U624 ( .A1(n611), .A2(n550), .ZN(n531) );
  XNOR2_X1 U625 ( .A(n531), .B(n530), .ZN(n534) );
  NOR2_X1 U626 ( .A1(n561), .A2(n552), .ZN(n730) );
  NAND2_X1 U627 ( .A1(n730), .A2(n615), .ZN(n533) );
  NAND2_X1 U628 ( .A1(n534), .A2(n587), .ZN(n620) );
  INV_X1 U629 ( .A(n620), .ZN(n543) );
  NAND2_X1 U630 ( .A1(G902), .A2(n535), .ZN(n536) );
  NOR2_X1 U631 ( .A1(G900), .A2(n536), .ZN(n537) );
  NAND2_X1 U632 ( .A1(G953), .A2(n537), .ZN(n538) );
  XNOR2_X1 U633 ( .A(n538), .B(KEYINPUT105), .ZN(n541) );
  NOR2_X1 U634 ( .A1(n754), .A2(n539), .ZN(n540) );
  NOR2_X1 U635 ( .A1(n541), .A2(n540), .ZN(n618) );
  NOR2_X1 U636 ( .A1(n618), .A2(n581), .ZN(n542) );
  NAND2_X1 U637 ( .A1(n543), .A2(n542), .ZN(n549) );
  NAND2_X1 U638 ( .A1(n675), .A2(n544), .ZN(n546) );
  INV_X1 U639 ( .A(n608), .ZN(n547) );
  INV_X1 U640 ( .A(n571), .ZN(n582) );
  NAND2_X1 U641 ( .A1(n547), .A2(n582), .ZN(n548) );
  NOR2_X1 U642 ( .A1(n549), .A2(n548), .ZN(n640) );
  XOR2_X1 U643 ( .A(G143), .B(n640), .Z(G45) );
  INV_X1 U644 ( .A(n550), .ZN(n739) );
  INV_X1 U645 ( .A(KEYINPUT6), .ZN(n551) );
  NOR2_X1 U646 ( .A1(n552), .A2(n618), .ZN(n553) );
  NAND2_X1 U647 ( .A1(n561), .A2(n553), .ZN(n610) );
  XNOR2_X1 U648 ( .A(n554), .B(KEYINPUT106), .ZN(n556) );
  INV_X1 U649 ( .A(n581), .ZN(n572) );
  NAND2_X1 U650 ( .A1(n572), .A2(n571), .ZN(n555) );
  XNOR2_X2 U651 ( .A(KEYINPUT101), .B(n555), .ZN(n717) );
  NAND2_X1 U652 ( .A1(n556), .A2(n717), .ZN(n637) );
  NOR2_X1 U653 ( .A1(n739), .A2(n637), .ZN(n557) );
  XNOR2_X1 U654 ( .A(n557), .B(KEYINPUT107), .ZN(n558) );
  NOR2_X1 U655 ( .A1(n729), .A2(n558), .ZN(n559) );
  NAND2_X1 U656 ( .A1(n418), .A2(n608), .ZN(n656) );
  XNOR2_X1 U657 ( .A(n656), .B(G140), .ZN(G42) );
  XNOR2_X1 U658 ( .A(n561), .B(KEYINPUT103), .ZN(n724) );
  INV_X1 U659 ( .A(n724), .ZN(n594) );
  AND2_X1 U660 ( .A1(n729), .A2(n594), .ZN(n562) );
  INV_X1 U661 ( .A(KEYINPUT78), .ZN(n563) );
  XOR2_X1 U662 ( .A(KEYINPUT35), .B(KEYINPUT77), .Z(n573) );
  NAND2_X1 U663 ( .A1(n564), .A2(n730), .ZN(n583) );
  XNOR2_X1 U664 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n566) );
  XNOR2_X1 U665 ( .A(n567), .B(n566), .ZN(n747) );
  NOR2_X1 U666 ( .A1(n747), .A2(n569), .ZN(n570) );
  INV_X1 U667 ( .A(KEYINPUT44), .ZN(n574) );
  INV_X1 U668 ( .A(KEYINPUT68), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n380), .A2(n602), .ZN(n575) );
  NAND2_X1 U670 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U671 ( .A(n601), .B(KEYINPUT84), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n578), .A2(n603), .ZN(n600) );
  INV_X1 U673 ( .A(n601), .ZN(n579) );
  NAND2_X1 U674 ( .A1(n579), .A2(KEYINPUT44), .ZN(n580) );
  NAND2_X1 U675 ( .A1(n580), .A2(KEYINPUT65), .ZN(n598) );
  AND2_X1 U676 ( .A1(n582), .A2(n581), .ZN(n720) );
  NOR2_X1 U677 ( .A1(n717), .A2(n720), .ZN(n641) );
  NOR2_X1 U678 ( .A1(n583), .A2(n728), .ZN(n735) );
  INV_X1 U679 ( .A(n569), .ZN(n585) );
  NAND2_X1 U680 ( .A1(n735), .A2(n585), .ZN(n586) );
  XNOR2_X1 U681 ( .A(n586), .B(KEYINPUT31), .ZN(n721) );
  NAND2_X1 U682 ( .A1(n587), .A2(n728), .ZN(n588) );
  NOR2_X1 U683 ( .A1(n588), .A2(n569), .ZN(n707) );
  NOR2_X1 U684 ( .A1(n721), .A2(n707), .ZN(n589) );
  NOR2_X1 U685 ( .A1(n641), .A2(n589), .ZN(n590) );
  XNOR2_X1 U686 ( .A(n590), .B(KEYINPUT102), .ZN(n596) );
  XOR2_X1 U687 ( .A(KEYINPUT83), .B(n593), .Z(n595) );
  NOR2_X1 U688 ( .A1(n595), .A2(n594), .ZN(n705) );
  NOR2_X1 U689 ( .A1(n596), .A2(n705), .ZN(n597) );
  INV_X1 U690 ( .A(n607), .ZN(n741) );
  NOR2_X1 U691 ( .A1(n740), .A2(n739), .ZN(n744) );
  NAND2_X1 U692 ( .A1(n741), .A2(n744), .ZN(n609) );
  XOR2_X1 U693 ( .A(n609), .B(KEYINPUT41), .Z(n758) );
  XOR2_X1 U694 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n613) );
  NAND2_X1 U695 ( .A1(n369), .A2(n611), .ZN(n612) );
  NAND2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n628) );
  OR2_X1 U697 ( .A1(n740), .A2(n618), .ZN(n619) );
  NOR2_X2 U698 ( .A1(n620), .A2(n619), .ZN(n622) );
  INV_X1 U699 ( .A(KEYINPUT39), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n622), .B(n621), .ZN(n655) );
  NAND2_X1 U701 ( .A1(n655), .A2(n717), .ZN(n624) );
  XOR2_X1 U702 ( .A(KEYINPUT40), .B(KEYINPUT111), .Z(n623) );
  NAND2_X1 U703 ( .A1(n808), .A2(n806), .ZN(n625) );
  XNOR2_X1 U704 ( .A(n625), .B(KEYINPUT46), .ZN(n653) );
  INV_X1 U705 ( .A(n626), .ZN(n627) );
  NOR2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n714) );
  INV_X1 U707 ( .A(n641), .ZN(n743) );
  NOR2_X1 U708 ( .A1(KEYINPUT81), .A2(n743), .ZN(n629) );
  NOR2_X1 U709 ( .A1(KEYINPUT73), .A2(n629), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n714), .A2(n630), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n631), .A2(KEYINPUT47), .ZN(n636) );
  XOR2_X1 U712 ( .A(KEYINPUT73), .B(n743), .Z(n633) );
  INV_X1 U713 ( .A(KEYINPUT47), .ZN(n632) );
  AND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n714), .A2(n634), .ZN(n635) );
  AND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n639), .B(KEYINPUT113), .ZN(n803) );
  INV_X1 U718 ( .A(n803), .ZN(n649) );
  INV_X1 U719 ( .A(n640), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n641), .A2(KEYINPUT47), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n645), .A2(n642), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n643), .A2(KEYINPUT81), .ZN(n647) );
  INV_X1 U723 ( .A(KEYINPUT81), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X2 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(KEYINPUT48), .ZN(n661) );
  NAND2_X1 U729 ( .A1(n655), .A2(n720), .ZN(n723) );
  AND2_X1 U730 ( .A1(n723), .A2(n656), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n661), .A2(n658), .ZN(n792) );
  INV_X1 U732 ( .A(KEYINPUT2), .ZN(n756) );
  INV_X1 U733 ( .A(n657), .ZN(n776) );
  NAND2_X1 U734 ( .A1(n756), .A2(KEYINPUT74), .ZN(n660) );
  INV_X1 U735 ( .A(n658), .ZN(n659) );
  NOR2_X1 U736 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U737 ( .A1(n662), .A2(n661), .ZN(n665) );
  INV_X1 U738 ( .A(KEYINPUT74), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n792), .A2(n663), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U741 ( .A1(n776), .A2(n666), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n670), .A2(n669), .ZN(n672) );
  INV_X1 U744 ( .A(KEYINPUT64), .ZN(n671) );
  XNOR2_X2 U745 ( .A(n672), .B(n671), .ZN(n699) );
  NAND2_X1 U746 ( .A1(n699), .A2(G210), .ZN(n677) );
  XNOR2_X1 U747 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n673) );
  XNOR2_X1 U748 ( .A(n673), .B(KEYINPUT55), .ZN(n674) );
  XNOR2_X1 U749 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U750 ( .A(n677), .B(n676), .ZN(n679) );
  INV_X1 U751 ( .A(G952), .ZN(n678) );
  NOR2_X2 U752 ( .A1(n679), .A2(n775), .ZN(n681) );
  XNOR2_X1 U753 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n680) );
  XNOR2_X1 U754 ( .A(n681), .B(n680), .ZN(G51) );
  NAND2_X1 U755 ( .A1(n699), .A2(G472), .ZN(n685) );
  XOR2_X1 U756 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n682) );
  XNOR2_X1 U757 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X2 U758 ( .A1(n686), .A2(n775), .ZN(n688) );
  XNOR2_X1 U759 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n687) );
  XNOR2_X1 U760 ( .A(n688), .B(n687), .ZN(G57) );
  NAND2_X1 U761 ( .A1(n699), .A2(G475), .ZN(n691) );
  XNOR2_X1 U762 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X2 U763 ( .A1(n692), .A2(n775), .ZN(n694) );
  XNOR2_X1 U764 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n693) );
  XNOR2_X1 U765 ( .A(n694), .B(n693), .ZN(G60) );
  NAND2_X1 U766 ( .A1(n699), .A2(G217), .ZN(n696) );
  XNOR2_X1 U767 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X2 U768 ( .A1(n697), .A2(n775), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n698), .B(KEYINPUT122), .ZN(G66) );
  NAND2_X1 U770 ( .A1(n770), .A2(G469), .ZN(n703) );
  XNOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n700) );
  XNOR2_X1 U772 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U773 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U774 ( .A1(n704), .A2(n775), .ZN(G54) );
  XOR2_X1 U775 ( .A(G101), .B(n374), .Z(G3) );
  NAND2_X1 U776 ( .A1(n707), .A2(n717), .ZN(n706) );
  XNOR2_X1 U777 ( .A(n706), .B(G104), .ZN(G6) );
  XNOR2_X1 U778 ( .A(G107), .B(KEYINPUT27), .ZN(n711) );
  XOR2_X1 U779 ( .A(KEYINPUT26), .B(KEYINPUT116), .Z(n709) );
  NAND2_X1 U780 ( .A1(n707), .A2(n720), .ZN(n708) );
  XNOR2_X1 U781 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U782 ( .A(n711), .B(n710), .ZN(G9) );
  XOR2_X1 U783 ( .A(G128), .B(KEYINPUT29), .Z(n713) );
  NAND2_X1 U784 ( .A1(n714), .A2(n720), .ZN(n712) );
  XNOR2_X1 U785 ( .A(n713), .B(n712), .ZN(G30) );
  XOR2_X1 U786 ( .A(G146), .B(KEYINPUT117), .Z(n716) );
  NAND2_X1 U787 ( .A1(n714), .A2(n717), .ZN(n715) );
  XNOR2_X1 U788 ( .A(n716), .B(n715), .ZN(G48) );
  NAND2_X1 U789 ( .A1(n721), .A2(n717), .ZN(n718) );
  XNOR2_X1 U790 ( .A(n718), .B(KEYINPUT118), .ZN(n719) );
  XNOR2_X1 U791 ( .A(G113), .B(n719), .ZN(G15) );
  NAND2_X1 U792 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U793 ( .A(n722), .B(G116), .ZN(G18) );
  XNOR2_X1 U794 ( .A(G134), .B(n723), .ZN(G36) );
  INV_X1 U795 ( .A(n758), .ZN(n738) );
  NOR2_X1 U796 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U797 ( .A(n726), .B(KEYINPUT49), .ZN(n727) );
  NAND2_X1 U798 ( .A1(n728), .A2(n727), .ZN(n733) );
  NOR2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U800 ( .A(n731), .B(KEYINPUT50), .ZN(n732) );
  NOR2_X1 U801 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U802 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U803 ( .A(KEYINPUT51), .B(n736), .ZN(n737) );
  NAND2_X1 U804 ( .A1(n738), .A2(n737), .ZN(n751) );
  NAND2_X1 U805 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U806 ( .A1(n742), .A2(n741), .ZN(n746) );
  NAND2_X1 U807 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U808 ( .A1(n746), .A2(n745), .ZN(n749) );
  INV_X1 U809 ( .A(n747), .ZN(n748) );
  NAND2_X1 U810 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U811 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U812 ( .A(KEYINPUT52), .B(n752), .Z(n753) );
  NOR2_X1 U813 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U814 ( .A1(n755), .A2(G952), .ZN(n767) );
  XOR2_X1 U815 ( .A(n360), .B(KEYINPUT80), .Z(n757) );
  NAND2_X1 U816 ( .A1(n757), .A2(n756), .ZN(n761) );
  NOR2_X1 U817 ( .A1(n747), .A2(n758), .ZN(n759) );
  NOR2_X1 U818 ( .A1(G953), .A2(n759), .ZN(n760) );
  NAND2_X1 U819 ( .A1(n761), .A2(n760), .ZN(n765) );
  INV_X1 U820 ( .A(n360), .ZN(n763) );
  NAND2_X1 U821 ( .A1(KEYINPUT2), .A2(KEYINPUT80), .ZN(n762) );
  NOR2_X1 U822 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U823 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U824 ( .A(n768), .B(KEYINPUT53), .ZN(n769) );
  XNOR2_X1 U825 ( .A(KEYINPUT119), .B(n769), .ZN(G75) );
  NAND2_X1 U826 ( .A1(n770), .A2(G478), .ZN(n773) );
  XOR2_X1 U827 ( .A(n771), .B(KEYINPUT121), .Z(n772) );
  XNOR2_X1 U828 ( .A(n773), .B(n772), .ZN(n774) );
  NOR2_X1 U829 ( .A1(n775), .A2(n774), .ZN(G63) );
  NAND2_X1 U830 ( .A1(n776), .A2(n796), .ZN(n777) );
  XOR2_X1 U831 ( .A(KEYINPUT123), .B(n777), .Z(n781) );
  NAND2_X1 U832 ( .A1(G953), .A2(G224), .ZN(n778) );
  XNOR2_X1 U833 ( .A(KEYINPUT61), .B(n778), .ZN(n779) );
  NAND2_X1 U834 ( .A1(n779), .A2(G898), .ZN(n780) );
  NAND2_X1 U835 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U836 ( .A(n782), .B(KEYINPUT126), .ZN(n783) );
  XNOR2_X1 U837 ( .A(KEYINPUT124), .B(n783), .ZN(n791) );
  XNOR2_X1 U838 ( .A(n784), .B(G101), .ZN(n785) );
  XOR2_X1 U839 ( .A(KEYINPUT125), .B(n785), .Z(n786) );
  XNOR2_X1 U840 ( .A(n787), .B(n786), .ZN(n788) );
  NOR2_X1 U841 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U842 ( .A(n791), .B(n790), .ZN(G69) );
  BUF_X1 U843 ( .A(n792), .Z(n795) );
  XOR2_X1 U844 ( .A(n794), .B(n793), .Z(n798) );
  XNOR2_X1 U845 ( .A(n795), .B(n798), .ZN(n797) );
  NAND2_X1 U846 ( .A1(n797), .A2(n796), .ZN(n802) );
  XNOR2_X1 U847 ( .A(G227), .B(n798), .ZN(n799) );
  NAND2_X1 U848 ( .A1(n799), .A2(G900), .ZN(n800) );
  NAND2_X1 U849 ( .A1(n800), .A2(G953), .ZN(n801) );
  NAND2_X1 U850 ( .A1(n802), .A2(n801), .ZN(G72) );
  XNOR2_X1 U851 ( .A(G125), .B(n803), .ZN(n804) );
  XNOR2_X1 U852 ( .A(n804), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U853 ( .A(G122), .B(n380), .Z(G24) );
  XOR2_X1 U854 ( .A(G131), .B(n806), .Z(n807) );
  XNOR2_X1 U855 ( .A(KEYINPUT127), .B(n807), .ZN(G33) );
  XNOR2_X1 U856 ( .A(G137), .B(n378), .ZN(G39) );
endmodule

