//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT95), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  AND2_X1   g003(.A1(new_n204), .A2(KEYINPUT92), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G8gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT89), .ZN(new_n215));
  OR3_X1    g014(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n217), .A2(KEYINPUT90), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(KEYINPUT90), .B2(new_n217), .ZN(new_n219));
  XNOR2_X1  g018(.A(G43gat), .B(G50gat), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n215), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n216), .B(KEYINPUT91), .ZN(new_n225));
  OAI221_X1 g024(.A(new_n223), .B1(KEYINPUT15), .B2(new_n220), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n213), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n222), .A2(new_n226), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(KEYINPUT17), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n212), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n228), .B(new_n229), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n236), .A2(KEYINPUT93), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n230), .A2(new_n212), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n228), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n229), .B(KEYINPUT13), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n234), .B2(new_n235), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT94), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT94), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n244), .B(new_n241), .C1(new_n234), .C2(new_n235), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n236), .A2(KEYINPUT93), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n237), .A2(new_n243), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G197gat), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT11), .B(G169gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n251), .B(KEYINPUT12), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n236), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n254), .A2(new_n242), .A3(new_n252), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n203), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  AOI211_X1 g056(.A(KEYINPUT95), .B(new_n255), .C1(new_n247), .C2(new_n252), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G120gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G113gat), .ZN(new_n261));
  INV_X1    g060(.A(G113gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G120gat), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT1), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G127gat), .B(G134gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G127gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G134gat), .ZN(new_n268));
  INV_X1    g067(.A(G134gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G127gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n270), .A3(KEYINPUT69), .ZN(new_n271));
  OR3_X1    g070(.A1(new_n269), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n273), .A2(new_n274), .A3(new_n264), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n269), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(new_n265), .B2(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n263), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT70), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n266), .B1(new_n275), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT71), .ZN(new_n283));
  INV_X1    g082(.A(new_n266), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n274), .B1(new_n273), .B2(new_n264), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n280), .A2(KEYINPUT70), .A3(new_n271), .A4(new_n272), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT26), .ZN(new_n292));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(new_n291), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT68), .B(G183gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT27), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G190gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT28), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT27), .B(G183gat), .Z(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n307), .A2(new_n308), .A3(G190gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n299), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT67), .B1(new_n291), .B2(KEYINPUT23), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n312), .B(new_n313), .C1(G169gat), .C2(G176gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n311), .A2(new_n295), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n293), .A2(KEYINPUT24), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT24), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(G183gat), .A3(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(G183gat), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n316), .A2(new_n318), .B1(new_n319), .B2(new_n305), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n313), .A2(G176gat), .ZN(new_n322));
  OR2_X1    g121(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT66), .ZN(new_n326));
  AND2_X1   g125(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT66), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(new_n322), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT25), .B1(new_n321), .B2(new_n332), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n302), .A2(new_n305), .B1(new_n316), .B2(new_n318), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n313), .A2(G176gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT25), .B1(new_n335), .B2(G169gat), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n334), .A2(new_n315), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n310), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n290), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT25), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n330), .B1(new_n329), .B2(new_n322), .ZN(new_n341));
  AND4_X1   g140(.A1(new_n330), .A2(new_n322), .A3(new_n323), .A4(new_n324), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n316), .A2(new_n318), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n319), .A2(new_n305), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n314), .A2(new_n295), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n311), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n340), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n337), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G183gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n300), .B1(new_n354), .B2(KEYINPUT27), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n308), .B1(new_n355), .B2(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n309), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n349), .A2(new_n350), .B1(new_n358), .B2(new_n299), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(new_n283), .A3(new_n289), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n339), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G227gat), .ZN(new_n362));
  INV_X1    g161(.A(G233gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT64), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT32), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT33), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G15gat), .B(G43gat), .Z(new_n370));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n367), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n366), .B(KEYINPUT32), .C1(new_n368), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OR3_X1    g175(.A1(new_n361), .A2(KEYINPUT34), .A3(new_n365), .ZN(new_n377));
  INV_X1    g176(.A(new_n364), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n339), .A2(new_n378), .A3(new_n360), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT72), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT34), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n379), .B2(KEYINPUT34), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n377), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n381), .A2(new_n382), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n385), .A2(new_n377), .A3(new_n375), .A4(new_n373), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G141gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G148gat), .ZN(new_n389));
  INV_X1    g188(.A(G148gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G141gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G155gat), .B(G162gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT2), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n395), .B2(new_n392), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G197gat), .B(G204gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT22), .ZN(new_n400));
  INV_X1    g199(.A(G211gat), .ZN(new_n401));
  INV_X1    g200(.A(G218gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G211gat), .B(G218gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n399), .A3(new_n403), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n398), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n407), .A2(KEYINPUT73), .A3(new_n408), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT73), .B1(new_n407), .B2(new_n408), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n398), .B2(new_n412), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n409), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n414), .B1(new_n421), .B2(new_n413), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n424), .A2(KEYINPUT83), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(KEYINPUT83), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(G22gat), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G78gat), .B(G106gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT82), .ZN(new_n429));
  XOR2_X1   g228(.A(KEYINPUT31), .B(G50gat), .Z(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n423), .A2(G22gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n433), .B2(KEYINPUT84), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n427), .B(new_n434), .C1(KEYINPUT84), .C2(new_n433), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n423), .A2(G22gat), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n431), .B1(new_n436), .B2(new_n432), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n387), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT35), .ZN(new_n441));
  XNOR2_X1  g240(.A(G8gat), .B(G36gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(G64gat), .B(G92gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  NAND2_X1  g243(.A1(G226gat), .A2(G233gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n410), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n321), .A2(new_n332), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n337), .B1(new_n447), .B2(new_n340), .ZN(new_n448));
  INV_X1    g247(.A(new_n299), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n356), .B2(new_n357), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n446), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n310), .B(new_n445), .C1(new_n333), .C2(new_n337), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n451), .A2(new_n452), .A3(new_n409), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n418), .B1(new_n451), .B2(new_n452), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT74), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI211_X1 g255(.A(KEYINPUT74), .B(new_n418), .C1(new_n451), .C2(new_n452), .ZN(new_n457));
  OAI211_X1 g256(.A(KEYINPUT30), .B(new_n444), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n446), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n452), .B1(new_n359), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n418), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n455), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n451), .A2(new_n452), .A3(new_n409), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n457), .ZN(new_n465));
  INV_X1    g264(.A(new_n444), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n458), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT75), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n457), .B1(new_n463), .B2(new_n462), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(new_n466), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT30), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT75), .B(new_n444), .C1(new_n456), .C2(new_n457), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT76), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n471), .A2(KEYINPUT76), .A3(new_n473), .A4(new_n472), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n287), .B(new_n398), .ZN(new_n480));
  NAND2_X1  g279(.A1(G225gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n479), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT3), .B1(new_n396), .B2(new_n397), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n392), .A2(new_n395), .ZN(new_n485));
  INV_X1    g284(.A(new_n393), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n412), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n481), .B1(new_n490), .B2(new_n287), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT4), .B1(new_n287), .B2(new_n398), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n283), .A2(KEYINPUT4), .A3(new_n398), .A4(new_n289), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n493), .B2(new_n494), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n483), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(G1gat), .B(G29gat), .Z(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G57gat), .B(G85gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n287), .A2(KEYINPUT4), .A3(new_n398), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n283), .A2(new_n398), .A3(new_n289), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT4), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n490), .A2(new_n287), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n508), .A2(new_n481), .A3(new_n510), .A4(new_n479), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n498), .A2(new_n503), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n503), .B1(new_n498), .B2(new_n511), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT87), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n515), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT87), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n517), .A2(new_n518), .A3(new_n513), .A4(new_n512), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n440), .A2(new_n441), .A3(new_n478), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n514), .A2(KEYINPUT80), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT80), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n512), .A2(new_n524), .A3(new_n513), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n520), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n527), .A2(new_n478), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n528), .B1(new_n527), .B2(new_n478), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n529), .A2(new_n530), .A3(new_n439), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n522), .B1(new_n531), .B2(new_n441), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n384), .A2(new_n386), .A3(KEYINPUT36), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT36), .B1(new_n384), .B2(new_n386), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n438), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n476), .A2(new_n477), .ZN(new_n538));
  INV_X1    g337(.A(new_n468), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT39), .ZN(new_n541));
  AOI211_X1 g340(.A(new_n509), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n542), .A2(KEYINPUT85), .A3(new_n481), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT85), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n506), .A2(new_n507), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n545), .A2(new_n510), .A3(new_n504), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n546), .B2(new_n482), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n541), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT85), .B1(new_n542), .B2(new_n481), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n544), .A3(new_n482), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n480), .A2(new_n482), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n549), .A2(KEYINPUT39), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n548), .A2(new_n552), .A3(new_n503), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n517), .ZN(new_n556));
  INV_X1    g355(.A(new_n503), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n549), .A2(new_n550), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(new_n541), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n554), .B1(new_n559), .B2(new_n552), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n537), .B1(new_n540), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n466), .A2(KEYINPUT37), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n467), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n470), .A2(KEYINPUT37), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT38), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n471), .A2(new_n473), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT37), .B1(new_n460), .B2(new_n418), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n460), .B2(new_n409), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT38), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n564), .A2(KEYINPUT88), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT88), .B1(new_n564), .B2(new_n571), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n567), .B(new_n568), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n574), .A2(new_n521), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n536), .B1(new_n562), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n537), .B1(new_n529), .B2(new_n530), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n202), .B(new_n259), .C1(new_n533), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n527), .A2(new_n478), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT81), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n527), .A2(new_n478), .A3(new_n528), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n440), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT35), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n585), .A2(new_n522), .B1(new_n577), .B2(new_n576), .ZN(new_n586));
  INV_X1    g385(.A(new_n259), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT96), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G99gat), .B(G106gat), .Z(new_n590));
  INV_X1    g389(.A(G85gat), .ZN(new_n591));
  INV_X1    g390(.A(G92gat), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT97), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n590), .A2(KEYINPUT98), .B1(new_n593), .B2(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n591), .B2(new_n592), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n594), .B(new_n596), .C1(KEYINPUT7), .C2(new_n593), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n590), .A2(KEYINPUT98), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(new_n227), .B2(new_n232), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n231), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n597), .B(new_n598), .Z(new_n604));
  AND2_X1   g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n227), .A2(new_n604), .B1(KEYINPUT41), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n607), .B(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G190gat), .B(G218gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT100), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n607), .B(new_n608), .ZN(new_n616));
  INV_X1    g415(.A(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G57gat), .B(G64gat), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G71gat), .B(G78gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT21), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n267), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n212), .B1(new_n626), .B2(new_n625), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G155gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G183gat), .B(G211gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n632), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n604), .A2(new_n624), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n599), .B2(new_n625), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n604), .A2(new_n640), .A3(new_n624), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT10), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n624), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n638), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n642), .A2(G230gat), .A3(G233gat), .A4(new_n643), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n619), .A2(new_n637), .A3(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n658), .A2(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(KEYINPUT102), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n526), .A2(KEYINPUT103), .A3(new_n520), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT103), .B1(new_n526), .B2(new_n520), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n589), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT104), .B(G1gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1324gat));
  INV_X1    g466(.A(new_n589), .ZN(new_n668));
  INV_X1    g467(.A(new_n661), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  NOR4_X1   g469(.A1(new_n668), .A2(new_n478), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n669), .A2(new_n478), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n211), .B1(new_n672), .B2(new_n589), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(KEYINPUT42), .B2(new_n671), .ZN(G1325gat));
  INV_X1    g474(.A(G15gat), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n589), .A2(new_n676), .A3(new_n387), .A4(new_n661), .ZN(new_n677));
  INV_X1    g476(.A(new_n536), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n668), .A2(new_n678), .A3(new_n669), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n679), .B2(new_n676), .ZN(G1326gat));
  NAND3_X1  g479(.A1(new_n589), .A2(new_n537), .A3(new_n661), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NOR2_X1   g482(.A1(new_n637), .A2(new_n656), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n619), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n589), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(G29gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n688), .A3(new_n664), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n255), .B1(new_n247), .B2(new_n252), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n619), .B1(new_n532), .B2(new_n578), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT105), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n697), .B(KEYINPUT44), .C1(new_n586), .C2(new_n619), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n438), .B1(new_n582), .B2(new_n583), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n548), .A2(new_n552), .A3(new_n503), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n553), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n517), .A3(new_n555), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n438), .B1(new_n478), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n574), .A2(new_n521), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n678), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n700), .A2(new_n706), .A3(KEYINPUT106), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n576), .B2(new_n577), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n532), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n712), .B(new_n532), .C1(new_n707), .C2(new_n709), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n619), .A2(KEYINPUT44), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n693), .B1(new_n699), .B2(new_n715), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n716), .A2(new_n664), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n690), .B1(new_n688), .B2(new_n717), .ZN(G1328gat));
  INV_X1    g517(.A(G36gat), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n687), .A2(new_n719), .A3(new_n540), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n716), .A2(new_n540), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n722), .B(new_n723), .C1(new_n719), .C2(new_n724), .ZN(G1329gat));
  INV_X1    g524(.A(G43gat), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n716), .B2(new_n536), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n687), .A2(new_n726), .A3(new_n387), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT47), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n727), .B2(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1330gat));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n736));
  INV_X1    g535(.A(G50gat), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n716), .B2(new_n537), .ZN(new_n738));
  AND4_X1   g537(.A1(new_n737), .A2(new_n589), .A3(new_n537), .A4(new_n686), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n735), .B(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n699), .A2(new_n715), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n537), .A3(new_n692), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G50gat), .ZN(new_n743));
  INV_X1    g542(.A(new_n739), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n743), .A2(KEYINPUT108), .A3(new_n734), .A4(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n740), .A2(new_n745), .ZN(G1331gat));
  AND2_X1   g545(.A1(new_n711), .A2(new_n713), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n615), .A2(new_n618), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n253), .A2(new_n256), .ZN(new_n749));
  INV_X1    g548(.A(new_n637), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n657), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n664), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n540), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT49), .B(G64gat), .Z(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n755), .B2(new_n757), .ZN(G1333gat));
  NAND3_X1  g557(.A1(new_n747), .A2(new_n387), .A3(new_n751), .ZN(new_n759));
  INV_X1    g558(.A(G71gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n678), .A2(new_n760), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n711), .A2(new_n713), .A3(new_n751), .A4(new_n762), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1334gat));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n537), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT111), .B(G78gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1335gat));
  NOR3_X1   g570(.A1(new_n619), .A2(new_n749), .A3(new_n637), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n710), .A2(KEYINPUT51), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT51), .B1(new_n710), .B2(new_n772), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n657), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n591), .A3(new_n664), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n750), .A2(new_n691), .A3(new_n656), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n699), .B2(new_n715), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n664), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n777), .B1(new_n780), .B2(new_n591), .ZN(G1336gat));
  AOI21_X1  g580(.A(new_n592), .B1(new_n779), .B2(new_n540), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n540), .A2(new_n592), .A3(new_n656), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT112), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n773), .B2(new_n774), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n782), .A2(KEYINPUT52), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT52), .B1(new_n782), .B2(new_n786), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1337gat));
  AND2_X1   g588(.A1(new_n779), .A2(new_n536), .ZN(new_n790));
  OAI21_X1  g589(.A(G99gat), .B1(new_n790), .B2(KEYINPUT113), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n779), .A2(KEYINPUT113), .A3(new_n536), .ZN(new_n792));
  INV_X1    g591(.A(G99gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n656), .A2(new_n793), .A3(new_n387), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT114), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n791), .A2(new_n792), .B1(new_n775), .B2(new_n795), .ZN(G1338gat));
  NOR2_X1   g595(.A1(new_n438), .A2(G106gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(G106gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n779), .B2(new_n537), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT53), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n779), .A2(new_n537), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n803), .B(new_n798), .C1(new_n804), .C2(new_n800), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(G1339gat));
  OAI21_X1  g605(.A(new_n228), .B1(new_n231), .B2(new_n233), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(G229gat), .A3(G233gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n239), .B2(new_n240), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n255), .B1(new_n251), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n656), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n638), .C1(new_n644), .C2(new_n645), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n652), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n646), .A2(KEYINPUT54), .ZN(new_n815));
  OR3_X1    g614(.A1(new_n644), .A2(new_n638), .A3(new_n645), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n653), .B1(new_n817), .B2(KEYINPUT55), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(KEYINPUT54), .A3(new_n646), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n821), .B2(new_n814), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n811), .B1(new_n823), .B2(new_n691), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n619), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n823), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n748), .A2(new_n810), .A3(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n828), .A2(new_n637), .B1(new_n749), .B2(new_n658), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n440), .ZN(new_n830));
  INV_X1    g629(.A(new_n664), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n540), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n749), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n587), .A2(new_n262), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n833), .B2(new_n835), .ZN(G1340gat));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n656), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g637(.A1(new_n833), .A2(new_n637), .ZN(new_n839));
  XNOR2_X1  g638(.A(KEYINPUT115), .B(G127gat), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n839), .B(new_n840), .ZN(G1342gat));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n619), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n830), .A2(new_n832), .A3(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT116), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(KEYINPUT116), .ZN(new_n846));
  AND4_X1   g645(.A1(new_n842), .A2(new_n845), .A3(new_n269), .A4(new_n846), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n845), .A2(new_n846), .B1(new_n842), .B2(new_n269), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(G1343gat));
  XOR2_X1   g648(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n850));
  NAND2_X1  g649(.A1(new_n678), .A2(new_n537), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT118), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n829), .A2(new_n832), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n259), .A2(new_n388), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n831), .A2(new_n540), .A3(new_n536), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n658), .A2(new_n749), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n820), .A2(KEYINPUT55), .A3(new_n652), .A4(new_n813), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n654), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n817), .B2(KEYINPUT55), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT117), .B(new_n819), .C1(new_n821), .C2(new_n814), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n259), .A2(new_n863), .B1(new_n656), .B2(new_n810), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n827), .B1(new_n864), .B2(new_n748), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n857), .B1(new_n865), .B2(new_n750), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n866), .A2(new_n867), .A3(new_n438), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n829), .B2(new_n537), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n259), .B(new_n856), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n855), .B1(new_n870), .B2(G141gat), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(KEYINPUT120), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n873), .B(new_n855), .C1(new_n870), .C2(G141gat), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n853), .A2(new_n854), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n749), .B(new_n856), .C1(new_n868), .C2(new_n869), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(G141gat), .ZN(new_n878));
  OAI22_X1  g677(.A1(new_n872), .A2(new_n874), .B1(new_n875), .B2(new_n878), .ZN(G1344gat));
  NOR3_X1   g678(.A1(new_n853), .A2(G148gat), .A3(new_n657), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n856), .B1(new_n868), .B2(new_n869), .ZN(new_n881));
  OAI21_X1  g680(.A(G148gat), .B1(new_n881), .B2(new_n657), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n856), .A2(new_n656), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n749), .A2(KEYINPUT95), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n691), .A2(new_n203), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n863), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n748), .B1(new_n889), .B2(new_n811), .ZN(new_n890));
  INV_X1    g689(.A(new_n827), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(KEYINPUT122), .B(new_n827), .C1(new_n864), .C2(new_n748), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(new_n750), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n659), .A2(new_n587), .A3(new_n660), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n537), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n867), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n829), .A2(new_n899), .A3(KEYINPUT57), .A4(new_n537), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n637), .B1(new_n825), .B2(new_n827), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT57), .B(new_n537), .C1(new_n857), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT121), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n885), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n884), .B1(new_n905), .B2(new_n906), .ZN(G1345gat));
  OAI21_X1  g706(.A(G155gat), .B1(new_n881), .B2(new_n750), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n750), .A2(G155gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n853), .B2(new_n909), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n881), .B2(new_n619), .ZN(new_n911));
  OR3_X1    g710(.A1(new_n853), .A2(G162gat), .A3(new_n619), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT123), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n664), .A2(new_n478), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n830), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n587), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n829), .A2(new_n831), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT124), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n439), .A2(new_n478), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n749), .A2(new_n329), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(G1348gat));
  OAI21_X1  g725(.A(G176gat), .B1(new_n919), .B2(new_n657), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n657), .A2(G176gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n924), .B2(new_n928), .ZN(G1349gat));
  NOR2_X1   g728(.A1(new_n750), .A2(new_n307), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n922), .A2(new_n923), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n354), .B1(new_n919), .B2(new_n750), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT60), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n931), .A2(new_n935), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n919), .B2(new_n619), .ZN(new_n938));
  XNOR2_X1  g737(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n938), .A2(new_n940), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n748), .A2(new_n305), .ZN(new_n943));
  OAI22_X1  g742(.A1(new_n941), .A2(new_n942), .B1(new_n924), .B2(new_n943), .ZN(G1351gat));
  NAND2_X1  g743(.A1(new_n918), .A2(new_n678), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT126), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n898), .B2(new_n904), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(G197gat), .A3(new_n259), .ZN(new_n948));
  INV_X1    g747(.A(G197gat), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n851), .A2(new_n478), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n922), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n949), .B1(new_n951), .B2(new_n691), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n948), .A2(new_n952), .ZN(G1352gat));
  NAND2_X1  g752(.A1(new_n947), .A2(new_n656), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G204gat), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n657), .A2(G204gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n922), .A2(new_n950), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(G1353gat));
  INV_X1    g759(.A(new_n946), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT57), .B1(new_n896), .B2(new_n537), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n900), .A2(new_n903), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n637), .B(new_n961), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n637), .A2(new_n401), .ZN(new_n967));
  OAI22_X1  g766(.A1(new_n965), .A2(new_n966), .B1(new_n951), .B2(new_n967), .ZN(G1354gat));
  AND2_X1   g767(.A1(new_n947), .A2(new_n748), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n748), .A2(new_n402), .ZN(new_n970));
  OAI22_X1  g769(.A1(new_n969), .A2(new_n402), .B1(new_n951), .B2(new_n970), .ZN(G1355gat));
endmodule


