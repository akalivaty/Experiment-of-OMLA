//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT83), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  OAI21_X1  g003(.A(G210), .B1(G237), .B2(G902), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT0), .B(G128), .Z(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT64), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT0), .A4(G128), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n191), .A2(new_n200), .A3(new_n196), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n196), .A2(new_n204), .A3(G128), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n193), .B(new_n195), .C1(KEYINPUT1), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT86), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT86), .ZN(new_n211));
  AOI211_X1 g025(.A(new_n211), .B(G125), .C1(new_n205), .C2(new_n207), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n203), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G224), .ZN(new_n215));
  XOR2_X1   g029(.A(new_n215), .B(KEYINPUT87), .Z(new_n216));
  XNOR2_X1  g030(.A(new_n213), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT5), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G116), .ZN(new_n221));
  XNOR2_X1  g035(.A(G116), .B(G119), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI211_X1 g037(.A(G113), .B(new_n221), .C1(new_n223), .C2(new_n219), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT2), .A2(G113), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT65), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT2), .A3(G113), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT2), .A2(G113), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AND4_X1   g046(.A1(new_n225), .A2(new_n230), .A3(new_n232), .A4(new_n222), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n231), .B1(new_n227), .B2(new_n229), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n225), .B1(new_n234), .B2(new_n222), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n224), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G107), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT81), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(KEYINPUT81), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n238), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G101), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n237), .A2(G107), .ZN(new_n245));
  INV_X1    g059(.A(G107), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G104), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n239), .B2(KEYINPUT3), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n245), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G101), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT84), .B1(new_n236), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n249), .A2(new_n251), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT84), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n230), .A2(new_n232), .A3(new_n222), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n234), .A2(new_n225), .A3(new_n222), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n254), .A2(new_n255), .A3(new_n259), .A4(new_n224), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n248), .B(new_n245), .C1(new_n262), .C2(new_n247), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G101), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT4), .A3(new_n249), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n266), .A3(G101), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n228), .B1(KEYINPUT2), .B2(G113), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n226), .A2(KEYINPUT65), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n232), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT66), .A3(new_n223), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n234), .B2(new_n222), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n259), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n259), .B2(new_n275), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n268), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G110), .B(G122), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n261), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n261), .A2(new_n279), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n280), .B(KEYINPUT85), .Z(new_n283));
  AOI22_X1  g097(.A1(new_n281), .A2(KEYINPUT6), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n265), .A2(new_n267), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT66), .B1(new_n271), .B2(new_n223), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n234), .A2(new_n273), .A3(new_n222), .ZN(new_n287));
  OAI22_X1  g101(.A1(new_n286), .A2(new_n287), .B1(new_n233), .B2(new_n235), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT68), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n259), .A2(new_n275), .A3(new_n276), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n285), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n253), .A2(new_n260), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT6), .B(new_n283), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n218), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT88), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n283), .B1(new_n291), .B2(new_n292), .ZN(new_n297));
  INV_X1    g111(.A(new_n280), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n291), .A2(new_n292), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT6), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n293), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT88), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(new_n218), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n215), .A2(KEYINPUT7), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n210), .B2(new_n212), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n203), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n210), .A2(new_n212), .A3(new_n308), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT90), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  OR3_X1    g128(.A1(new_n213), .A2(KEYINPUT91), .A3(new_n307), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n236), .B(new_n252), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n280), .B(KEYINPUT8), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT91), .B1(new_n213), .B2(new_n307), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n281), .A2(new_n315), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n306), .B1(new_n314), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n190), .B1(new_n305), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n190), .ZN(new_n324));
  AOI211_X1 g138(.A(new_n324), .B(new_n321), .C1(new_n296), .C2(new_n304), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n189), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n205), .A2(new_n207), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT11), .ZN(new_n328));
  INV_X1    g142(.A(G134), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(G137), .ZN(new_n330));
  INV_X1    g144(.A(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT11), .A3(G134), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n334), .A2(G131), .ZN(new_n335));
  INV_X1    g149(.A(new_n333), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n329), .A2(G137), .ZN(new_n337));
  OAI21_X1  g151(.A(G131), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n327), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G131), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n334), .B(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n339), .B1(new_n202), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT30), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n289), .A2(new_n290), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n342), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n277), .A2(new_n278), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT69), .B1(new_n289), .B2(new_n290), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G237), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(new_n214), .A3(G210), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n353), .B(KEYINPUT27), .Z(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT26), .B(G101), .ZN(new_n355));
  XOR2_X1   g169(.A(new_n354), .B(new_n355), .Z(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT31), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT31), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n345), .A2(new_n359), .A3(new_n350), .A4(new_n356), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n342), .B(KEYINPUT71), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n347), .B1(new_n277), .B2(new_n278), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n289), .A2(KEYINPUT69), .A3(new_n290), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT28), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n342), .B1(new_n277), .B2(new_n278), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT70), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n344), .A2(KEYINPUT70), .A3(new_n342), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n350), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n366), .B1(new_n371), .B2(KEYINPUT28), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT72), .B1(new_n372), .B2(new_n356), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n370), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n342), .B1(new_n363), .B2(new_n364), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT28), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n362), .A2(new_n365), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT28), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT72), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n357), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n361), .B1(new_n373), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(G472), .A2(G902), .ZN(new_n384));
  XOR2_X1   g198(.A(new_n384), .B(KEYINPUT73), .Z(new_n385));
  OAI21_X1  g199(.A(KEYINPUT32), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n358), .A2(new_n360), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n381), .B1(new_n380), .B2(new_n357), .ZN(new_n388));
  AOI211_X1 g202(.A(KEYINPUT72), .B(new_n356), .C1(new_n376), .C2(new_n379), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT32), .ZN(new_n391));
  INV_X1    g205(.A(new_n385), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n351), .B2(new_n357), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n380), .B2(new_n357), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n365), .B(new_n346), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n366), .B1(new_n397), .B2(KEYINPUT28), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n356), .A2(KEYINPUT29), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n399), .B1(new_n398), .B2(new_n401), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n306), .B(new_n396), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G472), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n326), .B1(new_n394), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n254), .A2(KEYINPUT10), .A3(new_n327), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n252), .B2(new_n208), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n411));
  INV_X1    g225(.A(new_n202), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n265), .A3(new_n267), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n410), .A2(new_n411), .A3(new_n341), .A4(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n413), .A2(new_n341), .A3(new_n409), .A4(new_n407), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT82), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n334), .B(G131), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n254), .A2(new_n327), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n252), .A2(new_n208), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT12), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(KEYINPUT12), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G140), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n214), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n414), .B2(new_n416), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n410), .A2(new_n413), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n418), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n426), .A2(new_n429), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G469), .B1(new_n433), .B2(G902), .ZN(new_n434));
  INV_X1    g248(.A(G469), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n430), .A2(new_n425), .ZN(new_n436));
  INV_X1    g250(.A(new_n429), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n417), .B2(new_n432), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n435), .B(new_n306), .C1(new_n436), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G217), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(G234), .B2(new_n306), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G902), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n220), .A2(G128), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n445), .A2(KEYINPUT23), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n206), .A2(G119), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT76), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT76), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(KEYINPUT23), .ZN(new_n450));
  OAI22_X1  g264(.A1(new_n446), .A2(new_n448), .B1(new_n450), .B2(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G110), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT77), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G125), .B(G140), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT16), .ZN(new_n456));
  OR3_X1    g270(.A1(new_n209), .A2(KEYINPUT16), .A3(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n192), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(G146), .A3(new_n457), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n447), .A2(new_n445), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT24), .B(G110), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT75), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n454), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n463), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT78), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(G110), .B2(new_n451), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n455), .A2(new_n192), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n460), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT22), .B(G137), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n466), .A2(new_n471), .A3(new_n475), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT79), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT79), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n444), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n306), .A3(new_n478), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT25), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n483), .B1(new_n486), .B2(new_n442), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT9), .B(G234), .ZN(new_n488));
  OAI21_X1  g302(.A(G221), .B1(new_n488), .B2(G902), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT80), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n440), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n352), .A2(new_n214), .A3(G214), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n194), .A2(KEYINPUT92), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n194), .A2(KEYINPUT92), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n494), .A2(G214), .A3(new_n352), .A4(new_n214), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(KEYINPUT18), .A2(G131), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT93), .B1(new_n455), .B2(new_n192), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n192), .B2(new_n455), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n497), .A2(new_n500), .A3(new_n498), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n506));
  OR3_X1    g320(.A1(new_n455), .A2(new_n506), .A3(new_n192), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n502), .A2(new_n504), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n497), .A2(new_n340), .A3(new_n498), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n340), .B1(new_n497), .B2(new_n498), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT19), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n455), .B(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n460), .B1(new_n514), .B2(G146), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n508), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G113), .B(G122), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(new_n237), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n510), .A2(KEYINPUT17), .A3(new_n511), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n499), .A2(KEYINPUT17), .A3(G131), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n460), .A3(new_n459), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n518), .B(new_n508), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT94), .ZN(new_n526));
  NOR2_X1   g340(.A1(G475), .A2(G902), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n520), .A2(new_n528), .A3(new_n524), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n527), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(KEYINPUT20), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n530), .A2(KEYINPUT20), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G475), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n521), .A2(new_n523), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n518), .B1(new_n535), .B2(new_n508), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT95), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n524), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(G902), .B1(new_n536), .B2(KEYINPUT95), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n534), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(G116), .B(G122), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n543), .A2(new_n246), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n194), .A2(G128), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n206), .A2(G143), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n329), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G134), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n544), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G116), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(KEYINPUT14), .A3(G122), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G107), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT14), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n554), .B2(new_n543), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n550), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n488), .A2(new_n441), .A3(G953), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT97), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT13), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n545), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n546), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n545), .A2(new_n563), .ZN(new_n566));
  OAI21_X1  g380(.A(G134), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n543), .A2(new_n246), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n567), .B(new_n547), .C1(new_n568), .C2(new_n544), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n559), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n562), .B1(new_n559), .B2(new_n569), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G478), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n306), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n306), .B1(new_n571), .B2(new_n572), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n575), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G952), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G953), .ZN(new_n582));
  INV_X1    g396(.A(G234), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n582), .B1(new_n583), .B2(new_n352), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI211_X1 g399(.A(new_n306), .B(new_n214), .C1(G234), .C2(G237), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT21), .B(G898), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR4_X1   g402(.A1(new_n533), .A2(new_n542), .A3(new_n580), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n492), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n406), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  AOI21_X1  g407(.A(new_n303), .B1(new_n302), .B2(new_n218), .ZN(new_n594));
  AOI211_X1 g408(.A(KEYINPUT88), .B(new_n217), .C1(new_n301), .C2(new_n293), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n322), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n324), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n190), .B(new_n322), .C1(new_n594), .C2(new_n595), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n188), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n588), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n574), .A2(new_n306), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n578), .B2(G478), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT33), .B1(new_n572), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n573), .B(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n603), .B1(new_n606), .B2(G478), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n533), .A2(new_n542), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n599), .A2(new_n600), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G472), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n390), .B2(new_n306), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n383), .A2(new_n385), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n613), .A2(new_n492), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  AND3_X1   g432(.A1(new_n520), .A2(new_n528), .A3(new_n524), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n528), .B1(new_n520), .B2(new_n524), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n619), .A2(new_n620), .A3(new_n531), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT20), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT99), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n530), .A2(new_n624), .A3(KEYINPUT20), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n526), .A2(new_n529), .A3(new_n532), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n623), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n535), .A2(new_n508), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(KEYINPUT95), .A3(new_n519), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n306), .ZN(new_n631));
  OAI21_X1  g445(.A(G475), .B1(new_n631), .B2(new_n539), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n580), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n628), .A2(new_n634), .A3(new_n600), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n530), .A2(KEYINPUT20), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n626), .B1(new_n638), .B2(KEYINPUT99), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n633), .B1(new_n639), .B2(new_n625), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(KEYINPUT100), .A3(new_n600), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n326), .A2(new_n642), .A3(KEYINPUT101), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT100), .B1(new_n640), .B2(new_n600), .ZN(new_n645));
  AND4_X1   g459(.A1(KEYINPUT100), .A2(new_n628), .A3(new_n600), .A4(new_n634), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n644), .B1(new_n647), .B2(new_n599), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n615), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NAND2_X1  g465(.A1(new_n486), .A2(new_n442), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n476), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT102), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n472), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n443), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n657), .A2(new_n440), .A3(new_n491), .A4(new_n589), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n326), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n613), .A2(new_n614), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT103), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT37), .B(G110), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  NAND3_X1  g478(.A1(new_n657), .A2(new_n440), .A3(new_n491), .ZN(new_n665));
  INV_X1    g479(.A(new_n586), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n584), .B1(new_n666), .B2(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n640), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n406), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  NAND2_X1  g485(.A1(new_n351), .A2(new_n356), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n672), .B(new_n306), .C1(new_n356), .C2(new_n397), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n394), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n657), .ZN(new_n676));
  INV_X1    g490(.A(new_n580), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n609), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n675), .A2(new_n189), .A3(new_n676), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n597), .A2(new_n598), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT38), .Z(new_n681));
  OR2_X1    g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n667), .B(KEYINPUT39), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AOI211_X1 g500(.A(new_n490), .B(new_n686), .C1(new_n434), .C2(new_n439), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT40), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n688), .B1(new_n682), .B2(new_n683), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n194), .ZN(G45));
  INV_X1    g505(.A(new_n609), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n607), .A3(new_n667), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n665), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n406), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  INV_X1    g510(.A(new_n487), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n394), .B2(new_n405), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n417), .A2(new_n432), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n699), .A2(new_n429), .B1(new_n430), .B2(new_n425), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n439), .A3(new_n489), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n611), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  OAI211_X1 g520(.A(new_n698), .B(new_n703), .C1(new_n643), .C2(new_n648), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NAND2_X1  g522(.A1(new_n394), .A2(new_n405), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n676), .A2(new_n590), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n188), .B(new_n702), .C1(new_n597), .C2(new_n598), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  XNOR2_X1  g527(.A(KEYINPUT105), .B(G472), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n390), .B2(new_n306), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n398), .A2(new_n356), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n385), .B1(new_n717), .B2(new_n387), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n716), .A2(new_n697), .A3(new_n718), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n188), .B(new_n588), .C1(new_n597), .C2(new_n598), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n678), .A4(new_n703), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NOR4_X1   g536(.A1(new_n716), .A2(new_n676), .A3(new_n718), .A4(new_n693), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n711), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(new_n693), .ZN(new_n726));
  INV_X1    g540(.A(new_n489), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n434), .B2(new_n439), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n597), .A2(new_n728), .A3(new_n189), .A4(new_n598), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n698), .B(new_n726), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n729), .B(new_n730), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(KEYINPUT42), .A3(new_n726), .A4(new_n698), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  INV_X1    g553(.A(new_n668), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n698), .B(new_n740), .C1(new_n731), .C2(new_n732), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  NOR2_X1   g556(.A1(new_n660), .A2(new_n676), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n743), .B(KEYINPUT107), .Z(new_n744));
  NAND2_X1  g558(.A1(new_n609), .A2(new_n607), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT43), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT44), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n597), .A2(new_n189), .A3(new_n598), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n433), .A2(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n433), .A2(KEYINPUT45), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(G469), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(G469), .A2(G902), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n754), .A2(KEYINPUT46), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n753), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n439), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n489), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n748), .A2(new_n686), .A3(new_n749), .A4(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n744), .A2(KEYINPUT44), .A3(new_n747), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  XNOR2_X1  g576(.A(new_n758), .B(KEYINPUT47), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n709), .A2(new_n487), .A3(new_n693), .A4(new_n749), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n763), .B1(KEYINPUT108), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(KEYINPUT108), .B2(new_n764), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  NAND3_X1  g581(.A1(new_n394), .A2(new_n487), .A3(new_n674), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n749), .A2(new_n584), .A3(new_n702), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT114), .Z(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n610), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n698), .A2(new_n747), .A3(new_n770), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT48), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n719), .A2(new_n585), .A3(new_n747), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n711), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n773), .A2(new_n582), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n772), .A2(new_n609), .A3(new_n608), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT115), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n770), .A2(new_n747), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n781), .A2(new_n676), .A3(new_n718), .A4(new_n716), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n776), .A2(new_n681), .A3(new_n188), .A4(new_n703), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT113), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n783), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n701), .A2(new_n439), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n763), .B1(new_n491), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n749), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n776), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT112), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n782), .B(new_n786), .C1(new_n788), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n780), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n778), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n780), .A2(new_n792), .A3(KEYINPUT51), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT116), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n406), .B1(new_n669), .B2(new_n694), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n680), .A2(new_n189), .A3(new_n678), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n676), .A2(new_n728), .A3(new_n667), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n675), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n724), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT110), .B1(new_n804), .B2(KEYINPUT111), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(KEYINPUT52), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n805), .B2(KEYINPUT52), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n723), .B1(new_n731), .B2(new_n732), .ZN(new_n809));
  INV_X1    g623(.A(new_n628), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n677), .A2(new_n632), .A3(new_n667), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n665), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n709), .A2(new_n789), .A3(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n741), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n738), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n609), .A2(new_n607), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n609), .B2(new_n677), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n615), .A2(new_n720), .A3(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n721), .A2(new_n712), .A3(new_n818), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n406), .A2(new_n591), .B1(new_n659), .B2(new_n660), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n704), .A3(new_n707), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n815), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n741), .A2(new_n809), .A3(new_n813), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n735), .B2(new_n737), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n707), .A2(new_n820), .A3(new_n704), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n721), .A2(new_n712), .A3(new_n818), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT109), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  OAI221_X1 g643(.A(new_n799), .B1(new_n806), .B2(new_n808), .C1(new_n823), .C2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n804), .B(KEYINPUT52), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n823), .B2(new_n829), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n831), .B1(KEYINPUT53), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT54), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n815), .A2(new_n821), .A3(new_n799), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(new_n806), .B2(new_n808), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n822), .B1(new_n815), .B2(new_n821), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n825), .A2(new_n828), .A3(KEYINPUT109), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n832), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n837), .B(new_n839), .C1(new_n842), .C2(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n836), .A2(new_n843), .ZN(new_n844));
  OAI22_X1  g658(.A1(new_n798), .A2(new_n844), .B1(G952), .B2(G953), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n787), .A2(KEYINPUT49), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n787), .A2(KEYINPUT49), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n491), .A2(new_n189), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n846), .A2(new_n847), .A3(new_n745), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n681), .A2(new_n769), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n845), .A2(new_n850), .ZN(G75));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n302), .B(new_n218), .ZN(new_n853));
  XNOR2_X1  g667(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n839), .B1(new_n842), .B2(KEYINPUT53), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(G902), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT119), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n852), .B(new_n855), .C1(new_n858), .C2(new_n190), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n214), .A2(G952), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n856), .A2(G210), .A3(G902), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n855), .B1(new_n862), .B2(new_n852), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n859), .B(new_n861), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(G51));
  NOR2_X1   g682(.A1(new_n857), .A2(KEYINPUT119), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n856), .B2(G902), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n869), .A2(new_n752), .A3(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n753), .B(KEYINPUT57), .Z(new_n873));
  NAND2_X1  g687(.A1(new_n834), .A2(new_n799), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n837), .B1(new_n874), .B2(new_n839), .ZN(new_n875));
  INV_X1    g689(.A(new_n843), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n700), .B1(new_n877), .B2(KEYINPUT120), .ZN(new_n878));
  INV_X1    g692(.A(new_n873), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n856), .A2(KEYINPUT54), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(new_n843), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n872), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT121), .B1(new_n884), .B2(new_n860), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n881), .A2(new_n882), .B1(new_n438), .B2(new_n436), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n877), .A2(KEYINPUT120), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n886), .A2(new_n887), .B1(new_n752), .B2(new_n858), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n861), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n890), .ZN(G54));
  NOR2_X1   g705(.A1(new_n869), .A2(new_n871), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n620), .B2(new_n619), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n619), .A2(new_n620), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .A4(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n894), .A2(new_n861), .A3(new_n896), .ZN(G60));
  XNOR2_X1  g711(.A(new_n606), .B(KEYINPUT122), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n601), .B(KEYINPUT59), .Z(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n844), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n880), .B2(new_n843), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n860), .A3(new_n902), .ZN(G63));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT60), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n874), .B2(new_n839), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n480), .A2(new_n482), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n861), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n911), .B2(new_n904), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n907), .A2(new_n655), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n911), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n913), .B(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n912), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n914), .B1(new_n915), .B2(new_n918), .ZN(G66));
  XNOR2_X1  g733(.A(new_n828), .B(KEYINPUT125), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n214), .ZN(new_n921));
  INV_X1    g735(.A(G224), .ZN(new_n922));
  OAI21_X1  g736(.A(G953), .B1(new_n587), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n301), .B(new_n293), .C1(G898), .C2(new_n214), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(G69));
  NAND2_X1  g740(.A1(G900), .A2(G953), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n800), .A2(new_n724), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n766), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n741), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n758), .A2(new_n686), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n698), .A2(new_n801), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n929), .A2(new_n761), .A3(new_n738), .A4(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n927), .B1(new_n934), .B2(G953), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n343), .B(new_n514), .Z(new_n936));
  NAND4_X1  g750(.A1(new_n698), .A2(new_n687), .A3(new_n789), .A4(new_n817), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n766), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n928), .B1(new_n684), .B2(new_n689), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n938), .A2(new_n761), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n936), .A2(G953), .ZN(new_n943));
  AOI22_X1  g757(.A1(new_n935), .A2(new_n936), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n214), .B1(G227), .B2(G900), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G72));
  XNOR2_X1  g760(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n612), .A2(new_n306), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n934), .B2(new_n920), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n351), .A2(new_n356), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n860), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n951), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n835), .A2(new_n672), .A3(new_n953), .A4(new_n949), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n949), .B1(new_n942), .B2(new_n920), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n351), .A3(new_n356), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n952), .A2(new_n954), .A3(new_n956), .ZN(G57));
endmodule


