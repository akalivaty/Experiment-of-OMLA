//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n452), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT70), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(new_n466), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(G125), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  XOR2_X1   g048(.A(new_n473), .B(KEYINPUT71), .Z(new_n474));
  AOI21_X1  g049(.A(new_n464), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n464), .A2(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(new_n469), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G160));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n464), .C2(G112), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT72), .Z(new_n483));
  OAI21_X1  g058(.A(new_n467), .B1(new_n463), .B2(new_n462), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n469), .A2(G2105), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n485), .A2(G124), .B1(G136), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n483), .A2(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n467), .A2(new_n489), .A3(G126), .A4(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT73), .B1(new_n469), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g068(.A1(KEYINPUT74), .A2(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT74), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n464), .A2(G138), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(new_n467), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n500), .A2(new_n468), .A3(new_n471), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n515), .A2(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n513), .A2(new_n523), .ZN(G166));
  NOR2_X1   g099(.A1(new_n518), .A2(new_n517), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n514), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  INV_X1    g105(.A(new_n520), .ZN(new_n531));
  NAND2_X1  g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n533), .A2(G51), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n529), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  OAI21_X1  g114(.A(G64), .B1(new_n518), .B2(new_n517), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n512), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n533), .A2(G52), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n510), .A2(new_n514), .A3(G90), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n546), .B(new_n547), .C1(new_n542), .C2(new_n543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n512), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n515), .A2(new_n552), .B1(new_n521), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n515), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n533), .A2(new_n563), .A3(G53), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n512), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n521), .A2(KEYINPUT77), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n510), .A2(new_n514), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(G91), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n565), .A2(new_n567), .A3(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G166), .ZN(G303));
  AND2_X1   g149(.A1(new_n568), .A2(new_n570), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G87), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n510), .A2(G74), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(new_n533), .B2(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(new_n575), .A2(G86), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n512), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n533), .A2(G48), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n580), .A2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n512), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n515), .A2(new_n589), .B1(new_n521), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  OR3_X1    g169(.A1(G171), .A2(KEYINPUT78), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT78), .B1(G171), .B2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n508), .B2(new_n509), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n533), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n568), .A2(G92), .A3(new_n570), .ZN(new_n605));
  XNOR2_X1  g180(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n568), .A2(G92), .A3(new_n570), .A4(new_n606), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n604), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n595), .B(new_n596), .C1(G868), .C2(new_n610), .ZN(G284));
  OAI211_X1 g186(.A(new_n595), .B(new_n596), .C1(G868), .C2(new_n610), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(new_n555), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n594), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n608), .A2(new_n609), .ZN(new_n621));
  INV_X1    g196(.A(new_n604), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n620), .B1(new_n624), .B2(new_n594), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g201(.A1(new_n468), .A2(new_n471), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n477), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n485), .A2(G123), .B1(G135), .B2(new_n486), .ZN(new_n634));
  OAI221_X1 g209(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT81), .ZN(G156));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT82), .Z(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n641), .B2(new_n642), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT83), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  INV_X1    g241(.A(new_n659), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n666), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT85), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n673), .A2(new_n676), .A3(new_n679), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1981), .B(G1986), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(G6), .ZN(new_n696));
  INV_X1    g271(.A(G305), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n690), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  OR2_X1    g275(.A1(new_n690), .A2(KEYINPUT86), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n690), .A2(KEYINPUT86), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1971), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n695), .A2(new_n700), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n485), .A2(G119), .ZN(new_n713));
  OAI221_X1 g288(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n486), .A2(G131), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n712), .B1(new_n717), .B2(new_n711), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n703), .A2(G24), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n592), .B2(new_n703), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT87), .B(G1986), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n709), .A2(new_n710), .A3(new_n720), .A4(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT36), .Z(new_n726));
  NOR2_X1   g301(.A1(G162), .A2(new_n711), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n711), .B2(G35), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n729));
  INV_X1    g304(.A(G2090), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G164), .A2(new_n711), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G27), .B2(new_n711), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n728), .A2(new_n731), .B1(G2078), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n728), .B2(new_n731), .ZN(new_n736));
  INV_X1    g311(.A(G2078), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT31), .B(G11), .Z(new_n739));
  INV_X1    g314(.A(G28), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(KEYINPUT30), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT95), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n740), .B2(KEYINPUT30), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n703), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n555), .B2(new_n745), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n744), .B1(new_n636), .B2(new_n711), .C1(new_n747), .C2(G1341), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G1341), .B2(new_n747), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n690), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n690), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n738), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n486), .A2(G139), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT91), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT90), .B(KEYINPUT25), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n627), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n756), .B(new_n759), .C1(new_n760), .C2(new_n464), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(new_n711), .ZN(new_n762));
  NOR2_X1   g337(.A1(G29), .A2(G33), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT89), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G2072), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  NOR2_X1   g342(.A1(G171), .A2(new_n690), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G5), .B2(new_n690), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n766), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n610), .A2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G4), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1348), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR4_X1   g349(.A1(new_n736), .A2(new_n754), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n765), .A2(G2072), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT92), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n769), .A2(new_n767), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT24), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n711), .B1(new_n779), .B2(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n779), .B2(G34), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G160), .B2(G29), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n778), .B1(G2084), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G2084), .B2(new_n782), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n775), .A2(new_n777), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n485), .A2(G129), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT93), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n486), .A2(G141), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT26), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n477), .A2(G105), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n787), .A2(new_n788), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G32), .B(new_n792), .S(G29), .Z(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT94), .Z(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT27), .B(G1996), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n795), .A2(new_n796), .B1(new_n773), .B2(new_n772), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n745), .A2(G20), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT23), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n614), .B2(new_n690), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT97), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n711), .A2(G26), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT28), .ZN(new_n806));
  OAI221_X1 g381(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n486), .A2(G140), .ZN(new_n808));
  INV_X1    g383(.A(G128), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n484), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n810), .A2(KEYINPUT88), .A3(G29), .ZN(new_n811));
  AOI21_X1  g386(.A(KEYINPUT88), .B1(new_n810), .B2(G29), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n806), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G2067), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n797), .A2(new_n798), .A3(new_n804), .A4(new_n815), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n726), .A2(new_n785), .A3(new_n816), .ZN(G311));
  INV_X1    g392(.A(G311), .ZN(G150));
  NAND2_X1  g393(.A1(new_n533), .A2(G55), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n510), .A2(new_n514), .A3(G93), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n510), .A2(G67), .ZN(new_n822));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n512), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n610), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n619), .A2(new_n831), .A3(new_n825), .ZN(new_n832));
  INV_X1    g407(.A(new_n824), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n833), .A2(KEYINPUT99), .A3(new_n820), .A4(new_n819), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n831), .B1(new_n821), .B2(new_n824), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(new_n555), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n830), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n840), .B2(KEYINPUT39), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n827), .B1(new_n841), .B2(new_n843), .ZN(G145));
  AND3_X1   g419(.A1(new_n502), .A2(KEYINPUT100), .A3(new_n504), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT100), .B1(new_n502), .B2(new_n504), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n499), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n810), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n761), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n792), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n485), .A2(G130), .B1(G142), .B2(new_n486), .ZN(new_n851));
  OAI221_X1 g426(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n629), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n716), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(G160), .B(new_n636), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G162), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n855), .B(KEYINPUT101), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n856), .B(new_n859), .C1(new_n850), .C2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n850), .B(new_n860), .Z(new_n863));
  OAI211_X1 g438(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n859), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g440(.A1(new_n825), .A2(new_n594), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n610), .A2(KEYINPUT102), .A3(G299), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n621), .A2(G299), .A3(new_n622), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT102), .B1(new_n610), .B2(G299), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT41), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n623), .A2(new_n872), .A3(new_n614), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n610), .A2(G299), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AND4_X1   g451(.A1(new_n870), .A2(new_n873), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n870), .A3(new_n874), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n624), .B(new_n837), .Z(new_n881));
  MUX2_X1   g456(.A(new_n878), .B(new_n880), .S(new_n881), .Z(new_n882));
  XNOR2_X1  g457(.A(G288), .B(G303), .ZN(new_n883));
  XNOR2_X1  g458(.A(G305), .B(G290), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT42), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n882), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n866), .B1(new_n889), .B2(new_n594), .ZN(G295));
  OAI21_X1  g465(.A(new_n866), .B1(new_n889), .B2(new_n594), .ZN(G331));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n535), .A2(new_n536), .ZN(new_n893));
  INV_X1    g468(.A(G51), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n515), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT105), .B1(new_n895), .B2(new_n528), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n529), .A2(new_n537), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(G171), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g474(.A(G286), .B(KEYINPUT105), .C1(new_n545), .C2(new_n548), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n837), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n899), .A2(new_n832), .A3(new_n836), .A4(new_n900), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n892), .B(new_n904), .C1(new_n871), .C2(new_n877), .ZN(new_n905));
  AND4_X1   g480(.A1(new_n832), .A2(new_n899), .A3(new_n836), .A4(new_n900), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n900), .A2(new_n899), .B1(new_n832), .B2(new_n836), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n869), .A2(new_n870), .A3(new_n876), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n879), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n908), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT106), .B1(new_n904), .B2(new_n880), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n905), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n887), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n879), .B1(new_n908), .B2(new_n875), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n879), .B2(new_n910), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n904), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n879), .A2(new_n918), .A3(new_n910), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n887), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n916), .A2(new_n923), .A3(new_n862), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n925), .A2(KEYINPUT111), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n905), .B(new_n887), .C1(new_n912), .C2(new_n913), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n862), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT107), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n930), .A3(new_n862), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n916), .A3(new_n931), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n925), .A2(KEYINPUT111), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n926), .A2(new_n933), .A3(KEYINPUT44), .A4(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n936));
  XNOR2_X1  g511(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n931), .A2(new_n916), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n930), .B1(new_n927), .B2(new_n862), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  AND4_X1   g517(.A1(new_n942), .A2(new_n916), .A3(new_n862), .A4(new_n923), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n938), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT108), .B1(new_n932), .B2(KEYINPUT43), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n936), .B(new_n937), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n938), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n943), .B1(new_n932), .B2(KEYINPUT43), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(new_n950), .B2(new_n938), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n936), .B1(new_n951), .B2(new_n937), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n935), .B1(new_n948), .B2(new_n952), .ZN(G397));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n847), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G160), .A2(G40), .ZN(new_n958));
  OR3_X1    g533(.A1(new_n957), .A2(KEYINPUT112), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT112), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1996), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n792), .B(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n810), .B(new_n814), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n717), .A2(new_n719), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n717), .A2(new_n719), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1986), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n592), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n961), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n958), .B1(new_n955), .B2(new_n956), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n499), .B2(new_n505), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT45), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(G2078), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n506), .A2(new_n954), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n958), .B1(new_n977), .B2(new_n956), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n847), .A2(KEYINPUT45), .A3(new_n954), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n737), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n974), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n958), .B1(new_n977), .B2(KEYINPUT50), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n847), .A2(new_n983), .A3(new_n954), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n976), .B(new_n981), .C1(G1961), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G171), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n979), .A2(new_n975), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n971), .A2(new_n988), .B1(new_n980), .B2(new_n974), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT125), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n985), .B2(G1961), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n982), .A2(new_n984), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(KEYINPUT125), .A3(new_n767), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n989), .A2(new_n991), .A3(G301), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G303), .A2(G8), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1971), .B1(new_n978), .B2(new_n979), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n1002));
  OAI22_X1  g577(.A1(new_n1001), .A2(new_n1002), .B1(new_n992), .B2(G2090), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  OAI211_X1 g579(.A(G8), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G40), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n475), .A2(new_n1006), .A3(new_n480), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n847), .A2(new_n954), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G305), .A2(G1981), .ZN(new_n1009));
  INV_X1    g584(.A(G1981), .ZN(new_n1010));
  INV_X1    g585(.A(G86), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n583), .B1(new_n1011), .B2(new_n521), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(KEYINPUT115), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n582), .B1(new_n1012), .B2(KEYINPUT115), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1008), .B(G8), .C1(new_n1016), .C2(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(KEYINPUT116), .A3(KEYINPUT49), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n692), .A2(G1976), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1008), .A2(G8), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n692), .A2(G1976), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1024), .A2(KEYINPUT52), .A3(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1024), .A2(KEYINPUT52), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1022), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n983), .B1(new_n847), .B2(new_n954), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1007), .B1(new_n977), .B2(KEYINPUT50), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1029), .A2(new_n1030), .A3(G2090), .ZN(new_n1031));
  OAI21_X1  g606(.A(G8), .B1(new_n1031), .B2(new_n1001), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1000), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1005), .A2(new_n1028), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n997), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT54), .B1(new_n986), .B2(G171), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n988), .A2(new_n971), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n991), .A2(new_n981), .A3(new_n1038), .A4(new_n993), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G171), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT126), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(KEYINPUT126), .A3(G171), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1037), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1036), .A2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT56), .B(G2072), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n978), .A2(new_n979), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT100), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n505), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n502), .A2(KEYINPUT100), .A3(new_n504), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n498), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT50), .B1(new_n1052), .B2(G1384), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n958), .B1(new_n983), .B2(new_n972), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1956), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT119), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n803), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n1047), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n1061));
  OAI21_X1  g636(.A(G299), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1056), .A2(new_n1059), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1348), .B1(new_n982), .B2(new_n984), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1008), .A2(G2067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1066), .B1(new_n623), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1057), .A2(new_n1047), .A3(new_n1064), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1066), .A2(KEYINPUT61), .A3(new_n1071), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n978), .A2(new_n979), .A3(new_n962), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT58), .B(G1341), .Z(new_n1075));
  NAND2_X1  g650(.A1(new_n1008), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n619), .B1(KEYINPUT120), .B2(KEYINPUT59), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1081), .A2(new_n1082), .B1(KEYINPUT120), .B2(KEYINPUT59), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n623), .B1(new_n1069), .B2(KEYINPUT60), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n1085));
  NOR4_X1   g660(.A1(new_n1067), .A2(new_n1068), .A3(new_n1085), .A4(new_n610), .ZN(new_n1086));
  OAI22_X1  g661(.A1(new_n1084), .A2(new_n1086), .B1(KEYINPUT60), .B2(new_n1069), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1082), .ZN(new_n1088));
  NOR2_X1   g663(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1080), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1073), .A2(new_n1083), .A3(new_n1087), .A4(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1065), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT61), .B1(new_n1092), .B2(new_n1071), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT122), .B(KEYINPUT61), .C1(new_n1092), .C2(new_n1071), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1072), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n957), .A2(new_n1007), .A3(new_n973), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n752), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n992), .A2(G2084), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(KEYINPUT123), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1966), .B1(new_n971), .B2(new_n973), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n992), .A2(G2084), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G8), .ZN(new_n1108));
  NOR2_X1   g683(.A1(G168), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(G8), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1109), .B(KEYINPUT124), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1115));
  AOI211_X1 g690(.A(KEYINPUT51), .B(new_n1109), .C1(new_n1115), .C2(G8), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1110), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1045), .A2(new_n1098), .A3(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1115), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1119));
  OAI21_X1  g694(.A(G8), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n1033), .B2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1005), .A2(new_n1028), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT117), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1108), .B(G286), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1035), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1121), .A2(new_n1129), .A3(new_n1122), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1124), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1022), .A2(G1976), .A3(G288), .ZN(new_n1132));
  OAI211_X1 g707(.A(G8), .B(new_n1008), .C1(new_n1132), .C2(new_n1009), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1028), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(new_n1005), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1118), .A2(new_n1131), .A3(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1035), .A2(G171), .A3(new_n986), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1108), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1113), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT51), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1116), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1141), .A2(new_n1142), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1138), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1146), .A2(new_n1144), .A3(new_n1110), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n970), .B1(new_n1137), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n961), .A2(new_n962), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT46), .ZN(new_n1151));
  INV_X1    g726(.A(new_n964), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n961), .B1(new_n792), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT47), .Z(new_n1155));
  NAND2_X1  g730(.A1(new_n963), .A2(new_n964), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n965), .B(KEYINPUT127), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1156), .A2(new_n1157), .B1(G2067), .B2(new_n810), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n961), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n961), .A2(new_n968), .A3(new_n592), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT48), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n961), .A2(new_n967), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1159), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1155), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1149), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g742(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n864), .A2(new_n657), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g744(.A(new_n951), .ZN(new_n1171));
  NOR2_X1   g745(.A1(new_n1170), .A2(new_n1171), .ZN(G308));
  OR2_X1    g746(.A1(new_n1170), .A2(new_n1171), .ZN(G225));
endmodule


