//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT21), .ZN(new_n209));
  NAND2_X1  g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  INV_X1    g009(.A(G71gat), .ZN(new_n211));
  INV_X1    g010(.A(G78gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G64gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G57gat), .ZN(new_n215));
  INV_X1    g014(.A(G57gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G64gat), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n210), .B(new_n213), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT92), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n214), .B2(G57gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n216), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n215), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n210), .B1(new_n213), .B2(new_n219), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT93), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n226), .B1(new_n224), .B2(new_n225), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n220), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n208), .B1(new_n209), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G183gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n209), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT94), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n235), .B2(new_n236), .ZN(new_n240));
  XNOR2_X1  g039(.A(G127gat), .B(G155gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(G211gat), .ZN(new_n242));
  AND2_X1   g041(.A1(G231gat), .A2(G233gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OR3_X1    g044(.A1(new_n239), .A2(new_n240), .A3(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n239), .B2(new_n240), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G190gat), .B(G218gat), .Z(new_n250));
  INV_X1    g049(.A(KEYINPUT96), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT95), .B(KEYINPUT97), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT90), .B(KEYINPUT17), .Z(new_n256));
  XOR2_X1   g055(.A(G43gat), .B(G50gat), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT87), .ZN(new_n258));
  XNOR2_X1  g057(.A(G43gat), .B(G50gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT87), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n258), .A2(KEYINPUT15), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G29gat), .ZN(new_n263));
  INV_X1    g062(.A(G36gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT14), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT14), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(G29gat), .B2(G36gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT88), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT88), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n270), .B(new_n271), .C1(new_n263), .C2(new_n264), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT15), .A3(new_n261), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT15), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n257), .A2(new_n275), .B1(G29gat), .B2(G36gat), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n274), .A2(new_n267), .A3(new_n265), .A4(new_n276), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n273), .A2(new_n277), .A3(KEYINPUT89), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT89), .B1(new_n273), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n256), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G85gat), .A2(G92gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT7), .ZN(new_n282));
  INV_X1    g081(.A(G85gat), .ZN(new_n283));
  INV_X1    g082(.A(G92gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G99gat), .ZN(new_n286));
  INV_X1    g085(.A(G106gat), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT8), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n282), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G99gat), .B(G106gat), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n292), .A2(new_n285), .A3(new_n282), .A4(new_n288), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n273), .A2(new_n277), .A3(KEYINPUT17), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT41), .ZN(new_n297));
  NAND2_X1  g096(.A1(G232gat), .A2(G233gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n278), .A2(new_n279), .ZN(new_n299));
  OAI221_X1 g098(.A(new_n296), .B1(new_n297), .B2(new_n298), .C1(new_n294), .C2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G134gat), .B(G162gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n297), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n250), .A2(new_n251), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n300), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n300), .B2(new_n305), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n255), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n300), .A2(new_n305), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n303), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n300), .A2(new_n304), .A3(new_n305), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n254), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G8gat), .B(G36gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(new_n284), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT78), .B(G64gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(KEYINPUT37), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT67), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n322), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT24), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT66), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n330), .A2(G169gat), .A3(G176gat), .ZN(new_n331));
  INV_X1    g130(.A(G169gat), .ZN(new_n332));
  INV_X1    g131(.A(G176gat), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT66), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT23), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n332), .A2(new_n333), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337));
  NOR2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n329), .A2(KEYINPUT25), .A3(new_n335), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n326), .ZN(new_n343));
  INV_X1    g142(.A(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n232), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n345), .A3(new_n320), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT65), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n338), .A2(KEYINPUT23), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT65), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n343), .A2(new_n345), .A3(new_n349), .A4(new_n320), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n347), .A2(new_n348), .A3(new_n350), .A4(new_n340), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n324), .B2(new_n328), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT68), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n340), .A4(new_n335), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n342), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT27), .B(G183gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n344), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n338), .A2(KEYINPUT66), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n330), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT26), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT69), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(new_n339), .B2(KEYINPUT26), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n361), .B(new_n327), .C1(new_n368), .C2(new_n336), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n357), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT77), .ZN(new_n371));
  AND2_X1   g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n373), .A3(new_n369), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G211gat), .B(G218gat), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT74), .B(G204gat), .ZN(new_n378));
  INV_X1    g177(.A(G197gat), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382));
  NAND2_X1  g181(.A1(G211gat), .A2(G218gat), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT75), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n377), .B1(new_n385), .B2(KEYINPUT76), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n377), .A2(KEYINPUT76), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n384), .B1(KEYINPUT75), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n372), .A2(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n375), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n357), .A2(new_n373), .A3(new_n369), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n373), .B1(new_n357), .B2(new_n369), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n370), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n372), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n389), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n317), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n319), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n389), .A3(new_n397), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n375), .A2(new_n391), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT37), .B(new_n402), .C1(new_n403), .C2(new_n389), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT38), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(G155gat), .A2(G162gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(G155gat), .A2(G162gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G141gat), .B(G148gat), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT2), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n412), .B1(G155gat), .B2(G162gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n410), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G148gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G141gat), .ZN(new_n416));
  INV_X1    g215(.A(G141gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G148gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G155gat), .B(G162gat), .ZN(new_n420));
  INV_X1    g219(.A(G155gat), .ZN(new_n421));
  INV_X1    g220(.A(G162gat), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT2), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n414), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT3), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(KEYINPUT3), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT79), .ZN(new_n429));
  XNOR2_X1  g228(.A(G127gat), .B(G134gat), .ZN(new_n430));
  INV_X1    g229(.A(G120gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G113gat), .ZN(new_n432));
  INV_X1    g231(.A(G113gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G120gat), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT1), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT70), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI211_X1 g236(.A(KEYINPUT70), .B(KEYINPUT1), .C1(new_n432), .C2(new_n434), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n430), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n430), .B1(new_n435), .B2(new_n436), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n429), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n430), .ZN(new_n443));
  XNOR2_X1  g242(.A(G113gat), .B(G120gat), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT70), .B1(new_n444), .B2(KEYINPUT1), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n432), .A2(new_n434), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT1), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n436), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n443), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n449), .A2(KEYINPUT79), .A3(new_n440), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n426), .B(new_n428), .C1(new_n442), .C2(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n414), .A2(new_n424), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n439), .A2(new_n452), .A3(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT4), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT4), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n439), .A2(new_n452), .A3(new_n455), .A4(new_n441), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G225gat), .A2(G233gat), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n451), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n458), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n439), .A2(new_n429), .A3(new_n441), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT79), .B1(new_n449), .B2(new_n440), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n452), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n453), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT5), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n468));
  XNOR2_X1  g267(.A(G57gat), .B(G85gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G1gat), .B(G29gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  INV_X1    g271(.A(KEYINPUT5), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n459), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n467), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476));
  INV_X1    g275(.A(new_n472), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n459), .B2(new_n465), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n427), .B1(new_n461), .B2(new_n462), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n479), .A2(new_n426), .B1(new_n454), .B2(new_n456), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT5), .B1(new_n480), .B2(new_n458), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n477), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n475), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n472), .A4(new_n474), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n317), .B1(new_n392), .B2(new_n398), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT85), .B1(new_n407), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n375), .A2(new_n389), .A3(new_n391), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n371), .A2(new_n374), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n489), .A2(new_n390), .B1(new_n372), .B2(new_n396), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n488), .B1(new_n490), .B2(new_n389), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(new_n318), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT38), .B1(new_n401), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n317), .B1(new_n491), .B2(new_n318), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(new_n405), .A3(new_n404), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT85), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n487), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT29), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n389), .B1(new_n500), .B2(new_n428), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(G228gat), .B2(G233gat), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n500), .B(new_n425), .C1(new_n384), .C2(new_n376), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n384), .A2(new_n376), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n426), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT83), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT3), .B1(new_n389), .B2(new_n500), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(new_n452), .ZN(new_n509));
  OAI211_X1 g308(.A(G228gat), .B(G233gat), .C1(new_n509), .C2(new_n501), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G22gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(G78gat), .B(G106gat), .ZN(new_n514));
  INV_X1    g313(.A(G50gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n513), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n511), .B(new_n517), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n480), .A2(KEYINPUT39), .A3(new_n458), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n472), .ZN(new_n520));
  OR3_X1    g319(.A1(new_n463), .A2(new_n460), .A3(new_n464), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n521), .B(KEYINPUT39), .C1(new_n458), .C2(new_n480), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT40), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT84), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n475), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(new_n524), .B2(new_n523), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n488), .B(new_n400), .C1(new_n490), .C2(new_n389), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n485), .A2(new_n527), .A3(KEYINPUT30), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n491), .A2(new_n529), .A3(new_n317), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n520), .A2(KEYINPUT40), .A3(new_n522), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n526), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n499), .A2(new_n518), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT71), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n439), .A2(new_n441), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n357), .A2(new_n537), .A3(new_n369), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n357), .B2(new_n369), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G227gat), .A2(G233gat), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n541), .B(KEYINPUT64), .Z(new_n542));
  AOI21_X1  g341(.A(new_n536), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n542), .ZN(new_n544));
  NOR4_X1   g343(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT71), .A4(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT32), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT72), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G15gat), .B(G43gat), .Z(new_n549));
  XNOR2_X1  g348(.A(G71gat), .B(G99gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT33), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n543), .B2(new_n545), .ZN(new_n553));
  OAI211_X1 g352(.A(KEYINPUT72), .B(KEYINPUT32), .C1(new_n543), .C2(new_n545), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n548), .A2(new_n551), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n551), .A2(KEYINPUT33), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n546), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n540), .A2(new_n542), .ZN(new_n559));
  NOR2_X1   g358(.A1(KEYINPUT73), .A2(KEYINPUT34), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(KEYINPUT73), .A2(KEYINPUT34), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n555), .A2(new_n563), .A3(new_n557), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(KEYINPUT36), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n555), .A2(new_n563), .A3(new_n557), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n563), .B1(new_n555), .B2(new_n557), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n518), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n483), .A2(KEYINPUT81), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT81), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n475), .A2(new_n482), .A3(new_n574), .A4(new_n476), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n484), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n531), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n535), .A2(new_n567), .A3(new_n571), .A4(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n518), .B1(new_n569), .B2(new_n570), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT35), .B1(new_n580), .B2(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n483), .A2(new_n484), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT86), .B1(new_n531), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(KEYINPUT35), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n566), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n531), .A2(KEYINPUT86), .A3(new_n582), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n518), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  AOI211_X1 g387(.A(new_n249), .B(new_n313), .C1(new_n579), .C2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n280), .A2(new_n208), .A3(new_n295), .ZN(new_n590));
  INV_X1    g389(.A(new_n208), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n278), .B2(new_n279), .ZN(new_n592));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT91), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n590), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n594), .B(KEYINPUT13), .ZN(new_n599));
  INV_X1    g398(.A(new_n299), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(new_n591), .ZN(new_n601));
  INV_X1    g400(.A(new_n592), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n590), .A2(KEYINPUT18), .A3(new_n592), .A4(new_n595), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n598), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G197gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT11), .B(G169gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT12), .Z(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n598), .A2(new_n603), .A3(new_n610), .A4(new_n604), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n230), .A2(new_n294), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n230), .A2(new_n294), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n230), .A2(new_n294), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT99), .B1(new_n619), .B2(KEYINPUT10), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NOR4_X1   g421(.A1(new_n230), .A2(new_n294), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n618), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G230gat), .ZN(new_n625));
  INV_X1    g424(.A(G233gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n615), .B2(new_n616), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OR3_X1    g432(.A1(new_n629), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n629), .B2(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n614), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n589), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n576), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT100), .B(G1gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1324gat));
  NOR2_X1   g440(.A1(new_n638), .A2(new_n531), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT16), .B(G8gat), .Z(new_n643));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(KEYINPUT42), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n645), .B1(KEYINPUT101), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n642), .A2(new_n644), .A3(KEYINPUT42), .A4(new_n643), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n647), .B(new_n648), .C1(new_n207), .C2(new_n642), .ZN(G1325gat));
  INV_X1    g448(.A(new_n638), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n571), .A2(new_n567), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n650), .A2(G15gat), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(G15gat), .B1(new_n650), .B2(new_n585), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(G1326gat));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n518), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT43), .B(G22gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  AND3_X1   g456(.A1(new_n499), .A2(new_n518), .A3(new_n534), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n571), .A2(new_n567), .A3(new_n578), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n518), .B(new_n586), .C1(new_n569), .C2(new_n570), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n576), .A2(new_n531), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n663), .B(new_n518), .C1(new_n569), .C2(new_n570), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n662), .A2(new_n584), .B1(new_n664), .B2(KEYINPUT35), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n313), .B1(new_n660), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n249), .A2(new_n637), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n576), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n263), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(KEYINPUT103), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n308), .A2(new_n312), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n579), .B2(new_n588), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(KEYINPUT103), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n675), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n666), .A2(new_n674), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n667), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684), .B2(new_n576), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n672), .A2(new_n685), .ZN(G1328gat));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n684), .B2(new_n531), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n667), .B1(new_n680), .B2(new_n681), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(KEYINPUT104), .A3(new_n532), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(G36gat), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n668), .A2(new_n264), .A3(new_n532), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT46), .Z(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(G1329gat));
  INV_X1    g493(.A(new_n651), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT107), .B1(new_n684), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n689), .A2(new_n697), .A3(new_n651), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n696), .A2(G43gat), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(G43gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n668), .A2(new_n700), .A3(new_n585), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT106), .Z(new_n702));
  NAND3_X1  g501(.A1(new_n699), .A2(KEYINPUT47), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n701), .B(KEYINPUT106), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n700), .B1(new_n689), .B2(new_n651), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n707), .ZN(G1330gat));
  AOI21_X1  g507(.A(new_n674), .B1(new_n666), .B2(new_n678), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n677), .A2(new_n675), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n572), .B(new_n683), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT109), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n689), .A2(new_n713), .A3(new_n572), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(G50gat), .A3(new_n714), .ZN(new_n715));
  NOR4_X1   g514(.A1(new_n666), .A2(G50gat), .A3(new_n518), .A4(new_n667), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(KEYINPUT48), .A3(new_n717), .ZN(new_n718));
  AOI211_X1 g517(.A(KEYINPUT108), .B(new_n515), .C1(new_n689), .C2(new_n572), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n711), .B2(G50gat), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n719), .A2(new_n721), .A3(new_n716), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n718), .B1(new_n722), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g522(.A1(new_n589), .A2(new_n636), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n614), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n576), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT110), .B(G57gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1332gat));
  NOR2_X1   g527(.A1(new_n725), .A2(new_n531), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  AND2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(G1333gat));
  OAI21_X1  g532(.A(G71gat), .B1(new_n725), .B2(new_n695), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n724), .A2(new_n211), .A3(new_n614), .A4(new_n585), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1334gat));
  NOR2_X1   g537(.A1(new_n725), .A2(new_n518), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n212), .ZN(G1335gat));
  INV_X1    g539(.A(new_n636), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n612), .A2(new_n613), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n248), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n677), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n677), .A2(KEYINPUT51), .A3(new_n743), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n741), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748), .B2(new_n669), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n682), .A2(new_n636), .A3(new_n743), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n576), .A2(new_n283), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n532), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n746), .A2(new_n747), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n531), .A2(new_n741), .A3(G92gat), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT111), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n753), .A2(G92gat), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n284), .B1(new_n750), .B2(new_n532), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n754), .A2(new_n755), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n758), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n757), .A2(new_n758), .B1(new_n759), .B2(new_n761), .ZN(G1337gat));
  AOI21_X1  g561(.A(G99gat), .B1(new_n748), .B2(new_n585), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n695), .A2(new_n286), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n750), .B2(new_n764), .ZN(G1338gat));
  OR2_X1    g564(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n682), .A2(new_n636), .A3(new_n572), .A4(new_n743), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G106gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n518), .A2(G106gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n748), .A2(new_n770), .ZN(new_n771));
  AND4_X1   g570(.A1(new_n766), .A2(new_n768), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n767), .A2(G106gat), .B1(new_n748), .B2(new_n770), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n766), .B1(new_n773), .B2(new_n769), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n772), .A2(new_n774), .ZN(G1339gat));
  NOR4_X1   g574(.A1(new_n249), .A2(new_n313), .A3(new_n636), .A4(new_n742), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n620), .A2(new_n623), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n778), .A2(new_n779), .A3(new_n627), .A4(new_n618), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT113), .B1(new_n624), .B2(new_n628), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n624), .A2(new_n628), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n780), .B(KEYINPUT54), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n633), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n629), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n783), .A2(new_n786), .A3(KEYINPUT55), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n634), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n590), .A2(new_n592), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT114), .B1(new_n792), .B2(new_n594), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794));
  AOI211_X1 g593(.A(new_n794), .B(new_n595), .C1(new_n590), .C2(new_n592), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n601), .A2(new_n602), .A3(new_n599), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n613), .B1(new_n797), .B2(new_n609), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n676), .A2(new_n791), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n742), .A2(new_n634), .A3(new_n789), .A4(new_n790), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n636), .B(new_n613), .C1(new_n797), .C2(new_n609), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n313), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n249), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n580), .B1(new_n777), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n532), .A2(new_n576), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G113gat), .B1(new_n807), .B2(new_n614), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n669), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n809), .A2(KEYINPUT115), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(KEYINPUT115), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n531), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n742), .A2(new_n433), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n808), .B1(new_n812), .B2(new_n813), .ZN(G1340gat));
  OAI21_X1  g613(.A(G120gat), .B1(new_n807), .B2(new_n741), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n636), .A2(new_n431), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n812), .B2(new_n816), .ZN(G1341gat));
  INV_X1    g616(.A(G127gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n807), .A2(new_n818), .A3(new_n249), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n812), .A2(new_n249), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n818), .ZN(G1342gat));
  OAI21_X1  g620(.A(G134gat), .B1(new_n807), .B2(new_n676), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT116), .Z(new_n823));
  NOR2_X1   g622(.A1(new_n812), .A2(G134gat), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(KEYINPUT56), .A3(new_n313), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n824), .B2(new_n313), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(G1343gat));
  NOR3_X1   g626(.A1(new_n651), .A2(new_n576), .A3(new_n532), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n777), .A2(new_n803), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n830), .A3(new_n572), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n791), .A2(KEYINPUT117), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n789), .A2(new_n833), .A3(new_n634), .A4(new_n790), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n742), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n313), .B1(new_n835), .B2(new_n801), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n249), .B1(new_n836), .B2(new_n799), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n518), .B1(new_n837), .B2(new_n777), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n828), .B(new_n831), .C1(new_n838), .C2(new_n830), .ZN(new_n839));
  OAI21_X1  g638(.A(G141gat), .B1(new_n839), .B2(new_n614), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n829), .A2(new_n572), .A3(new_n828), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n417), .A3(new_n742), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n415), .A3(new_n636), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT118), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n828), .B(KEYINPUT119), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n838), .A2(KEYINPUT57), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n801), .B1(new_n791), .B2(new_n614), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n676), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n791), .A2(new_n798), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n313), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n248), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(KEYINPUT57), .B(new_n572), .C1(new_n854), .C2(new_n776), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n829), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n572), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n636), .B(new_n848), .C1(new_n849), .C2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n847), .B1(new_n860), .B2(G148gat), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n847), .B(G148gat), .C1(new_n839), .C2(new_n741), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n846), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT121), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n866), .B(new_n846), .C1(new_n861), .C2(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1345gat));
  AOI21_X1  g667(.A(G155gat), .B1(new_n841), .B2(new_n248), .ZN(new_n869));
  INV_X1    g668(.A(new_n839), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n249), .A2(new_n421), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(G1346gat));
  AOI21_X1  g671(.A(G162gat), .B1(new_n841), .B2(new_n313), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n676), .A2(new_n422), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n870), .B2(new_n874), .ZN(G1347gat));
  AOI21_X1  g674(.A(new_n572), .B1(new_n777), .B2(new_n803), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n669), .A2(new_n531), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n585), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n332), .A3(new_n742), .ZN(new_n882));
  INV_X1    g681(.A(new_n876), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n878), .B(KEYINPUT122), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n742), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n886), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT123), .B1(new_n886), .B2(G169gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n882), .B1(new_n887), .B2(new_n888), .ZN(G1348gat));
  OAI21_X1  g688(.A(new_n333), .B1(new_n880), .B2(new_n741), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n741), .A2(new_n333), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n892), .A2(new_n893), .B1(new_n885), .B2(new_n894), .ZN(G1349gat));
  NAND3_X1  g694(.A1(new_n881), .A2(new_n248), .A3(new_n358), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n883), .A2(new_n249), .A3(new_n884), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n232), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n881), .A2(new_n344), .A3(new_n313), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n313), .ZN(new_n901));
  XNOR2_X1  g700(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n901), .A2(G190gat), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n901), .B2(G190gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(G1351gat));
  NAND2_X1  g704(.A1(new_n695), .A2(new_n877), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n849), .B2(new_n859), .ZN(new_n908));
  OAI21_X1  g707(.A(G197gat), .B1(new_n908), .B2(new_n614), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n907), .A2(new_n572), .A3(new_n829), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n379), .A3(new_n742), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1352gat));
  INV_X1    g711(.A(G204gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n913), .A3(new_n636), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n915));
  NAND2_X1  g714(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n915), .B(new_n916), .Z(new_n917));
  OAI21_X1  g716(.A(new_n636), .B1(new_n849), .B2(new_n859), .ZN(new_n918));
  OAI21_X1  g717(.A(G204gat), .B1(new_n918), .B2(new_n906), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1353gat));
  INV_X1    g719(.A(G211gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n910), .A2(new_n921), .A3(new_n248), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n908), .A2(new_n249), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n923), .B2(G211gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1354gat));
  OAI21_X1  g725(.A(G218gat), .B1(new_n908), .B2(new_n676), .ZN(new_n927));
  INV_X1    g726(.A(G218gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n928), .A3(new_n313), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n930), .B(new_n931), .ZN(G1355gat));
endmodule


