

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U324 ( .A(n453), .B(KEYINPUT123), .ZN(n454) );
  XOR2_X1 U325 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n292) );
  XOR2_X1 U326 ( .A(n339), .B(n338), .Z(n293) );
  XNOR2_X1 U327 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n392) );
  XNOR2_X1 U328 ( .A(n393), .B(n392), .ZN(n395) );
  XNOR2_X1 U329 ( .A(n377), .B(n292), .ZN(n378) );
  XNOR2_X1 U330 ( .A(n340), .B(n293), .ZN(n341) );
  XNOR2_X1 U331 ( .A(n379), .B(n378), .ZN(n383) );
  XNOR2_X1 U332 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U333 ( .A(KEYINPUT36), .B(n557), .Z(n586) );
  XNOR2_X1 U334 ( .A(n353), .B(n352), .ZN(n557) );
  XNOR2_X1 U335 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n456) );
  XNOR2_X1 U336 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U337 ( .A(G190GAT), .B(G99GAT), .Z(n295) );
  XOR2_X1 U338 ( .A(G15GAT), .B(G127GAT), .Z(n360) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G71GAT), .Z(n374) );
  XNOR2_X1 U340 ( .A(n360), .B(n374), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U342 ( .A(n296), .B(G134GAT), .Z(n303) );
  XOR2_X1 U343 ( .A(KEYINPUT0), .B(KEYINPUT88), .Z(n298) );
  XNOR2_X1 U344 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n423) );
  XOR2_X1 U346 ( .A(n423), .B(KEYINPUT20), .Z(n300) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(n301), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U351 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n305) );
  XNOR2_X1 U352 ( .A(G113GAT), .B(KEYINPUT94), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U354 ( .A(n307), .B(n306), .Z(n315) );
  XOR2_X1 U355 ( .A(KEYINPUT93), .B(KEYINPUT17), .Z(n309) );
  XNOR2_X1 U356 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U358 ( .A(G169GAT), .B(n310), .Z(n401) );
  XOR2_X1 U359 ( .A(G183GAT), .B(KEYINPUT65), .Z(n312) );
  XNOR2_X1 U360 ( .A(KEYINPUT95), .B(G176GAT), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n401), .B(n313), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n530) );
  XOR2_X1 U364 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n317) );
  XNOR2_X1 U365 ( .A(KEYINPUT69), .B(KEYINPUT71), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n330) );
  XOR2_X1 U367 ( .A(G22GAT), .B(G197GAT), .Z(n319) );
  XNOR2_X1 U368 ( .A(G36GAT), .B(G50GAT), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U370 ( .A(G8GAT), .B(G15GAT), .Z(n321) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(G141GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U373 ( .A(n323), .B(n322), .Z(n328) );
  XOR2_X1 U374 ( .A(G113GAT), .B(G1GAT), .Z(n426) );
  XOR2_X1 U375 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n325) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n426), .B(n326), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U381 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n332) );
  XNOR2_X1 U382 ( .A(G43GAT), .B(G29GAT), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U384 ( .A(KEYINPUT72), .B(n333), .ZN(n347) );
  XOR2_X1 U385 ( .A(n334), .B(n347), .Z(n547) );
  INV_X1 U386 ( .A(n547), .ZN(n573) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G85GAT), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n335), .B(KEYINPUT75), .ZN(n386) );
  XOR2_X1 U389 ( .A(G134GAT), .B(KEYINPUT82), .Z(n427) );
  XOR2_X1 U390 ( .A(n386), .B(n427), .Z(n337) );
  NAND2_X1 U391 ( .A1(G232GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U393 ( .A(G50GAT), .B(G162GAT), .Z(n450) );
  XOR2_X1 U394 ( .A(G36GAT), .B(G190GAT), .Z(n405) );
  XNOR2_X1 U395 ( .A(n450), .B(n405), .ZN(n340) );
  XOR2_X1 U396 ( .A(KEYINPUT83), .B(KEYINPUT79), .Z(n339) );
  XNOR2_X1 U397 ( .A(G106GAT), .B(G218GAT), .ZN(n338) );
  XOR2_X1 U398 ( .A(KEYINPUT10), .B(KEYINPUT81), .Z(n344) );
  XNOR2_X1 U399 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n353) );
  INV_X1 U402 ( .A(n347), .ZN(n351) );
  XOR2_X1 U403 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n349) );
  XNOR2_X1 U404 ( .A(KEYINPUT67), .B(KEYINPUT80), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U406 ( .A(n351), .B(n350), .Z(n352) );
  XOR2_X1 U407 ( .A(G57GAT), .B(KEYINPUT13), .Z(n377) );
  XOR2_X1 U408 ( .A(G8GAT), .B(G183GAT), .Z(n400) );
  XOR2_X1 U409 ( .A(n377), .B(n400), .Z(n355) );
  XNOR2_X1 U410 ( .A(G78GAT), .B(G211GAT), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U412 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n357) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U415 ( .A(n359), .B(n358), .Z(n362) );
  XNOR2_X1 U416 ( .A(G22GAT), .B(G155GAT), .ZN(n451) );
  XOR2_X1 U417 ( .A(n360), .B(n451), .Z(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n370) );
  XOR2_X1 U419 ( .A(KEYINPUT12), .B(G64GAT), .Z(n364) );
  XNOR2_X1 U420 ( .A(G1GAT), .B(G71GAT), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U422 ( .A(KEYINPUT15), .B(KEYINPUT84), .Z(n366) );
  XNOR2_X1 U423 ( .A(KEYINPUT14), .B(KEYINPUT87), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U425 ( .A(n368), .B(n367), .Z(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n554) );
  NOR2_X1 U427 ( .A1(n586), .A2(n554), .ZN(n371) );
  XNOR2_X1 U428 ( .A(KEYINPUT45), .B(n371), .ZN(n389) );
  XOR2_X1 U429 ( .A(G64GAT), .B(G92GAT), .Z(n373) );
  XNOR2_X1 U430 ( .A(G176GAT), .B(G204GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n410) );
  XOR2_X1 U432 ( .A(n410), .B(n374), .Z(n376) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n379) );
  XOR2_X1 U435 ( .A(KEYINPUT77), .B(KEYINPUT33), .Z(n381) );
  XNOR2_X1 U436 ( .A(KEYINPUT73), .B(KEYINPUT32), .ZN(n380) );
  XOR2_X1 U437 ( .A(n381), .B(n380), .Z(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n388) );
  XOR2_X1 U439 ( .A(G78GAT), .B(G148GAT), .Z(n385) );
  XNOR2_X1 U440 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n446) );
  XNOR2_X1 U442 ( .A(n446), .B(n386), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n578) );
  NAND2_X1 U444 ( .A1(n389), .A2(n578), .ZN(n390) );
  XOR2_X1 U445 ( .A(KEYINPUT115), .B(n390), .Z(n391) );
  NOR2_X1 U446 ( .A1(n573), .A2(n391), .ZN(n398) );
  XOR2_X1 U447 ( .A(n578), .B(KEYINPUT41), .Z(n549) );
  OR2_X1 U448 ( .A1(n549), .A2(n547), .ZN(n393) );
  INV_X1 U449 ( .A(n554), .ZN(n581) );
  NOR2_X1 U450 ( .A1(n557), .A2(n581), .ZN(n394) );
  AND2_X1 U451 ( .A1(n395), .A2(n394), .ZN(n396) );
  XOR2_X1 U452 ( .A(n396), .B(KEYINPUT47), .Z(n397) );
  NOR2_X1 U453 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U454 ( .A(KEYINPUT48), .B(n399), .ZN(n527) );
  XOR2_X1 U455 ( .A(n400), .B(KEYINPUT99), .Z(n403) );
  XNOR2_X1 U456 ( .A(n401), .B(KEYINPUT100), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U458 ( .A(n405), .B(n404), .Z(n407) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n412) );
  XOR2_X1 U461 ( .A(G211GAT), .B(KEYINPUT21), .Z(n409) );
  XNOR2_X1 U462 ( .A(G197GAT), .B(G218GAT), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n438) );
  XOR2_X1 U464 ( .A(n438), .B(n410), .Z(n411) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n494) );
  NOR2_X1 U466 ( .A1(n527), .A2(n494), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n413), .B(KEYINPUT54), .ZN(n436) );
  XOR2_X1 U468 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n415) );
  XNOR2_X1 U469 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n435) );
  XOR2_X1 U471 ( .A(G148GAT), .B(G155GAT), .Z(n417) );
  XNOR2_X1 U472 ( .A(G127GAT), .B(G162GAT), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U474 ( .A(KEYINPUT1), .B(KEYINPUT98), .Z(n419) );
  XNOR2_X1 U475 ( .A(G120GAT), .B(KEYINPUT6), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U477 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n422), .B(KEYINPUT2), .ZN(n445) );
  XNOR2_X1 U480 ( .A(n423), .B(n445), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n431) );
  XOR2_X1 U482 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U485 ( .A(n431), .B(n430), .Z(n433) );
  XNOR2_X1 U486 ( .A(G29GAT), .B(G85GAT), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n528) );
  NAND2_X1 U489 ( .A1(n436), .A2(n528), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n437), .B(KEYINPUT64), .ZN(n572) );
  XOR2_X1 U491 ( .A(KEYINPUT23), .B(n438), .Z(n440) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U494 ( .A(G204GAT), .B(KEYINPUT22), .Z(n442) );
  XNOR2_X1 U495 ( .A(KEYINPUT96), .B(KEYINPUT24), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U497 ( .A(n444), .B(n443), .Z(n448) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U501 ( .A(n452), .B(n451), .ZN(n467) );
  NOR2_X1 U502 ( .A1(n572), .A2(n467), .ZN(n455) );
  INV_X1 U503 ( .A(KEYINPUT55), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n455), .B(n454), .ZN(n563) );
  NOR2_X1 U505 ( .A1(n530), .A2(n563), .ZN(n569) );
  NAND2_X1 U506 ( .A1(n569), .A2(n557), .ZN(n457) );
  NAND2_X1 U507 ( .A1(n569), .A2(n573), .ZN(n459) );
  XNOR2_X1 U508 ( .A(KEYINPUT124), .B(G169GAT), .ZN(n458) );
  XNOR2_X1 U509 ( .A(n459), .B(n458), .ZN(G1348GAT) );
  NAND2_X1 U510 ( .A1(n573), .A2(n578), .ZN(n460) );
  XNOR2_X1 U511 ( .A(n460), .B(KEYINPUT78), .ZN(n488) );
  NOR2_X1 U512 ( .A1(n557), .A2(n554), .ZN(n461) );
  XNOR2_X1 U513 ( .A(KEYINPUT16), .B(n461), .ZN(n475) );
  XNOR2_X1 U514 ( .A(KEYINPUT27), .B(n494), .ZN(n465) );
  XNOR2_X1 U515 ( .A(KEYINPUT28), .B(n467), .ZN(n523) );
  NOR2_X1 U516 ( .A1(n465), .A2(n523), .ZN(n529) );
  NAND2_X1 U517 ( .A1(n530), .A2(n529), .ZN(n462) );
  INV_X1 U518 ( .A(n528), .ZN(n516) );
  NAND2_X1 U519 ( .A1(n462), .A2(n516), .ZN(n473) );
  XOR2_X1 U520 ( .A(KEYINPUT101), .B(KEYINPUT26), .Z(n464) );
  NAND2_X1 U521 ( .A1(n530), .A2(n467), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(n571) );
  NOR2_X1 U523 ( .A1(n571), .A2(n465), .ZN(n545) );
  NOR2_X1 U524 ( .A1(n530), .A2(n494), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U526 ( .A(n468), .B(KEYINPUT25), .Z(n469) );
  XNOR2_X1 U527 ( .A(KEYINPUT102), .B(n469), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n545), .A2(n470), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n471), .A2(n528), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n485) );
  INV_X1 U531 ( .A(n485), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n504) );
  NOR2_X1 U533 ( .A1(n488), .A2(n504), .ZN(n483) );
  NAND2_X1 U534 ( .A1(n483), .A2(n516), .ZN(n479) );
  XOR2_X1 U535 ( .A(KEYINPUT104), .B(KEYINPUT34), .Z(n477) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(KEYINPUT103), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(G1324GAT) );
  INV_X1 U539 ( .A(n494), .ZN(n518) );
  NAND2_X1 U540 ( .A1(n483), .A2(n518), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n480), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .Z(n482) );
  INV_X1 U543 ( .A(n530), .ZN(n562) );
  NAND2_X1 U544 ( .A1(n483), .A2(n562), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n482), .B(n481), .ZN(G1326GAT) );
  NAND2_X1 U546 ( .A1(n483), .A2(n523), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n484), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U548 ( .A1(n586), .A2(n485), .ZN(n486) );
  NAND2_X1 U549 ( .A1(n486), .A2(n554), .ZN(n487) );
  XOR2_X1 U550 ( .A(KEYINPUT37), .B(n487), .Z(n515) );
  NOR2_X1 U551 ( .A1(n488), .A2(n515), .ZN(n490) );
  XNOR2_X1 U552 ( .A(KEYINPUT105), .B(KEYINPUT38), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(n502) );
  NOR2_X1 U554 ( .A1(n502), .A2(n528), .ZN(n492) );
  XNOR2_X1 U555 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n502), .A2(n494), .ZN(n496) );
  XNOR2_X1 U559 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n499) );
  NOR2_X1 U563 ( .A1(n530), .A2(n502), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  INV_X1 U566 ( .A(n523), .ZN(n501) );
  NOR2_X1 U567 ( .A1(n502), .A2(n501), .ZN(n503) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n506) );
  INV_X1 U570 ( .A(n549), .ZN(n561) );
  NAND2_X1 U571 ( .A1(n547), .A2(n561), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n514), .A2(n504), .ZN(n511) );
  NAND2_X1 U573 ( .A1(n511), .A2(n516), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n507), .Z(G1332GAT) );
  NAND2_X1 U576 ( .A1(n511), .A2(n518), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U578 ( .A(G71GAT), .B(KEYINPUT111), .Z(n510) );
  NAND2_X1 U579 ( .A1(n511), .A2(n562), .ZN(n509) );
  XNOR2_X1 U580 ( .A(n510), .B(n509), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U582 ( .A1(n511), .A2(n523), .ZN(n512) );
  XNOR2_X1 U583 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n515), .A2(n514), .ZN(n524) );
  NAND2_X1 U585 ( .A1(n516), .A2(n524), .ZN(n517) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n518), .A2(n524), .ZN(n519) );
  XNOR2_X1 U588 ( .A(G92GAT), .B(n519), .ZN(G1337GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n521) );
  NAND2_X1 U590 ( .A1(n524), .A2(n562), .ZN(n520) );
  XNOR2_X1 U591 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(n522), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n525), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT117), .Z(n534) );
  NOR2_X1 U597 ( .A1(n528), .A2(n527), .ZN(n546) );
  NAND2_X1 U598 ( .A1(n546), .A2(n529), .ZN(n531) );
  NOR2_X1 U599 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n532), .B(KEYINPUT116), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n542), .A2(n573), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n536) );
  NAND2_X1 U604 ( .A1(n542), .A2(n561), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT118), .Z(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n540) );
  NAND2_X1 U609 ( .A1(n581), .A2(n542), .ZN(n539) );
  XNOR2_X1 U610 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U613 ( .A1(n557), .A2(n542), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n546), .A2(n545), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n547), .A2(n558), .ZN(n548) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n548), .Z(G1344GAT) );
  NOR2_X1 U618 ( .A1(n558), .A2(n549), .ZN(n553) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n551) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U621 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n554), .A2(n558), .ZN(n555) );
  XOR2_X1 U624 ( .A(KEYINPUT122), .B(n555), .Z(n556) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n556), .ZN(G1346GAT) );
  INV_X1 U626 ( .A(n557), .ZN(n559) );
  NOR2_X1 U627 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n566) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n564) );
  OR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n568) );
  XOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT56), .Z(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n581), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n573), .A2(n582), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  INV_X1 U644 ( .A(n582), .ZN(n585) );
  OR2_X1 U645 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

