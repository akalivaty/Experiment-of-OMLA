

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U554 ( .A1(G164), .A2(G1384), .ZN(n721) );
  NOR2_X1 U555 ( .A1(G651), .A2(G543), .ZN(n781) );
  NOR2_X1 U556 ( .A1(G651), .A2(n561), .ZN(n782) );
  INV_X1 U557 ( .A(G651), .ZN(n523) );
  NOR2_X1 U558 ( .A1(G543), .A2(n523), .ZN(n520) );
  XOR2_X1 U559 ( .A(KEYINPUT1), .B(n520), .Z(n786) );
  NAND2_X1 U560 ( .A1(G61), .A2(n786), .ZN(n522) );
  NAND2_X1 U561 ( .A1(G86), .A2(n781), .ZN(n521) );
  NAND2_X1 U562 ( .A1(n522), .A2(n521), .ZN(n527) );
  XOR2_X1 U563 ( .A(G543), .B(KEYINPUT0), .Z(n561) );
  OR2_X1 U564 ( .A1(n523), .A2(n561), .ZN(n524) );
  XOR2_X2 U565 ( .A(KEYINPUT68), .B(n524), .Z(n783) );
  NAND2_X1 U566 ( .A1(G73), .A2(n783), .ZN(n525) );
  XOR2_X1 U567 ( .A(KEYINPUT2), .B(n525), .Z(n526) );
  NOR2_X1 U568 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U569 ( .A(KEYINPUT81), .B(n528), .Z(n530) );
  NAND2_X1 U570 ( .A1(n782), .A2(G48), .ZN(n529) );
  NAND2_X1 U571 ( .A1(n530), .A2(n529), .ZN(G305) );
  NAND2_X1 U572 ( .A1(G64), .A2(n786), .ZN(n532) );
  NAND2_X1 U573 ( .A1(G52), .A2(n782), .ZN(n531) );
  NAND2_X1 U574 ( .A1(n532), .A2(n531), .ZN(n537) );
  NAND2_X1 U575 ( .A1(n781), .A2(G90), .ZN(n534) );
  NAND2_X1 U576 ( .A1(G77), .A2(n783), .ZN(n533) );
  NAND2_X1 U577 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U578 ( .A(KEYINPUT9), .B(n535), .Z(n536) );
  NOR2_X1 U579 ( .A1(n537), .A2(n536), .ZN(G171) );
  NAND2_X1 U580 ( .A1(n781), .A2(G89), .ZN(n538) );
  XNOR2_X1 U581 ( .A(n538), .B(KEYINPUT4), .ZN(n540) );
  NAND2_X1 U582 ( .A1(G76), .A2(n783), .ZN(n539) );
  NAND2_X1 U583 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U584 ( .A(KEYINPUT5), .B(n541), .ZN(n547) );
  NAND2_X1 U585 ( .A1(n786), .A2(G63), .ZN(n542) );
  XOR2_X1 U586 ( .A(KEYINPUT73), .B(n542), .Z(n544) );
  NAND2_X1 U587 ( .A1(n782), .A2(G51), .ZN(n543) );
  NAND2_X1 U588 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U589 ( .A(KEYINPUT6), .B(n545), .Z(n546) );
  NAND2_X1 U590 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U591 ( .A(KEYINPUT7), .B(n548), .ZN(G168) );
  XOR2_X1 U592 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U593 ( .A1(G50), .A2(n782), .ZN(n550) );
  NAND2_X1 U594 ( .A1(G88), .A2(n781), .ZN(n549) );
  NAND2_X1 U595 ( .A1(n550), .A2(n549), .ZN(n555) );
  NAND2_X1 U596 ( .A1(G75), .A2(n783), .ZN(n551) );
  XNOR2_X1 U597 ( .A(n551), .B(KEYINPUT82), .ZN(n553) );
  NAND2_X1 U598 ( .A1(G62), .A2(n786), .ZN(n552) );
  NAND2_X1 U599 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U600 ( .A1(n555), .A2(n554), .ZN(G166) );
  XOR2_X1 U601 ( .A(KEYINPUT88), .B(G166), .Z(G303) );
  NAND2_X1 U602 ( .A1(n782), .A2(G49), .ZN(n556) );
  XOR2_X1 U603 ( .A(KEYINPUT79), .B(n556), .Z(n558) );
  NAND2_X1 U604 ( .A1(G651), .A2(G74), .ZN(n557) );
  NAND2_X1 U605 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U606 ( .A(KEYINPUT80), .B(n559), .ZN(n560) );
  NOR2_X1 U607 ( .A1(n786), .A2(n560), .ZN(n563) );
  NAND2_X1 U608 ( .A1(n561), .A2(G87), .ZN(n562) );
  NAND2_X1 U609 ( .A1(n563), .A2(n562), .ZN(G288) );
  NAND2_X1 U610 ( .A1(G60), .A2(n786), .ZN(n565) );
  NAND2_X1 U611 ( .A1(G47), .A2(n782), .ZN(n564) );
  NAND2_X1 U612 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U613 ( .A1(G72), .A2(n783), .ZN(n566) );
  XNOR2_X1 U614 ( .A(KEYINPUT69), .B(n566), .ZN(n567) );
  NOR2_X1 U615 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U616 ( .A1(n781), .A2(G85), .ZN(n569) );
  NAND2_X1 U617 ( .A1(n570), .A2(n569), .ZN(G290) );
  XNOR2_X1 U618 ( .A(G1981), .B(KEYINPUT102), .ZN(n571) );
  XNOR2_X1 U619 ( .A(n571), .B(G305), .ZN(n970) );
  XNOR2_X1 U620 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n573) );
  NOR2_X1 U621 ( .A1(G2105), .A2(G2104), .ZN(n572) );
  XNOR2_X2 U622 ( .A(n573), .B(n572), .ZN(n874) );
  NAND2_X1 U623 ( .A1(G137), .A2(n874), .ZN(n575) );
  AND2_X1 U624 ( .A1(G2105), .A2(G2104), .ZN(n878) );
  NAND2_X1 U625 ( .A1(G113), .A2(n878), .ZN(n574) );
  AND2_X1 U626 ( .A1(n575), .A2(n574), .ZN(n756) );
  AND2_X1 U627 ( .A1(n756), .A2(G40), .ZN(n583) );
  INV_X1 U628 ( .A(G2105), .ZN(n578) );
  XNOR2_X1 U629 ( .A(G2104), .B(KEYINPUT64), .ZN(n577) );
  NOR2_X4 U630 ( .A1(n578), .A2(n577), .ZN(n879) );
  NAND2_X1 U631 ( .A1(n879), .A2(G125), .ZN(n576) );
  XNOR2_X1 U632 ( .A(n576), .B(KEYINPUT65), .ZN(n581) );
  AND2_X1 U633 ( .A1(n578), .A2(n577), .ZN(n703) );
  NAND2_X1 U634 ( .A1(n703), .A2(G101), .ZN(n579) );
  XNOR2_X1 U635 ( .A(n579), .B(KEYINPUT23), .ZN(n580) );
  NOR2_X1 U636 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U637 ( .A(n582), .B(KEYINPUT66), .ZN(n755) );
  NAND2_X1 U638 ( .A1(n583), .A2(n755), .ZN(n720) );
  XNOR2_X1 U639 ( .A(n720), .B(KEYINPUT95), .ZN(n593) );
  NAND2_X1 U640 ( .A1(n874), .A2(G138), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n703), .A2(G102), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U643 ( .A(KEYINPUT86), .B(n586), .ZN(n590) );
  NAND2_X1 U644 ( .A1(G114), .A2(n878), .ZN(n588) );
  NAND2_X1 U645 ( .A1(G126), .A2(n879), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U647 ( .A1(n590), .A2(n589), .ZN(n592) );
  INV_X1 U648 ( .A(KEYINPUT87), .ZN(n591) );
  XNOR2_X1 U649 ( .A(n592), .B(n591), .ZN(G164) );
  NAND2_X2 U650 ( .A1(n593), .A2(n721), .ZN(n667) );
  NAND2_X1 U651 ( .A1(G8), .A2(n667), .ZN(n693) );
  NOR2_X1 U652 ( .A1(G1966), .A2(n693), .ZN(n660) );
  INV_X2 U653 ( .A(n667), .ZN(n644) );
  NAND2_X1 U654 ( .A1(G1996), .A2(n644), .ZN(n594) );
  XOR2_X1 U655 ( .A(n594), .B(KEYINPUT26), .Z(n608) );
  NAND2_X1 U656 ( .A1(n667), .A2(G1341), .ZN(n595) );
  XNOR2_X1 U657 ( .A(n595), .B(KEYINPUT98), .ZN(n606) );
  NAND2_X1 U658 ( .A1(n786), .A2(G56), .ZN(n596) );
  XNOR2_X1 U659 ( .A(n596), .B(KEYINPUT14), .ZN(n598) );
  NAND2_X1 U660 ( .A1(G43), .A2(n782), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(n605) );
  NAND2_X1 U662 ( .A1(n781), .A2(G81), .ZN(n599) );
  XNOR2_X1 U663 ( .A(n599), .B(KEYINPUT12), .ZN(n601) );
  NAND2_X1 U664 ( .A1(G68), .A2(n783), .ZN(n600) );
  NAND2_X1 U665 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U666 ( .A(KEYINPUT13), .B(n602), .Z(n603) );
  XNOR2_X1 U667 ( .A(KEYINPUT70), .B(n603), .ZN(n604) );
  NOR2_X2 U668 ( .A1(n605), .A2(n604), .ZN(n974) );
  NAND2_X1 U669 ( .A1(n606), .A2(n974), .ZN(n607) );
  NOR2_X1 U670 ( .A1(n608), .A2(n607), .ZN(n622) );
  NAND2_X1 U671 ( .A1(n781), .A2(G92), .ZN(n609) );
  XOR2_X1 U672 ( .A(KEYINPUT71), .B(n609), .Z(n611) );
  NAND2_X1 U673 ( .A1(n786), .A2(G66), .ZN(n610) );
  NAND2_X1 U674 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U675 ( .A(KEYINPUT72), .B(n612), .ZN(n616) );
  NAND2_X1 U676 ( .A1(n782), .A2(G54), .ZN(n614) );
  NAND2_X1 U677 ( .A1(G79), .A2(n783), .ZN(n613) );
  NAND2_X1 U678 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U679 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U680 ( .A(KEYINPUT15), .B(n617), .Z(n982) );
  NAND2_X1 U681 ( .A1(n622), .A2(n982), .ZN(n621) );
  NAND2_X1 U682 ( .A1(G1348), .A2(n667), .ZN(n619) );
  NAND2_X1 U683 ( .A1(G2067), .A2(n644), .ZN(n618) );
  NAND2_X1 U684 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U685 ( .A1(n621), .A2(n620), .ZN(n624) );
  OR2_X1 U686 ( .A1(n622), .A2(n982), .ZN(n623) );
  NAND2_X1 U687 ( .A1(n624), .A2(n623), .ZN(n636) );
  XOR2_X1 U688 ( .A(KEYINPUT27), .B(KEYINPUT97), .Z(n626) );
  NAND2_X1 U689 ( .A1(G2072), .A2(n644), .ZN(n625) );
  XNOR2_X1 U690 ( .A(n626), .B(n625), .ZN(n628) );
  INV_X1 U691 ( .A(G1956), .ZN(n1003) );
  NOR2_X1 U692 ( .A1(n644), .A2(n1003), .ZN(n627) );
  NOR2_X1 U693 ( .A1(n628), .A2(n627), .ZN(n637) );
  NAND2_X1 U694 ( .A1(G65), .A2(n786), .ZN(n630) );
  NAND2_X1 U695 ( .A1(G53), .A2(n782), .ZN(n629) );
  NAND2_X1 U696 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U697 ( .A1(n781), .A2(G91), .ZN(n632) );
  NAND2_X1 U698 ( .A1(G78), .A2(n783), .ZN(n631) );
  NAND2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U700 ( .A1(n634), .A2(n633), .ZN(n981) );
  NAND2_X1 U701 ( .A1(n637), .A2(n981), .ZN(n635) );
  NAND2_X1 U702 ( .A1(n636), .A2(n635), .ZN(n641) );
  NOR2_X1 U703 ( .A1(n637), .A2(n981), .ZN(n638) );
  XNOR2_X1 U704 ( .A(n638), .B(KEYINPUT28), .ZN(n639) );
  INV_X1 U705 ( .A(n639), .ZN(n640) );
  NAND2_X1 U706 ( .A1(n641), .A2(n640), .ZN(n643) );
  INV_X1 U707 ( .A(KEYINPUT29), .ZN(n642) );
  XNOR2_X1 U708 ( .A(n643), .B(n642), .ZN(n648) );
  XNOR2_X1 U709 ( .A(KEYINPUT25), .B(G2078), .ZN(n916) );
  NOR2_X1 U710 ( .A1(n667), .A2(n916), .ZN(n646) );
  INV_X1 U711 ( .A(G1961), .ZN(n1008) );
  NOR2_X1 U712 ( .A1(n644), .A2(n1008), .ZN(n645) );
  NOR2_X1 U713 ( .A1(n646), .A2(n645), .ZN(n652) );
  NAND2_X1 U714 ( .A1(G171), .A2(n652), .ZN(n647) );
  NAND2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n658) );
  NOR2_X1 U716 ( .A1(G2084), .A2(n667), .ZN(n662) );
  NOR2_X1 U717 ( .A1(n660), .A2(n662), .ZN(n649) );
  NAND2_X1 U718 ( .A1(G8), .A2(n649), .ZN(n650) );
  XNOR2_X1 U719 ( .A(KEYINPUT30), .B(n650), .ZN(n651) );
  NOR2_X1 U720 ( .A1(G168), .A2(n651), .ZN(n654) );
  NOR2_X1 U721 ( .A1(G171), .A2(n652), .ZN(n653) );
  NOR2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n656) );
  XNOR2_X1 U723 ( .A(KEYINPUT31), .B(KEYINPUT99), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n666) );
  INV_X1 U726 ( .A(n666), .ZN(n659) );
  XNOR2_X1 U727 ( .A(KEYINPUT100), .B(n661), .ZN(n665) );
  NAND2_X1 U728 ( .A1(G8), .A2(n662), .ZN(n663) );
  XNOR2_X1 U729 ( .A(KEYINPUT96), .B(n663), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n676) );
  NAND2_X1 U731 ( .A1(n666), .A2(G286), .ZN(n672) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n693), .ZN(n669) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n667), .ZN(n668) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U735 ( .A1(G303), .A2(n670), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U737 ( .A1(n673), .A2(G8), .ZN(n674) );
  XNOR2_X1 U738 ( .A(n674), .B(KEYINPUT32), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n691) );
  NOR2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n682) );
  NOR2_X1 U741 ( .A1(G303), .A2(G1971), .ZN(n677) );
  NOR2_X1 U742 ( .A1(n682), .A2(n677), .ZN(n973) );
  NAND2_X1 U743 ( .A1(n691), .A2(n973), .ZN(n678) );
  NAND2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n972) );
  NAND2_X1 U745 ( .A1(n678), .A2(n972), .ZN(n679) );
  NOR2_X1 U746 ( .A1(n679), .A2(n693), .ZN(n680) );
  NOR2_X1 U747 ( .A1(KEYINPUT33), .A2(n680), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n970), .A2(n681), .ZN(n686) );
  NAND2_X1 U749 ( .A1(KEYINPUT33), .A2(n682), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n693), .A2(n683), .ZN(n684) );
  XNOR2_X1 U751 ( .A(n684), .B(KEYINPUT101), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n698) );
  NOR2_X1 U753 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XOR2_X1 U754 ( .A(n687), .B(KEYINPUT24), .Z(n688) );
  OR2_X1 U755 ( .A1(n693), .A2(n688), .ZN(n696) );
  NOR2_X1 U756 ( .A1(G303), .A2(G2090), .ZN(n689) );
  XOR2_X1 U757 ( .A(KEYINPUT103), .B(n689), .Z(n690) );
  NAND2_X1 U758 ( .A1(G8), .A2(n690), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n734) );
  NAND2_X1 U763 ( .A1(n878), .A2(G107), .ZN(n699) );
  XOR2_X1 U764 ( .A(KEYINPUT89), .B(n699), .Z(n701) );
  NAND2_X1 U765 ( .A1(n879), .A2(G119), .ZN(n700) );
  NAND2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U767 ( .A(KEYINPUT90), .B(n702), .ZN(n706) );
  BUF_X1 U768 ( .A(n703), .Z(n875) );
  NAND2_X1 U769 ( .A1(G95), .A2(n875), .ZN(n704) );
  XNOR2_X1 U770 ( .A(KEYINPUT91), .B(n704), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n874), .A2(G131), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n886) );
  AND2_X1 U774 ( .A1(n886), .A2(G1991), .ZN(n719) );
  NAND2_X1 U775 ( .A1(G105), .A2(n875), .ZN(n709) );
  XNOR2_X1 U776 ( .A(n709), .B(KEYINPUT38), .ZN(n717) );
  NAND2_X1 U777 ( .A1(G129), .A2(n879), .ZN(n710) );
  XNOR2_X1 U778 ( .A(n710), .B(KEYINPUT92), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n878), .A2(G117), .ZN(n711) );
  NAND2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U781 ( .A1(G141), .A2(n874), .ZN(n713) );
  XNOR2_X1 U782 ( .A(KEYINPUT93), .B(n713), .ZN(n714) );
  NOR2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U784 ( .A1(n717), .A2(n716), .ZN(n871) );
  AND2_X1 U785 ( .A1(n871), .A2(G1996), .ZN(n718) );
  NOR2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n941) );
  NOR2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n749) );
  XOR2_X1 U788 ( .A(n749), .B(KEYINPUT94), .Z(n722) );
  NOR2_X1 U789 ( .A1(n941), .A2(n722), .ZN(n740) );
  INV_X1 U790 ( .A(n740), .ZN(n732) );
  XNOR2_X1 U791 ( .A(G2067), .B(KEYINPUT37), .ZN(n746) );
  NAND2_X1 U792 ( .A1(G140), .A2(n874), .ZN(n724) );
  NAND2_X1 U793 ( .A1(G104), .A2(n875), .ZN(n723) );
  NAND2_X1 U794 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U795 ( .A(KEYINPUT34), .B(n725), .ZN(n730) );
  NAND2_X1 U796 ( .A1(G116), .A2(n878), .ZN(n727) );
  NAND2_X1 U797 ( .A1(G128), .A2(n879), .ZN(n726) );
  NAND2_X1 U798 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U799 ( .A(KEYINPUT35), .B(n728), .Z(n729) );
  NOR2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U801 ( .A(KEYINPUT36), .B(n731), .ZN(n889) );
  NOR2_X1 U802 ( .A1(n746), .A2(n889), .ZN(n959) );
  NAND2_X1 U803 ( .A1(n749), .A2(n959), .ZN(n744) );
  NAND2_X1 U804 ( .A1(n732), .A2(n744), .ZN(n733) );
  NOR2_X2 U805 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U806 ( .A(n735), .B(KEYINPUT104), .ZN(n737) );
  XNOR2_X1 U807 ( .A(G1986), .B(G290), .ZN(n986) );
  NAND2_X1 U808 ( .A1(n986), .A2(n749), .ZN(n736) );
  NAND2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n752) );
  NOR2_X1 U810 ( .A1(G1996), .A2(n871), .ZN(n945) );
  NOR2_X1 U811 ( .A1(G1986), .A2(G290), .ZN(n738) );
  NOR2_X1 U812 ( .A1(G1991), .A2(n886), .ZN(n943) );
  NOR2_X1 U813 ( .A1(n738), .A2(n943), .ZN(n739) );
  NOR2_X1 U814 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U815 ( .A1(n945), .A2(n741), .ZN(n742) );
  XOR2_X1 U816 ( .A(n742), .B(KEYINPUT105), .Z(n743) );
  XNOR2_X1 U817 ( .A(KEYINPUT39), .B(n743), .ZN(n745) );
  NAND2_X1 U818 ( .A1(n745), .A2(n744), .ZN(n747) );
  NAND2_X1 U819 ( .A1(n746), .A2(n889), .ZN(n956) );
  NAND2_X1 U820 ( .A1(n747), .A2(n956), .ZN(n748) );
  XNOR2_X1 U821 ( .A(KEYINPUT106), .B(n748), .ZN(n750) );
  NAND2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U823 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U824 ( .A(n753), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U825 ( .A1(n756), .A2(n755), .ZN(G160) );
  AND2_X1 U826 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U827 ( .A(G57), .ZN(G237) );
  INV_X1 U828 ( .A(G132), .ZN(G219) );
  INV_X1 U829 ( .A(G82), .ZN(G220) );
  NAND2_X1 U830 ( .A1(G7), .A2(G661), .ZN(n757) );
  XNOR2_X1 U831 ( .A(n757), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U832 ( .A(G223), .ZN(n818) );
  NAND2_X1 U833 ( .A1(n818), .A2(G567), .ZN(n758) );
  XOR2_X1 U834 ( .A(KEYINPUT11), .B(n758), .Z(G234) );
  NAND2_X1 U835 ( .A1(n974), .A2(G860), .ZN(G153) );
  INV_X1 U836 ( .A(G171), .ZN(G301) );
  NAND2_X1 U837 ( .A1(G868), .A2(G301), .ZN(n760) );
  INV_X1 U838 ( .A(n982), .ZN(n766) );
  INV_X1 U839 ( .A(G868), .ZN(n801) );
  NAND2_X1 U840 ( .A1(n766), .A2(n801), .ZN(n759) );
  NAND2_X1 U841 ( .A1(n760), .A2(n759), .ZN(G284) );
  INV_X1 U842 ( .A(n981), .ZN(G299) );
  NOR2_X1 U843 ( .A1(G286), .A2(n801), .ZN(n762) );
  NOR2_X1 U844 ( .A1(G868), .A2(G299), .ZN(n761) );
  NOR2_X1 U845 ( .A1(n762), .A2(n761), .ZN(G297) );
  INV_X1 U846 ( .A(G860), .ZN(n824) );
  NAND2_X1 U847 ( .A1(n824), .A2(G559), .ZN(n763) );
  NAND2_X1 U848 ( .A1(n763), .A2(n982), .ZN(n764) );
  XNOR2_X1 U849 ( .A(n764), .B(KEYINPUT74), .ZN(n765) );
  XNOR2_X1 U850 ( .A(KEYINPUT16), .B(n765), .ZN(G148) );
  NOR2_X1 U851 ( .A1(n766), .A2(n801), .ZN(n767) );
  XNOR2_X1 U852 ( .A(n767), .B(KEYINPUT75), .ZN(n768) );
  NOR2_X1 U853 ( .A1(G559), .A2(n768), .ZN(n770) );
  AND2_X1 U854 ( .A1(n801), .A2(n974), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n770), .A2(n769), .ZN(G282) );
  NAND2_X1 U856 ( .A1(G135), .A2(n874), .ZN(n772) );
  NAND2_X1 U857 ( .A1(G111), .A2(n878), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n778) );
  NAND2_X1 U859 ( .A1(G123), .A2(n879), .ZN(n773) );
  XNOR2_X1 U860 ( .A(n773), .B(KEYINPUT18), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G99), .A2(n875), .ZN(n774) );
  XNOR2_X1 U862 ( .A(n774), .B(KEYINPUT76), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n939) );
  XNOR2_X1 U865 ( .A(G2096), .B(n939), .ZN(n780) );
  INV_X1 U866 ( .A(G2100), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(G156) );
  XNOR2_X1 U868 ( .A(G305), .B(G288), .ZN(n798) );
  NAND2_X1 U869 ( .A1(G93), .A2(n781), .ZN(n791) );
  NAND2_X1 U870 ( .A1(n782), .A2(G55), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G80), .A2(n783), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U873 ( .A1(G67), .A2(n786), .ZN(n787) );
  XNOR2_X1 U874 ( .A(KEYINPUT77), .B(n787), .ZN(n788) );
  NOR2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U876 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U877 ( .A(n792), .B(KEYINPUT78), .ZN(n825) );
  XOR2_X1 U878 ( .A(n825), .B(KEYINPUT83), .Z(n794) );
  XNOR2_X1 U879 ( .A(n981), .B(KEYINPUT19), .ZN(n793) );
  XNOR2_X1 U880 ( .A(n794), .B(n793), .ZN(n795) );
  XNOR2_X1 U881 ( .A(G166), .B(n795), .ZN(n796) );
  XNOR2_X1 U882 ( .A(n796), .B(G290), .ZN(n797) );
  XNOR2_X1 U883 ( .A(n798), .B(n797), .ZN(n893) );
  NAND2_X1 U884 ( .A1(G559), .A2(n982), .ZN(n799) );
  XNOR2_X1 U885 ( .A(n799), .B(n974), .ZN(n823) );
  XNOR2_X1 U886 ( .A(n893), .B(n823), .ZN(n800) );
  NAND2_X1 U887 ( .A1(n800), .A2(G868), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n801), .A2(n825), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n803), .A2(n802), .ZN(G295) );
  NAND2_X1 U890 ( .A1(G2078), .A2(G2084), .ZN(n805) );
  XOR2_X1 U891 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n804) );
  XNOR2_X1 U892 ( .A(n805), .B(n804), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G2090), .A2(n806), .ZN(n807) );
  XNOR2_X1 U894 ( .A(KEYINPUT21), .B(n807), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n808), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U896 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U897 ( .A1(G220), .A2(G219), .ZN(n809) );
  XNOR2_X1 U898 ( .A(KEYINPUT22), .B(n809), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n810), .A2(G96), .ZN(n811) );
  NOR2_X1 U900 ( .A1(n811), .A2(G218), .ZN(n812) );
  XNOR2_X1 U901 ( .A(n812), .B(KEYINPUT85), .ZN(n828) );
  NAND2_X1 U902 ( .A1(n828), .A2(G2106), .ZN(n816) );
  NAND2_X1 U903 ( .A1(G69), .A2(G120), .ZN(n813) );
  NOR2_X1 U904 ( .A1(G237), .A2(n813), .ZN(n814) );
  NAND2_X1 U905 ( .A1(G108), .A2(n814), .ZN(n827) );
  NAND2_X1 U906 ( .A1(n827), .A2(G567), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n830) );
  NAND2_X1 U908 ( .A1(G483), .A2(G661), .ZN(n817) );
  NOR2_X1 U909 ( .A1(n830), .A2(n817), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n821), .A2(G36), .ZN(G176) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n818), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U913 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n820) );
  XNOR2_X1 U915 ( .A(KEYINPUT108), .B(n820), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(G188) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n826), .B(n825), .ZN(G145) );
  INV_X1 U920 ( .A(G120), .ZN(G236) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  INV_X1 U922 ( .A(G69), .ZN(G235) );
  NOR2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U924 ( .A(n829), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U925 ( .A(G261), .ZN(G325) );
  INV_X1 U926 ( .A(n830), .ZN(G319) );
  XOR2_X1 U927 ( .A(G2096), .B(KEYINPUT43), .Z(n832) );
  XNOR2_X1 U928 ( .A(G2090), .B(G2678), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U930 ( .A(n833), .B(KEYINPUT110), .Z(n835) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2072), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U933 ( .A(KEYINPUT42), .B(G2100), .Z(n837) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2084), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(G227) );
  XOR2_X1 U937 ( .A(G1976), .B(G1971), .Z(n841) );
  XNOR2_X1 U938 ( .A(G1986), .B(G1961), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U940 ( .A(n842), .B(G2474), .Z(n844) );
  XNOR2_X1 U941 ( .A(G1966), .B(G1981), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U943 ( .A(KEYINPUT41), .B(G1956), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U947 ( .A1(n879), .A2(G124), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U949 ( .A1(G136), .A2(n874), .ZN(n850) );
  NAND2_X1 U950 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(KEYINPUT111), .B(n852), .Z(n858) );
  NAND2_X1 U952 ( .A1(n878), .A2(G112), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n853), .B(KEYINPUT112), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G100), .A2(n875), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U956 ( .A(KEYINPUT113), .B(n856), .Z(n857) );
  NOR2_X1 U957 ( .A1(n858), .A2(n857), .ZN(G162) );
  XOR2_X1 U958 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n860) );
  XNOR2_X1 U959 ( .A(n939), .B(KEYINPUT48), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n870) );
  NAND2_X1 U961 ( .A1(G142), .A2(n874), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G106), .A2(n875), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n863), .B(KEYINPUT45), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G118), .A2(n878), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n868) );
  NAND2_X1 U967 ( .A1(n879), .A2(G130), .ZN(n866) );
  XOR2_X1 U968 ( .A(KEYINPUT114), .B(n866), .Z(n867) );
  NOR2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(n870), .B(n869), .Z(n873) );
  XOR2_X1 U971 ( .A(n871), .B(G162), .Z(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n885) );
  NAND2_X1 U973 ( .A1(G139), .A2(n874), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G103), .A2(n875), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n884) );
  NAND2_X1 U976 ( .A1(G115), .A2(n878), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G127), .A2(n879), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n950) );
  XOR2_X1 U981 ( .A(n885), .B(n950), .Z(n888) );
  XOR2_X1 U982 ( .A(G160), .B(n886), .Z(n887) );
  XNOR2_X1 U983 ( .A(n888), .B(n887), .ZN(n891) );
  XNOR2_X1 U984 ( .A(n889), .B(G164), .ZN(n890) );
  XNOR2_X1 U985 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U986 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U987 ( .A(n893), .B(KEYINPUT116), .ZN(n895) );
  XNOR2_X1 U988 ( .A(n974), .B(G286), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U990 ( .A(n982), .B(G171), .Z(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G397) );
  XOR2_X1 U993 ( .A(G2454), .B(G2435), .Z(n900) );
  XNOR2_X1 U994 ( .A(G2438), .B(G2427), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n907) );
  XOR2_X1 U996 ( .A(KEYINPUT107), .B(G2446), .Z(n902) );
  XNOR2_X1 U997 ( .A(G2443), .B(G2430), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U999 ( .A(n903), .B(G2451), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G1348), .B(G1341), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1003 ( .A1(n908), .A2(G14), .ZN(n915) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n915), .ZN(n912) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n909) );
  XOR2_X1 U1006 ( .A(KEYINPUT49), .B(n909), .Z(n910) );
  XNOR2_X1 U1007 ( .A(n910), .B(KEYINPUT117), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(n915), .ZN(G401) );
  XNOR2_X1 U1014 ( .A(G27), .B(n916), .ZN(n927) );
  XNOR2_X1 U1015 ( .A(KEYINPUT121), .B(G2072), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n917), .B(G33), .ZN(n922) );
  XOR2_X1 U1017 ( .A(G25), .B(G1991), .Z(n918) );
  NAND2_X1 U1018 ( .A1(n918), .A2(G28), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(G26), .B(G2067), .ZN(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(G32), .B(G1996), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(KEYINPUT122), .B(n923), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n928), .B(KEYINPUT53), .ZN(n931) );
  XOR2_X1 U1027 ( .A(G2084), .B(G34), .Z(n929) );
  XNOR2_X1 U1028 ( .A(KEYINPUT54), .B(n929), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(G35), .B(G2090), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(KEYINPUT55), .B(n934), .ZN(n936) );
  INV_X1 U1033 ( .A(G29), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n937), .A2(G11), .ZN(n966) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n961) );
  XOR2_X1 U1037 ( .A(G2084), .B(G160), .Z(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n949) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n944) );
  XNOR2_X1 U1042 ( .A(KEYINPUT118), .B(n944), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1044 ( .A(KEYINPUT51), .B(n947), .Z(n948) );
  NAND2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n955) );
  XOR2_X1 U1046 ( .A(G2072), .B(n950), .Z(n952) );
  XOR2_X1 U1047 ( .A(G164), .B(G2078), .Z(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1049 ( .A(KEYINPUT50), .B(n953), .Z(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n961), .B(n960), .ZN(n962) );
  OR2_X1 U1054 ( .A1(KEYINPUT55), .A2(n962), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n963), .A2(G29), .ZN(n964) );
  XOR2_X1 U1056 ( .A(KEYINPUT120), .B(n964), .Z(n965) );
  NOR2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n1021) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XNOR2_X1 U1059 ( .A(G171), .B(G1961), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(G1971), .A2(G303), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n980) );
  XOR2_X1 U1062 ( .A(G168), .B(G1966), .Z(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1064 ( .A(KEYINPUT57), .B(n971), .Z(n978) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1066 ( .A(n974), .B(G1341), .Z(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n988) );
  XNOR2_X1 U1070 ( .A(n981), .B(G1956), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(G1348), .B(n982), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1075 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1076 ( .A(KEYINPUT123), .B(n991), .ZN(n1019) );
  XOR2_X1 U1077 ( .A(G1986), .B(G24), .Z(n993) );
  XOR2_X1 U1078 ( .A(G1971), .B(G22), .Z(n992) );
  NAND2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1080 ( .A(G23), .B(G1976), .ZN(n994) );
  NOR2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1082 ( .A(KEYINPUT58), .B(n996), .Z(n1015) );
  XOR2_X1 U1083 ( .A(KEYINPUT125), .B(G4), .Z(n998) );
  XNOR2_X1 U1084 ( .A(G1348), .B(KEYINPUT59), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(n998), .B(n997), .ZN(n1002) );
  XNOR2_X1 U1086 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G1981), .B(G6), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1006) );
  XOR2_X1 U1090 ( .A(G20), .B(n1003), .Z(n1004) );
  XNOR2_X1 U1091 ( .A(KEYINPUT124), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(KEYINPUT60), .B(n1007), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(n1008), .B(G5), .ZN(n1009) );
  NAND2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(G21), .B(G1966), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1013), .Z(n1014) );
  NOR2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1100 ( .A(KEYINPUT61), .B(n1016), .Z(n1017) );
  NOR2_X1 U1101 ( .A1(G16), .A2(n1017), .ZN(n1018) );
  NOR2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1103 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1104 ( .A(KEYINPUT127), .B(n1022), .ZN(n1023) );
  XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1023), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

