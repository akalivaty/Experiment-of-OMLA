//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  AND2_X1   g003(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n206));
  OAI211_X1 g005(.A(KEYINPUT23), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n207), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT25), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(KEYINPUT24), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n219), .A2(KEYINPUT24), .ZN(new_n221));
  OR2_X1    g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n207), .A2(new_n214), .A3(new_n224), .A4(new_n215), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n217), .A2(new_n218), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n227));
  NOR3_X1   g026(.A1(new_n227), .A2(G169gat), .A3(G176gat), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT67), .B1(new_n204), .B2(new_n208), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT23), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n223), .A2(new_n230), .A3(new_n215), .A4(new_n214), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT25), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT27), .B(G183gat), .ZN(new_n234));
  INV_X1    g033(.A(G190gat), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT28), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n238));
  OAI211_X1 g037(.A(KEYINPUT28), .B(new_n235), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n219), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n204), .A2(new_n208), .A3(KEYINPUT67), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n227), .B1(G169gat), .B2(G176gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT26), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n215), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI211_X1 g045(.A(KEYINPUT68), .B(KEYINPUT26), .C1(new_n242), .C2(new_n243), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n209), .A2(KEYINPUT26), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n241), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n203), .B1(new_n233), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(KEYINPUT74), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n233), .B2(new_n250), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT74), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n249), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n246), .A2(new_n258), .A3(new_n247), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n226), .B(new_n232), .C1(new_n259), .C2(new_n241), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n254), .B1(new_n260), .B2(new_n203), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n253), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G197gat), .B(G204gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT22), .ZN(new_n264));
  INV_X1    g063(.A(G211gat), .ZN(new_n265));
  INV_X1    g064(.A(G218gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G211gat), .B(G218gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT75), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n225), .A2(new_n223), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT25), .B1(new_n216), .B2(KEYINPUT66), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n273), .A2(new_n274), .B1(KEYINPUT25), .B2(new_n231), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n228), .B2(new_n229), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n244), .A2(new_n245), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n278), .A2(new_n215), .A3(new_n249), .A4(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n236), .A2(new_n240), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n219), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT29), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n255), .B(new_n272), .C1(new_n283), .C2(new_n254), .ZN(new_n284));
  INV_X1    g083(.A(new_n270), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n251), .A2(KEYINPUT75), .A3(new_n252), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G8gat), .B(G36gat), .ZN(new_n289));
  INV_X1    g088(.A(G64gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G92gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT76), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n296));
  AOI211_X1 g095(.A(new_n296), .B(new_n293), .C1(new_n271), .C2(new_n287), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n202), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n293), .B1(new_n271), .B2(new_n287), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT30), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n271), .A2(new_n287), .A3(new_n293), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT77), .B(G155gat), .ZN(new_n303));
  INV_X1    g102(.A(G162gat), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT2), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G141gat), .B(G148gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G155gat), .B(G162gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT78), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n306), .A2(KEYINPUT2), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n312), .A2(new_n308), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n305), .A2(KEYINPUT78), .A3(new_n307), .A4(new_n308), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G127gat), .B(G134gat), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G113gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(G120gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT69), .B(G113gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(G120gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n317), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT1), .B1(new_n321), .B2(new_n322), .ZN(new_n325));
  XOR2_X1   g124(.A(G113gat), .B(G120gat), .Z(new_n326));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n324), .A2(new_n325), .B1(new_n328), .B2(new_n316), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n316), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n321), .A2(new_n322), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n327), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n335), .B2(new_n323), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT4), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n332), .A2(KEYINPUT3), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n311), .A2(new_n340), .A3(new_n313), .A4(new_n314), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n315), .A2(new_n329), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n332), .A2(new_n336), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n346), .B(KEYINPUT39), .C1(new_n345), .C2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT82), .B(KEYINPUT39), .Z(new_n351));
  NAND3_X1  g150(.A1(new_n343), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT0), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(G57gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G85gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT81), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n350), .A2(new_n352), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT40), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n350), .A2(new_n362), .A3(KEYINPUT40), .A4(new_n352), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT5), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n338), .A2(new_n344), .A3(new_n342), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n341), .A2(new_n336), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n337), .A2(new_n331), .B1(new_n371), .B2(new_n339), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT5), .A3(new_n344), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n361), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n365), .A2(new_n366), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n302), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT37), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n255), .B(new_n256), .C1(new_n283), .C2(new_n254), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n285), .B1(new_n379), .B2(new_n253), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n377), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n284), .A2(new_n286), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n270), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(new_n285), .A3(new_n253), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(KEYINPUT37), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT38), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n381), .A2(new_n385), .A3(new_n386), .A4(new_n293), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n373), .A3(new_n356), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT6), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n372), .A2(new_n344), .B1(new_n367), .B2(KEYINPUT5), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT5), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n369), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n357), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n374), .A3(new_n389), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n387), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n271), .A2(KEYINPUT37), .A3(new_n287), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n397), .A3(new_n293), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT38), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT83), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n295), .A2(new_n297), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(new_n402), .A3(KEYINPUT38), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n396), .A2(new_n400), .A3(new_n401), .A4(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G78gat), .B(G106gat), .Z(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT31), .B(G50gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n340), .B1(new_n270), .B2(KEYINPUT29), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n332), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n341), .A2(new_n203), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(new_n270), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(G228gat), .B(G233gat), .C1(new_n410), .C2(KEYINPUT79), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G228gat), .ZN(new_n415));
  INV_X1    g214(.A(G233gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n417));
  AOI211_X1 g216(.A(new_n415), .B(new_n416), .C1(new_n409), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n411), .A2(new_n270), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n409), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(G22gat), .B1(new_n414), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n407), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G22gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n412), .A2(new_n413), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n418), .A2(new_n420), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n414), .A2(new_n421), .A3(G22gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n428), .A2(new_n423), .A3(new_n429), .A4(new_n407), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n376), .A2(new_n404), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n260), .A2(new_n329), .ZN(new_n436));
  NAND2_X1  g235(.A1(G227gat), .A2(G233gat), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n275), .A2(new_n336), .A3(new_n282), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n440), .B1(KEYINPUT32), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G15gat), .B(G43gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(G71gat), .ZN(new_n444));
  INV_X1    g243(.A(G99gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n446), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n441), .B1(new_n448), .B2(KEYINPUT71), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(KEYINPUT71), .B2(new_n448), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT32), .A3(new_n440), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n439), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(new_n437), .ZN(new_n455));
  NAND2_X1  g254(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n454), .A2(KEYINPUT72), .A3(KEYINPUT34), .A4(new_n437), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n447), .A2(new_n457), .A3(new_n451), .A4(new_n458), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n463));
  OR2_X1    g262(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT73), .A4(KEYINPUT36), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n394), .A2(new_n388), .A3(new_n389), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n370), .A2(new_n373), .A3(KEYINPUT6), .A4(new_n356), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n298), .A2(new_n470), .A3(new_n300), .A4(new_n301), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n467), .B1(new_n471), .B2(new_n433), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n431), .A2(new_n462), .A3(new_n432), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT35), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n298), .A2(new_n301), .ZN(new_n475));
  INV_X1    g274(.A(new_n473), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT35), .B1(new_n395), .B2(new_n390), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n300), .A4(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n435), .A2(new_n472), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n480));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(G29gat), .A2(G36gat), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n482), .A2(KEYINPUT14), .ZN(new_n483));
  INV_X1    g282(.A(new_n482), .ZN(new_n484));
  INV_X1    g283(.A(G29gat), .ZN(new_n485));
  INV_X1    g284(.A(G36gat), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n483), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT15), .ZN(new_n490));
  AOI211_X1 g289(.A(new_n490), .B(new_n483), .C1(new_n484), .C2(new_n487), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n481), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n493));
  INV_X1    g292(.A(new_n481), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT17), .ZN(new_n497));
  INV_X1    g296(.A(G8gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(G15gat), .B(G22gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT16), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(G1gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(G1gat), .B2(new_n499), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI221_X1 g304(.A(new_n501), .B1(new_n502), .B2(new_n498), .C1(G1gat), .C2(new_n499), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n508), .A3(new_n495), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n497), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n496), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(KEYINPUT85), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n506), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G229gat), .A2(G233gat), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n510), .A2(new_n516), .A3(KEYINPUT18), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n512), .A2(new_n515), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n496), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n520), .A2(new_n516), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n517), .B(KEYINPUT13), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n480), .B(new_n518), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(G197gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT11), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(new_n204), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n527), .B(KEYINPUT12), .Z(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n521), .A2(new_n522), .ZN(new_n530));
  INV_X1    g329(.A(new_n518), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n516), .A3(new_n517), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n535), .B(new_n518), .C1(new_n521), .C2(new_n522), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(new_n523), .A3(new_n528), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(new_n538), .A3(KEYINPUT87), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n479), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT96), .B(KEYINPUT7), .ZN(new_n546));
  INV_X1    g345(.A(G85gat), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n547), .A2(new_n292), .A3(KEYINPUT95), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n546), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT97), .B(G85gat), .Z(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT98), .B(G92gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n550), .A2(new_n551), .B1(KEYINPUT8), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G99gat), .B(G106gat), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n549), .A2(new_n557), .A3(new_n553), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(KEYINPUT99), .A3(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n558), .A2(KEYINPUT99), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n511), .ZN(new_n562));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n563), .B(KEYINPUT93), .Z(new_n564));
  INV_X1    g363(.A(KEYINPUT41), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n497), .A2(new_n509), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n562), .B(new_n566), .C1(new_n567), .C2(new_n561), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n568), .A2(G190gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(G190gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n266), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n569), .A2(G218gat), .A3(new_n570), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n564), .A2(new_n565), .ZN(new_n576));
  XOR2_X1   g375(.A(G134gat), .B(G162gat), .Z(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G183gat), .B(G211gat), .Z(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT20), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT9), .ZN(new_n588));
  INV_X1    g387(.A(G71gat), .ZN(new_n589));
  INV_X1    g388(.A(G78gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G71gat), .B(G78gat), .ZN(new_n592));
  INV_X1    g391(.A(G57gat), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT89), .B1(new_n593), .B2(G64gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT89), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n290), .A3(G57gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n290), .A2(G57gat), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n591), .B(new_n592), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT90), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n592), .B(KEYINPUT88), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n593), .A2(G64gat), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n591), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT92), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n519), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n608), .B1(new_n519), .B2(new_n607), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n587), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n519), .A2(new_n607), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT92), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(KEYINPUT20), .A3(new_n609), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n612), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n615), .B1(new_n612), .B2(new_n618), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n586), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(new_n619), .A3(new_n585), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n578), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n606), .B1(new_n560), .B2(new_n559), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n601), .A2(new_n605), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n558), .B2(new_n556), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n627), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n561), .A2(KEYINPUT10), .A3(new_n606), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n628), .A2(new_n630), .ZN(new_n636));
  INV_X1    g435(.A(new_n634), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n208), .ZN(new_n640));
  INV_X1    g439(.A(G204gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n635), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n635), .A2(KEYINPUT100), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n637), .B1(new_n631), .B2(new_n632), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n638), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n644), .B1(new_n649), .B2(new_n642), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n580), .A2(new_n625), .A3(new_n626), .A4(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n545), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n470), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT101), .B(G1gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1324gat));
  INV_X1    g455(.A(new_n653), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n657), .B(new_n302), .C1(new_n500), .C2(new_n498), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659));
  NOR2_X1   g458(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT102), .ZN(new_n665));
  INV_X1    g464(.A(new_n302), .ZN(new_n666));
  OAI21_X1  g465(.A(G8gat), .B1(new_n653), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n665), .A3(new_n667), .ZN(G1325gat));
  INV_X1    g467(.A(G15gat), .ZN(new_n669));
  INV_X1    g468(.A(new_n467), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n653), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n657), .A2(new_n462), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n669), .B2(new_n672), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n653), .A2(new_n434), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT43), .B(G22gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  NAND2_X1  g475(.A1(new_n435), .A2(new_n472), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n478), .A2(new_n474), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n580), .A2(new_n626), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n650), .ZN(new_n682));
  NOR4_X1   g481(.A1(new_n681), .A2(new_n625), .A3(new_n682), .A4(new_n544), .ZN(new_n683));
  INV_X1    g482(.A(new_n470), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n485), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT45), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n679), .A2(new_n687), .A3(new_n680), .ZN(new_n688));
  INV_X1    g487(.A(new_n680), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT44), .B1(new_n479), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n625), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n691), .A2(new_n692), .A3(new_n650), .A4(new_n539), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n470), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n686), .A2(new_n694), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n683), .A2(new_n486), .A3(new_n302), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT46), .Z(new_n697));
  OAI21_X1  g496(.A(G36gat), .B1(new_n693), .B2(new_n666), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1329gat));
  OAI21_X1  g498(.A(G43gat), .B1(new_n693), .B2(new_n670), .ZN(new_n700));
  INV_X1    g499(.A(G43gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n683), .A2(new_n701), .A3(new_n462), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT47), .Z(G1330gat));
  OR2_X1    g503(.A1(new_n693), .A2(new_n434), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n434), .A2(G50gat), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n705), .A2(G50gat), .B1(new_n683), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g507(.A1(new_n479), .A2(new_n539), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n680), .A2(new_n692), .A3(new_n650), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n470), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(new_n593), .ZN(G1332gat));
  INV_X1    g512(.A(new_n711), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n666), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT104), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n717), .B(new_n718), .Z(G1333gat));
  NAND3_X1  g518(.A1(new_n714), .A2(new_n589), .A3(new_n462), .ZN(new_n720));
  OAI21_X1  g519(.A(G71gat), .B1(new_n711), .B2(new_n670), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g524(.A1(new_n711), .A2(new_n434), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT106), .B(G78gat), .Z(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1335gat));
  INV_X1    g527(.A(new_n550), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n470), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n689), .B1(new_n677), .B2(new_n678), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n625), .A2(new_n539), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT51), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  INV_X1    g534(.A(new_n733), .ZN(new_n736));
  NOR4_X1   g535(.A1(new_n479), .A2(new_n735), .A3(new_n689), .A4(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n731), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n681), .B2(new_n736), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT108), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n738), .A2(new_n740), .A3(KEYINPUT109), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT109), .B1(new_n738), .B2(new_n740), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n682), .B(new_n730), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n733), .A2(new_n682), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n744), .B1(new_n691), .B2(new_n746), .ZN(new_n747));
  AOI211_X1 g546(.A(KEYINPUT107), .B(new_n745), .C1(new_n688), .C2(new_n690), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n684), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n729), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n743), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n743), .A2(KEYINPUT110), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1336gat));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n756));
  INV_X1    g555(.A(new_n738), .ZN(new_n757));
  INV_X1    g556(.A(new_n740), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n666), .A2(G92gat), .A3(new_n650), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n756), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  INV_X1    g562(.A(new_n551), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n687), .B1(new_n679), .B2(new_n680), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n479), .A2(KEYINPUT44), .A3(new_n689), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n746), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n764), .B1(new_n767), .B2(new_n666), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT112), .B(new_n760), .C1(new_n757), .C2(new_n758), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n762), .A2(new_n763), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n302), .B1(new_n747), .B2(new_n748), .ZN(new_n771));
  INV_X1    g570(.A(new_n737), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n739), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n771), .A2(new_n764), .B1(new_n773), .B2(new_n760), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n774), .A2(new_n775), .A3(new_n763), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n760), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n767), .A2(KEYINPUT107), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n691), .A2(new_n744), .A3(new_n746), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n666), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n777), .B1(new_n780), .B2(new_n551), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT111), .B1(new_n781), .B2(KEYINPUT52), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n770), .B1(new_n776), .B2(new_n782), .ZN(G1337gat));
  OAI21_X1  g582(.A(new_n682), .B1(new_n741), .B2(new_n742), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n462), .A2(new_n445), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n670), .B1(new_n778), .B2(new_n779), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n784), .A2(new_n785), .B1(new_n445), .B2(new_n786), .ZN(G1338gat));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n434), .A2(new_n650), .A3(G106gat), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n759), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(G106gat), .ZN(new_n792));
  INV_X1    g591(.A(new_n767), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(new_n433), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n433), .B1(new_n747), .B2(new_n748), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n795), .A2(G106gat), .B1(new_n773), .B2(new_n789), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n791), .A2(new_n794), .B1(new_n796), .B2(new_n788), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  INV_X1    g597(.A(new_n539), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n652), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT113), .B1(new_n651), .B2(new_n539), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n646), .A2(new_n647), .ZN(new_n804));
  AOI211_X1 g603(.A(KEYINPUT100), .B(new_n637), .C1(new_n631), .C2(new_n632), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n631), .A2(new_n637), .A3(new_n632), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n635), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(new_n642), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT55), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n806), .A2(new_n811), .A3(new_n642), .A4(new_n808), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n644), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n520), .A2(new_n516), .A3(new_n522), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n510), .A2(new_n516), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(G229gat), .A3(G233gat), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n520), .A2(KEYINPUT114), .A3(new_n516), .A4(new_n522), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n820), .A2(KEYINPUT115), .A3(new_n527), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT115), .B1(new_n820), .B2(new_n527), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n537), .A2(new_n528), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n813), .A2(new_n680), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n822), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n537), .A2(new_n528), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n820), .A2(KEYINPUT115), .A3(new_n527), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n650), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n813), .B2(new_n539), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n825), .B1(new_n831), .B2(new_n680), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n802), .B1(new_n832), .B2(new_n692), .ZN(new_n833));
  NOR4_X1   g632(.A1(new_n833), .A2(new_n470), .A3(new_n302), .A4(new_n473), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n320), .A3(new_n539), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT116), .B1(new_n833), .B2(new_n433), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837));
  AOI211_X1 g636(.A(new_n644), .B(new_n799), .C1(new_n810), .C2(new_n812), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n689), .B1(new_n838), .B2(new_n830), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n625), .B1(new_n839), .B2(new_n825), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n837), .B(new_n434), .C1(new_n840), .C2(new_n802), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n302), .A2(new_n470), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n836), .A2(new_n841), .A3(new_n462), .A4(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n844), .A2(new_n845), .A3(new_n544), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n835), .B1(new_n846), .B2(new_n318), .ZN(G1340gat));
  INV_X1    g646(.A(G120gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n834), .A2(new_n848), .A3(new_n682), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n844), .A2(new_n845), .A3(new_n650), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n848), .ZN(G1341gat));
  AOI21_X1  g650(.A(G127gat), .B1(new_n834), .B2(new_n625), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n844), .A2(new_n845), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n625), .A2(G127gat), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(G1342gat));
  INV_X1    g654(.A(G134gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n834), .A2(new_n856), .A3(new_n680), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT56), .Z(new_n858));
  NOR3_X1   g657(.A1(new_n844), .A2(new_n845), .A3(new_n689), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n856), .ZN(G1343gat));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n861), .B(new_n433), .C1(new_n840), .C2(new_n802), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n467), .A2(new_n302), .A3(new_n470), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n810), .A2(new_n812), .ZN(new_n864));
  INV_X1    g663(.A(new_n644), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n543), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n649), .A2(new_n642), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n868), .B(new_n824), .C1(new_n869), .C2(new_n644), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT118), .B1(new_n829), .B2(new_n650), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n689), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(KEYINPUT119), .A3(new_n825), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n870), .A2(new_n871), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n866), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n689), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n692), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n802), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n434), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n862), .B(new_n863), .C1(new_n881), .C2(new_n861), .ZN(new_n882));
  OAI21_X1  g681(.A(G141gat), .B1(new_n882), .B2(new_n544), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n833), .B2(new_n470), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT120), .B(new_n684), .C1(new_n840), .C2(new_n802), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n302), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(G141gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n467), .A2(new_n434), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT121), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n887), .A2(new_n888), .A3(new_n543), .A4(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n883), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT119), .B(new_n680), .C1(new_n875), .C2(new_n866), .ZN(new_n894));
  INV_X1    g693(.A(new_n825), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n876), .B2(new_n689), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n896), .B2(KEYINPUT119), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n802), .B1(new_n897), .B2(new_n692), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT57), .B1(new_n898), .B2(new_n434), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n899), .A2(new_n539), .A3(new_n862), .A4(new_n863), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n900), .A2(G141gat), .B1(new_n901), .B2(new_n543), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n893), .B1(new_n902), .B2(new_n903), .ZN(G1344gat));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n905), .B(G148gat), .C1(new_n882), .C2(new_n650), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n625), .B1(new_n873), .B2(new_n825), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n651), .A2(new_n543), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n861), .B(new_n433), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT57), .B1(new_n833), .B2(new_n434), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n909), .A2(new_n910), .A3(new_n682), .A4(new_n863), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G148gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT123), .B1(new_n912), .B2(KEYINPUT59), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  AOI211_X1 g713(.A(new_n914), .B(new_n905), .C1(new_n911), .C2(G148gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n906), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n650), .A2(G148gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n887), .A2(new_n890), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1345gat));
  NOR3_X1   g718(.A1(new_n882), .A2(new_n303), .A3(new_n692), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n887), .A2(new_n625), .A3(new_n890), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n303), .B2(new_n921), .ZN(G1346gat));
  NOR3_X1   g721(.A1(new_n882), .A2(new_n304), .A3(new_n689), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n887), .A2(new_n680), .A3(new_n890), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n304), .B2(new_n924), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n666), .A2(new_n684), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n836), .A2(new_n841), .A3(new_n462), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n544), .ZN(new_n928));
  NOR4_X1   g727(.A1(new_n833), .A2(new_n684), .A3(new_n666), .A4(new_n473), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n204), .A3(new_n539), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1348gat));
  AOI21_X1  g730(.A(G176gat), .B1(new_n929), .B2(new_n682), .ZN(new_n932));
  INV_X1    g731(.A(new_n927), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n650), .A2(new_n206), .A3(new_n205), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G1349gat));
  NOR2_X1   g734(.A1(new_n833), .A2(new_n473), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n936), .A2(new_n625), .A3(new_n234), .A4(new_n926), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT124), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n929), .A2(new_n939), .A3(new_n625), .A4(new_n234), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G183gat), .B1(new_n927), .B2(new_n692), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(KEYINPUT125), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT60), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT60), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n941), .A2(new_n942), .A3(KEYINPUT125), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1350gat));
  OAI21_X1  g746(.A(G190gat), .B1(new_n927), .B2(new_n689), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g749(.A(KEYINPUT126), .B(G190gat), .C1(new_n927), .C2(new_n689), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(KEYINPUT61), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n929), .A2(new_n235), .A3(new_n680), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n948), .A2(new_n949), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(G1351gat));
  NAND2_X1  g755(.A1(new_n926), .A2(new_n670), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n833), .A2(new_n434), .A3(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(G197gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(new_n959), .A3(new_n539), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n909), .A2(new_n910), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n957), .B(KEYINPUT127), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n961), .A2(new_n544), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n963), .B2(new_n959), .ZN(G1352gat));
  NAND3_X1  g763(.A1(new_n958), .A2(new_n641), .A3(new_n682), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT62), .Z(new_n966));
  NOR3_X1   g765(.A1(new_n961), .A2(new_n650), .A3(new_n962), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n641), .B2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n958), .A2(new_n265), .A3(new_n625), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n961), .A2(new_n962), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(new_n625), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  AOI21_X1  g773(.A(G218gat), .B1(new_n958), .B2(new_n680), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n689), .A2(new_n266), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n970), .B2(new_n976), .ZN(G1355gat));
endmodule


