

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(G651), .A2(n575), .ZN(n799) );
  NOR2_X2 U552 ( .A1(G299), .A2(n645), .ZN(n640) );
  AND2_X1 U553 ( .A1(n703), .A2(n702), .ZN(n735) );
  AND2_X1 U554 ( .A1(n679), .A2(n678), .ZN(n680) );
  INV_X4 U555 ( .A(n672), .ZN(n650) );
  BUF_X1 U556 ( .A(n586), .Z(n895) );
  NOR2_X1 U557 ( .A1(n735), .A2(n734), .ZN(n737) );
  XNOR2_X1 U558 ( .A(n680), .B(KEYINPUT32), .ZN(n681) );
  NOR2_X2 U559 ( .A1(G164), .A2(G1384), .ZN(n705) );
  NOR2_X1 U560 ( .A1(n689), .A2(n520), .ZN(n517) );
  OR2_X1 U561 ( .A1(n517), .A2(n518), .ZN(n692) );
  AND2_X1 U562 ( .A1(n519), .A2(KEYINPUT33), .ZN(n518) );
  INV_X1 U563 ( .A(n691), .ZN(n519) );
  OR2_X1 U564 ( .A1(n700), .A2(n691), .ZN(n520) );
  OR2_X1 U565 ( .A1(n1010), .A2(n631), .ZN(n632) );
  OR2_X1 U566 ( .A1(n600), .A2(n599), .ZN(n601) );
  INV_X1 U567 ( .A(KEYINPUT97), .ZN(n683) );
  AND2_X1 U568 ( .A1(n701), .A2(n521), .ZN(n702) );
  INV_X1 U569 ( .A(KEYINPUT17), .ZN(n539) );
  NOR2_X2 U570 ( .A1(G2104), .A2(G2105), .ZN(n540) );
  XOR2_X1 U571 ( .A(KEYINPUT15), .B(n625), .Z(n1010) );
  OR2_X1 U572 ( .A1(n700), .A2(n699), .ZN(n521) );
  INV_X1 U573 ( .A(KEYINPUT27), .ZN(n634) );
  INV_X1 U574 ( .A(KEYINPUT96), .ZN(n664) );
  NOR2_X1 U575 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U576 ( .A1(n799), .A2(G54), .ZN(n621) );
  INV_X1 U577 ( .A(KEYINPUT99), .ZN(n736) );
  XNOR2_X1 U578 ( .A(n532), .B(KEYINPUT6), .ZN(n533) );
  AND2_X2 U579 ( .A1(n543), .A2(G2104), .ZN(n902) );
  NOR2_X1 U580 ( .A1(G543), .A2(n528), .ZN(n529) );
  NOR2_X2 U581 ( .A1(n575), .A2(n528), .ZN(n792) );
  XNOR2_X1 U582 ( .A(n534), .B(n533), .ZN(n535) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n575) );
  NOR2_X2 U585 ( .A1(n614), .A2(n613), .ZN(n1011) );
  XNOR2_X1 U586 ( .A(KEYINPUT72), .B(n538), .ZN(G168) );
  NOR2_X1 U587 ( .A1(G543), .A2(G651), .ZN(n522) );
  XNOR2_X2 U588 ( .A(n522), .B(KEYINPUT64), .ZN(n795) );
  NAND2_X1 U589 ( .A1(G89), .A2(n795), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n523), .B(KEYINPUT4), .ZN(n525) );
  INV_X1 U591 ( .A(G651), .ZN(n528) );
  NAND2_X1 U592 ( .A1(G76), .A2(n792), .ZN(n524) );
  NAND2_X1 U593 ( .A1(n525), .A2(n524), .ZN(n527) );
  XOR2_X1 U594 ( .A(KEYINPUT5), .B(KEYINPUT69), .Z(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(n536) );
  XOR2_X2 U596 ( .A(KEYINPUT1), .B(n529), .Z(n791) );
  NAND2_X1 U597 ( .A1(G63), .A2(n791), .ZN(n531) );
  NAND2_X1 U598 ( .A1(G51), .A2(n799), .ZN(n530) );
  NAND2_X1 U599 ( .A1(n531), .A2(n530), .ZN(n534) );
  XNOR2_X1 U600 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n532) );
  NAND2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT7), .ZN(n538) );
  INV_X1 U603 ( .A(G2105), .ZN(n543) );
  NAND2_X1 U604 ( .A1(G102), .A2(n902), .ZN(n542) );
  XNOR2_X2 U605 ( .A(n540), .B(n539), .ZN(n899) );
  NAND2_X1 U606 ( .A1(G138), .A2(n899), .ZN(n541) );
  AND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G114), .A2(n894), .ZN(n545) );
  NOR2_X1 U609 ( .A1(G2104), .A2(n543), .ZN(n586) );
  NAND2_X1 U610 ( .A1(G126), .A2(n586), .ZN(n544) );
  NAND2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT89), .ZN(n547) );
  AND2_X2 U613 ( .A1(n548), .A2(n547), .ZN(G164) );
  NAND2_X1 U614 ( .A1(G65), .A2(n791), .ZN(n550) );
  NAND2_X1 U615 ( .A1(G91), .A2(n795), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G78), .A2(n792), .ZN(n552) );
  NAND2_X1 U618 ( .A1(G53), .A2(n799), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  OR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(G299) );
  NAND2_X1 U621 ( .A1(G64), .A2(n791), .ZN(n556) );
  NAND2_X1 U622 ( .A1(G52), .A2(n799), .ZN(n555) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G90), .A2(n795), .ZN(n557) );
  XNOR2_X1 U625 ( .A(KEYINPUT65), .B(n557), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n792), .A2(G77), .ZN(n558) );
  XOR2_X1 U627 ( .A(KEYINPUT66), .B(n558), .Z(n559) );
  NOR2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(KEYINPUT9), .ZN(n562) );
  NOR2_X1 U630 ( .A1(n563), .A2(n562), .ZN(G171) );
  INV_X1 U631 ( .A(G171), .ZN(G301) );
  XOR2_X1 U632 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U633 ( .A1(G62), .A2(n791), .ZN(n564) );
  XNOR2_X1 U634 ( .A(n564), .B(KEYINPUT81), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n792), .A2(G75), .ZN(n566) );
  NAND2_X1 U636 ( .A1(G88), .A2(n795), .ZN(n565) );
  NAND2_X1 U637 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U638 ( .A(KEYINPUT82), .B(n567), .Z(n569) );
  NAND2_X1 U639 ( .A1(n799), .A2(G50), .ZN(n568) );
  NAND2_X1 U640 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U641 ( .A1(n571), .A2(n570), .ZN(G166) );
  INV_X1 U642 ( .A(G166), .ZN(G303) );
  NAND2_X1 U643 ( .A1(G49), .A2(n799), .ZN(n573) );
  NAND2_X1 U644 ( .A1(G74), .A2(G651), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U646 ( .A1(n791), .A2(n574), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n575), .A2(G87), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(G288) );
  NAND2_X1 U649 ( .A1(G61), .A2(n791), .ZN(n578) );
  XNOR2_X1 U650 ( .A(n578), .B(KEYINPUT80), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n799), .A2(G48), .ZN(n580) );
  NAND2_X1 U652 ( .A1(G86), .A2(n795), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n792), .A2(G73), .ZN(n581) );
  XOR2_X1 U655 ( .A(KEYINPUT2), .B(n581), .Z(n582) );
  NOR2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(G305) );
  NAND2_X1 U658 ( .A1(G137), .A2(n899), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G125), .A2(n895), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G101), .A2(n902), .ZN(n589) );
  XOR2_X1 U662 ( .A(KEYINPUT23), .B(n589), .Z(n591) );
  NAND2_X1 U663 ( .A1(n894), .A2(G113), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n602) );
  NOR2_X1 U665 ( .A1(n599), .A2(n602), .ZN(G160) );
  NAND2_X1 U666 ( .A1(n792), .A2(G72), .ZN(n593) );
  NAND2_X1 U667 ( .A1(G85), .A2(n795), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G60), .A2(n791), .ZN(n595) );
  NAND2_X1 U670 ( .A1(G47), .A2(n799), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n596) );
  OR2_X1 U672 ( .A1(n597), .A2(n596), .ZN(G290) );
  INV_X1 U673 ( .A(G40), .ZN(n600) );
  NAND2_X2 U674 ( .A1(n705), .A2(n603), .ZN(n672) );
  NAND2_X1 U675 ( .A1(G8), .A2(n672), .ZN(n700) );
  NOR2_X1 U676 ( .A1(G1966), .A2(n700), .ZN(n667) );
  NAND2_X1 U677 ( .A1(n650), .A2(G1996), .ZN(n604) );
  XNOR2_X1 U678 ( .A(n604), .B(KEYINPUT26), .ZN(n615) );
  NAND2_X1 U679 ( .A1(G81), .A2(n795), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n605), .B(KEYINPUT12), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G68), .A2(n792), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT13), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G43), .A2(n799), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n614) );
  XOR2_X1 U686 ( .A(KEYINPUT14), .B(KEYINPUT68), .Z(n612) );
  NAND2_X1 U687 ( .A1(G56), .A2(n791), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n612), .B(n611), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n615), .A2(n1011), .ZN(n618) );
  NAND2_X1 U690 ( .A1(G1341), .A2(n672), .ZN(n616) );
  XNOR2_X1 U691 ( .A(KEYINPUT93), .B(n616), .ZN(n617) );
  NOR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n631) );
  NAND2_X1 U693 ( .A1(G66), .A2(n791), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G92), .A2(n795), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U696 ( .A1(G79), .A2(n792), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n631), .A2(n1010), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n672), .A2(G1348), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(KEYINPUT94), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n650), .A2(G2067), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n644) );
  NAND2_X1 U706 ( .A1(n650), .A2(G2072), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n635), .B(n634), .ZN(n637) );
  NAND2_X1 U708 ( .A1(G1956), .A2(n672), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n645) );
  INV_X1 U710 ( .A(n640), .ZN(n639) );
  INV_X1 U711 ( .A(KEYINPUT95), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n640), .A2(KEYINPUT95), .ZN(n641) );
  NAND2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U716 ( .A1(G299), .A2(n645), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(KEYINPUT28), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n649), .B(KEYINPUT29), .ZN(n654) );
  XOR2_X1 U720 ( .A(G2078), .B(KEYINPUT25), .Z(n973) );
  NOR2_X1 U721 ( .A1(n973), .A2(n672), .ZN(n652) );
  NOR2_X1 U722 ( .A1(n650), .A2(G1961), .ZN(n651) );
  NOR2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n658) );
  NOR2_X1 U724 ( .A1(G301), .A2(n658), .ZN(n653) );
  NOR2_X1 U725 ( .A1(n654), .A2(n653), .ZN(n663) );
  NOR2_X1 U726 ( .A1(G2084), .A2(n672), .ZN(n668) );
  NOR2_X1 U727 ( .A1(n667), .A2(n668), .ZN(n655) );
  NAND2_X1 U728 ( .A1(G8), .A2(n655), .ZN(n656) );
  XNOR2_X1 U729 ( .A(KEYINPUT30), .B(n656), .ZN(n657) );
  NOR2_X1 U730 ( .A1(G168), .A2(n657), .ZN(n660) );
  AND2_X1 U731 ( .A1(G301), .A2(n658), .ZN(n659) );
  NOR2_X1 U732 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U733 ( .A(n661), .B(KEYINPUT31), .ZN(n662) );
  NOR2_X1 U734 ( .A1(n663), .A2(n662), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n665), .B(n664), .ZN(n671) );
  INV_X1 U736 ( .A(n671), .ZN(n666) );
  NOR2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U738 ( .A1(G8), .A2(n668), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n682) );
  NAND2_X1 U740 ( .A1(n671), .A2(G286), .ZN(n679) );
  INV_X1 U741 ( .A(G8), .ZN(n677) );
  NOR2_X1 U742 ( .A1(G1971), .A2(n700), .ZN(n674) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n672), .ZN(n673) );
  NOR2_X1 U744 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U745 ( .A1(n675), .A2(G303), .ZN(n676) );
  OR2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n684) );
  XNOR2_X1 U748 ( .A(n684), .B(n683), .ZN(n693) );
  NOR2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n994) );
  NOR2_X1 U750 ( .A1(G1971), .A2(G303), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n994), .A2(n685), .ZN(n686) );
  NAND2_X1 U752 ( .A1(n693), .A2(n686), .ZN(n687) );
  NAND2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n995) );
  NAND2_X1 U754 ( .A1(n687), .A2(n995), .ZN(n688) );
  XNOR2_X1 U755 ( .A(KEYINPUT98), .B(n688), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n994), .A2(KEYINPUT33), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n690), .A2(n700), .ZN(n691) );
  XOR2_X1 U758 ( .A(G1981), .B(G305), .Z(n1004) );
  NAND2_X1 U759 ( .A1(n692), .A2(n1004), .ZN(n703) );
  NOR2_X1 U760 ( .A1(G2090), .A2(G303), .ZN(n694) );
  NAND2_X1 U761 ( .A1(G8), .A2(n694), .ZN(n695) );
  NAND2_X1 U762 ( .A1(n693), .A2(n695), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n696), .A2(n700), .ZN(n701) );
  NOR2_X1 U764 ( .A1(G1981), .A2(G305), .ZN(n697) );
  XOR2_X1 U765 ( .A(n697), .B(KEYINPUT92), .Z(n698) );
  XNOR2_X1 U766 ( .A(KEYINPUT24), .B(n698), .ZN(n699) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n704) );
  NOR2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n749) );
  NAND2_X1 U769 ( .A1(G104), .A2(n902), .ZN(n707) );
  NAND2_X1 U770 ( .A1(G140), .A2(n899), .ZN(n706) );
  NAND2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n708), .ZN(n713) );
  NAND2_X1 U773 ( .A1(G116), .A2(n894), .ZN(n710) );
  NAND2_X1 U774 ( .A1(G128), .A2(n895), .ZN(n709) );
  NAND2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U776 ( .A(n711), .B(KEYINPUT35), .Z(n712) );
  NOR2_X1 U777 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U778 ( .A(KEYINPUT36), .B(n714), .Z(n715) );
  XOR2_X1 U779 ( .A(KEYINPUT90), .B(n715), .Z(n908) );
  XNOR2_X1 U780 ( .A(KEYINPUT37), .B(G2067), .ZN(n747) );
  NOR2_X1 U781 ( .A1(n908), .A2(n747), .ZN(n940) );
  NAND2_X1 U782 ( .A1(n749), .A2(n940), .ZN(n745) );
  NAND2_X1 U783 ( .A1(G107), .A2(n894), .ZN(n717) );
  NAND2_X1 U784 ( .A1(G95), .A2(n902), .ZN(n716) );
  NAND2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n721) );
  NAND2_X1 U786 ( .A1(G119), .A2(n895), .ZN(n719) );
  NAND2_X1 U787 ( .A1(G131), .A2(n899), .ZN(n718) );
  NAND2_X1 U788 ( .A1(n719), .A2(n718), .ZN(n720) );
  OR2_X1 U789 ( .A1(n721), .A2(n720), .ZN(n889) );
  NAND2_X1 U790 ( .A1(G1991), .A2(n889), .ZN(n722) );
  XNOR2_X1 U791 ( .A(n722), .B(KEYINPUT91), .ZN(n731) );
  NAND2_X1 U792 ( .A1(G117), .A2(n894), .ZN(n724) );
  NAND2_X1 U793 ( .A1(G129), .A2(n895), .ZN(n723) );
  NAND2_X1 U794 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U795 ( .A1(n902), .A2(G105), .ZN(n725) );
  XOR2_X1 U796 ( .A(KEYINPUT38), .B(n725), .Z(n726) );
  NOR2_X1 U797 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n899), .A2(G141), .ZN(n728) );
  NAND2_X1 U799 ( .A1(n729), .A2(n728), .ZN(n885) );
  AND2_X1 U800 ( .A1(G1996), .A2(n885), .ZN(n730) );
  NOR2_X1 U801 ( .A1(n731), .A2(n730), .ZN(n926) );
  INV_X1 U802 ( .A(n749), .ZN(n732) );
  NOR2_X1 U803 ( .A1(n926), .A2(n732), .ZN(n742) );
  INV_X1 U804 ( .A(n742), .ZN(n733) );
  NAND2_X1 U805 ( .A1(n745), .A2(n733), .ZN(n734) );
  XNOR2_X1 U806 ( .A(n737), .B(n736), .ZN(n739) );
  XNOR2_X1 U807 ( .A(G1986), .B(G290), .ZN(n1017) );
  NAND2_X1 U808 ( .A1(n1017), .A2(n749), .ZN(n738) );
  NAND2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n752) );
  NOR2_X1 U810 ( .A1(G1996), .A2(n885), .ZN(n932) );
  NOR2_X1 U811 ( .A1(G1991), .A2(n889), .ZN(n924) );
  NOR2_X1 U812 ( .A1(G1986), .A2(G290), .ZN(n740) );
  NOR2_X1 U813 ( .A1(n924), .A2(n740), .ZN(n741) );
  NOR2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U815 ( .A1(n932), .A2(n743), .ZN(n744) );
  XNOR2_X1 U816 ( .A(n744), .B(KEYINPUT39), .ZN(n746) );
  NAND2_X1 U817 ( .A1(n746), .A2(n745), .ZN(n748) );
  NAND2_X1 U818 ( .A1(n908), .A2(n747), .ZN(n929) );
  NAND2_X1 U819 ( .A1(n748), .A2(n929), .ZN(n750) );
  NAND2_X1 U820 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U821 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U822 ( .A(n753), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U823 ( .A(G2443), .B(G2446), .Z(n755) );
  XNOR2_X1 U824 ( .A(G2427), .B(G2451), .ZN(n754) );
  XNOR2_X1 U825 ( .A(n755), .B(n754), .ZN(n761) );
  XOR2_X1 U826 ( .A(G2430), .B(G2454), .Z(n757) );
  XNOR2_X1 U827 ( .A(G1348), .B(G1341), .ZN(n756) );
  XNOR2_X1 U828 ( .A(n757), .B(n756), .ZN(n759) );
  XOR2_X1 U829 ( .A(G2435), .B(G2438), .Z(n758) );
  XNOR2_X1 U830 ( .A(n759), .B(n758), .ZN(n760) );
  XOR2_X1 U831 ( .A(n761), .B(n760), .Z(n762) );
  AND2_X1 U832 ( .A1(G14), .A2(n762), .ZN(G401) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U834 ( .A(G108), .ZN(G238) );
  INV_X1 U835 ( .A(G132), .ZN(G219) );
  INV_X1 U836 ( .A(G82), .ZN(G220) );
  NAND2_X1 U837 ( .A1(G7), .A2(G661), .ZN(n763) );
  XNOR2_X1 U838 ( .A(n763), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U839 ( .A(G223), .ZN(n833) );
  NAND2_X1 U840 ( .A1(n833), .A2(G567), .ZN(n764) );
  XNOR2_X1 U841 ( .A(n764), .B(KEYINPUT67), .ZN(n765) );
  XNOR2_X1 U842 ( .A(KEYINPUT11), .B(n765), .ZN(G234) );
  NAND2_X1 U843 ( .A1(n1011), .A2(G860), .ZN(G153) );
  NAND2_X1 U844 ( .A1(G868), .A2(G301), .ZN(n767) );
  INV_X1 U845 ( .A(n1010), .ZN(n774) );
  INV_X1 U846 ( .A(G868), .ZN(n814) );
  NAND2_X1 U847 ( .A1(n774), .A2(n814), .ZN(n766) );
  NAND2_X1 U848 ( .A1(n767), .A2(n766), .ZN(G284) );
  NAND2_X1 U849 ( .A1(G868), .A2(G286), .ZN(n769) );
  NAND2_X1 U850 ( .A1(G299), .A2(n814), .ZN(n768) );
  NAND2_X1 U851 ( .A1(n769), .A2(n768), .ZN(G297) );
  INV_X1 U852 ( .A(G559), .ZN(n770) );
  NOR2_X1 U853 ( .A1(G860), .A2(n770), .ZN(n771) );
  XNOR2_X1 U854 ( .A(KEYINPUT73), .B(n771), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n772), .A2(n1010), .ZN(n773) );
  XNOR2_X1 U856 ( .A(n773), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U857 ( .A1(n774), .A2(n814), .ZN(n775) );
  XOR2_X1 U858 ( .A(KEYINPUT74), .B(n775), .Z(n776) );
  NOR2_X1 U859 ( .A1(G559), .A2(n776), .ZN(n777) );
  XOR2_X1 U860 ( .A(KEYINPUT75), .B(n777), .Z(n779) );
  AND2_X1 U861 ( .A1(n814), .A2(n1011), .ZN(n778) );
  NOR2_X1 U862 ( .A1(n779), .A2(n778), .ZN(G282) );
  NAND2_X1 U863 ( .A1(G111), .A2(n894), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G99), .A2(n902), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U866 ( .A(KEYINPUT76), .B(n782), .ZN(n787) );
  NAND2_X1 U867 ( .A1(n895), .A2(G123), .ZN(n783) );
  XNOR2_X1 U868 ( .A(n783), .B(KEYINPUT18), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G135), .A2(n899), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n923) );
  XNOR2_X1 U872 ( .A(n923), .B(G2096), .ZN(n788) );
  XNOR2_X1 U873 ( .A(n788), .B(KEYINPUT77), .ZN(n789) );
  NOR2_X1 U874 ( .A1(G2100), .A2(n789), .ZN(n790) );
  XOR2_X1 U875 ( .A(KEYINPUT78), .B(n790), .Z(G156) );
  NAND2_X1 U876 ( .A1(G67), .A2(n791), .ZN(n794) );
  NAND2_X1 U877 ( .A1(G80), .A2(n792), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U879 ( .A1(G93), .A2(n795), .ZN(n796) );
  XNOR2_X1 U880 ( .A(KEYINPUT79), .B(n796), .ZN(n797) );
  NOR2_X1 U881 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U882 ( .A1(n799), .A2(G55), .ZN(n800) );
  NAND2_X1 U883 ( .A1(n801), .A2(n800), .ZN(n815) );
  NAND2_X1 U884 ( .A1(G559), .A2(n1010), .ZN(n802) );
  XOR2_X1 U885 ( .A(n1011), .B(n802), .Z(n811) );
  NOR2_X1 U886 ( .A1(G860), .A2(n811), .ZN(n803) );
  XOR2_X1 U887 ( .A(n815), .B(n803), .Z(G145) );
  XNOR2_X1 U888 ( .A(G299), .B(G288), .ZN(n809) );
  XNOR2_X1 U889 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n805) );
  XNOR2_X1 U890 ( .A(G290), .B(KEYINPUT19), .ZN(n804) );
  XNOR2_X1 U891 ( .A(n805), .B(n804), .ZN(n806) );
  XOR2_X1 U892 ( .A(n806), .B(G305), .Z(n807) );
  XNOR2_X1 U893 ( .A(n815), .B(n807), .ZN(n808) );
  XNOR2_X1 U894 ( .A(n809), .B(n808), .ZN(n810) );
  XNOR2_X1 U895 ( .A(G166), .B(n810), .ZN(n841) );
  XNOR2_X1 U896 ( .A(n841), .B(n811), .ZN(n812) );
  NAND2_X1 U897 ( .A1(n812), .A2(G868), .ZN(n813) );
  XOR2_X1 U898 ( .A(KEYINPUT85), .B(n813), .Z(n817) );
  NAND2_X1 U899 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U900 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n818) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n818), .Z(n819) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n819), .ZN(n820) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n820), .ZN(n821) );
  NAND2_X1 U905 ( .A1(n821), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(KEYINPUT86), .B(G44), .ZN(n822) );
  XNOR2_X1 U907 ( .A(n822), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n823) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n823), .Z(n824) );
  NOR2_X1 U910 ( .A1(G218), .A2(n824), .ZN(n825) );
  NAND2_X1 U911 ( .A1(G96), .A2(n825), .ZN(n838) );
  NAND2_X1 U912 ( .A1(n838), .A2(G2106), .ZN(n831) );
  NAND2_X1 U913 ( .A1(G120), .A2(G69), .ZN(n826) );
  XOR2_X1 U914 ( .A(KEYINPUT87), .B(n826), .Z(n827) );
  NOR2_X1 U915 ( .A1(G238), .A2(n827), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G57), .A2(n828), .ZN(n837) );
  NAND2_X1 U917 ( .A1(G567), .A2(n837), .ZN(n829) );
  XNOR2_X1 U918 ( .A(KEYINPUT88), .B(n829), .ZN(n830) );
  NAND2_X1 U919 ( .A1(n831), .A2(n830), .ZN(n918) );
  NAND2_X1 U920 ( .A1(G661), .A2(G483), .ZN(n832) );
  NOR2_X1 U921 ( .A1(n918), .A2(n832), .ZN(n836) );
  NAND2_X1 U922 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U925 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n836), .A2(n835), .ZN(G188) );
  XOR2_X1 U928 ( .A(G69), .B(KEYINPUT100), .Z(G235) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U934 ( .A(G286), .B(KEYINPUT111), .ZN(n840) );
  XNOR2_X1 U935 ( .A(G171), .B(n1010), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n843) );
  XOR2_X1 U937 ( .A(n1011), .B(n841), .Z(n842) );
  XNOR2_X1 U938 ( .A(n843), .B(n842), .ZN(n844) );
  NOR2_X1 U939 ( .A1(G37), .A2(n844), .ZN(G397) );
  XNOR2_X1 U940 ( .A(G1956), .B(KEYINPUT41), .ZN(n854) );
  XOR2_X1 U941 ( .A(G1976), .B(G1981), .Z(n846) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1966), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U944 ( .A(G1971), .B(G1961), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U947 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U948 ( .A(KEYINPUT104), .B(G2474), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(G229) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2090), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n855), .B(KEYINPUT103), .ZN(n865) );
  XOR2_X1 U953 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n857) );
  XNOR2_X1 U954 ( .A(KEYINPUT42), .B(G2096), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(G2100), .B(G2084), .Z(n859) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2072), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U960 ( .A(G2678), .B(KEYINPUT43), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(G227) );
  NAND2_X1 U963 ( .A1(G124), .A2(n895), .ZN(n866) );
  XOR2_X1 U964 ( .A(KEYINPUT44), .B(n866), .Z(n867) );
  XNOR2_X1 U965 ( .A(n867), .B(KEYINPUT105), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G136), .A2(n899), .ZN(n868) );
  NAND2_X1 U967 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U968 ( .A(KEYINPUT106), .B(n870), .ZN(n875) );
  NAND2_X1 U969 ( .A1(G112), .A2(n894), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G100), .A2(n902), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(KEYINPUT107), .B(n873), .Z(n874) );
  NOR2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(KEYINPUT108), .B(n876), .ZN(G162) );
  XNOR2_X1 U975 ( .A(G160), .B(G162), .ZN(n888) );
  NAND2_X1 U976 ( .A1(G106), .A2(n902), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G142), .A2(n899), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U979 ( .A(n879), .B(KEYINPUT45), .ZN(n884) );
  NAND2_X1 U980 ( .A1(G118), .A2(n894), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G130), .A2(n895), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U983 ( .A(KEYINPUT109), .B(n882), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n893) );
  XNOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n889), .B(n923), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(n893), .B(n892), .Z(n907) );
  NAND2_X1 U991 ( .A1(G115), .A2(n894), .ZN(n897) );
  NAND2_X1 U992 ( .A1(G127), .A2(n895), .ZN(n896) );
  NAND2_X1 U993 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n898), .B(KEYINPUT47), .ZN(n901) );
  NAND2_X1 U995 ( .A1(G139), .A2(n899), .ZN(n900) );
  NAND2_X1 U996 ( .A1(n901), .A2(n900), .ZN(n905) );
  NAND2_X1 U997 ( .A1(n902), .A2(G103), .ZN(n903) );
  XOR2_X1 U998 ( .A(KEYINPUT110), .B(n903), .Z(n904) );
  NOR2_X1 U999 ( .A1(n905), .A2(n904), .ZN(n919) );
  XNOR2_X1 U1000 ( .A(G164), .B(n919), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n910), .ZN(G395) );
  NOR2_X1 U1004 ( .A1(G401), .A2(n918), .ZN(n915) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G397), .A2(n913), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(n916), .A2(G395), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(n917), .B(KEYINPUT113), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n918), .ZN(G319) );
  INV_X1 U1014 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1015 ( .A(G2072), .B(n919), .Z(n921) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT50), .B(n922), .ZN(n938) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1020 ( .A1(n926), .A2(n925), .ZN(n928) );
  XOR2_X1 U1021 ( .A(G160), .B(G2084), .Z(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n930) );
  NAND2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n936) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(KEYINPUT51), .B(n933), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(KEYINPUT114), .B(n934), .ZN(n935) );
  NOR2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1029 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1030 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n941), .ZN(n943) );
  INV_X1 U1032 ( .A(KEYINPUT55), .ZN(n942) );
  NAND2_X1 U1033 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1034 ( .A1(n944), .A2(G29), .ZN(n1027) );
  XNOR2_X1 U1035 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(n945), .B(KEYINPUT60), .ZN(n955) );
  XNOR2_X1 U1037 ( .A(G1956), .B(G20), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(G6), .B(G1981), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n953) );
  XOR2_X1 U1040 ( .A(G1348), .B(KEYINPUT59), .Z(n948) );
  XNOR2_X1 U1041 ( .A(G4), .B(n948), .ZN(n951) );
  XOR2_X1 U1042 ( .A(G1341), .B(KEYINPUT123), .Z(n949) );
  XNOR2_X1 U1043 ( .A(G19), .B(n949), .ZN(n950) );
  NOR2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(n955), .B(n954), .ZN(n959) );
  XNOR2_X1 U1047 ( .A(G1966), .B(G21), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(G5), .B(G1961), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n967) );
  XNOR2_X1 U1051 ( .A(G1986), .B(G24), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(G23), .B(G1976), .ZN(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1054 ( .A(G1971), .B(KEYINPUT126), .Z(n962) );
  XNOR2_X1 U1055 ( .A(G22), .B(n962), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(KEYINPUT58), .B(n965), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1059 ( .A(KEYINPUT61), .B(n968), .Z(n970) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT122), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n1025) );
  INV_X1 U1062 ( .A(G29), .ZN(n991) );
  XOR2_X1 U1063 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n989) );
  XNOR2_X1 U1064 ( .A(G2090), .B(G35), .ZN(n984) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G26), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G2072), .B(G33), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(G1996), .B(G32), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(G27), .B(n973), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n981) );
  XOR2_X1 U1072 ( .A(G1991), .B(G25), .Z(n978) );
  NAND2_X1 U1073 ( .A1(n978), .A2(G28), .ZN(n979) );
  XOR2_X1 U1074 ( .A(KEYINPUT115), .B(n979), .Z(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT53), .B(n982), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1078 ( .A(G2084), .B(G34), .Z(n985) );
  XNOR2_X1 U1079 ( .A(KEYINPUT54), .B(n985), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(n989), .B(n988), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n992), .A2(G11), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n993), .B(KEYINPUT117), .ZN(n1023) );
  XNOR2_X1 U1085 ( .A(G16), .B(KEYINPUT56), .ZN(n1021) );
  XNOR2_X1 U1086 ( .A(G171), .B(G1961), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(G166), .B(G1971), .ZN(n999) );
  INV_X1 U1088 ( .A(n994), .ZN(n996) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1090 ( .A(KEYINPUT120), .B(n997), .Z(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(n1000), .B(KEYINPUT121), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(KEYINPUT119), .B(KEYINPUT57), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(G1966), .B(KEYINPUT118), .ZN(n1003) );
  XNOR2_X1 U1096 ( .A(n1003), .B(G168), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1098 ( .A(n1007), .B(n1006), .Z(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1019) );
  XNOR2_X1 U1100 ( .A(G1348), .B(n1010), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(n1011), .B(G1341), .Z(n1013) );
  XNOR2_X1 U1102 ( .A(G299), .B(G1956), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

