//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n538, new_n539, new_n540, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n557, new_n558, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n584, new_n585, new_n586, new_n587, new_n590,
    new_n592, new_n593, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1103, new_n1104, new_n1105;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G221), .A3(G220), .A4(G218), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n460), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n460), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n464), .A2(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G112), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n460), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n480));
  AOI211_X1 g055(.A(new_n474), .B(new_n479), .C1(G136), .C2(new_n480), .ZN(G162));
  OAI211_X1 g056(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n482));
  OR2_X1    g057(.A1(G102), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(new_n485), .A3(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n465), .B2(new_n466), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n492), .C1(new_n466), .C2(new_n465), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n491), .B2(new_n493), .ZN(G164));
  XNOR2_X1  g069(.A(KEYINPUT5), .B(G543), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT6), .B(G651), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G88), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G50), .ZN(new_n500));
  OAI22_X1  g075(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n495), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n501), .A2(new_n504), .ZN(G166));
  NAND3_X1  g080(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n506), .B(KEYINPUT7), .ZN(new_n507));
  INV_X1    g082(.A(G51), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n499), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n495), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n496), .A2(G89), .ZN(new_n511));
  NAND2_X1  g086(.A1(G63), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n514));
  OR3_X1    g089(.A1(new_n509), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n509), .B2(new_n513), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(G168));
  NAND2_X1  g092(.A1(new_n495), .A2(G64), .ZN(new_n518));
  NAND2_X1  g093(.A1(G77), .A2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n503), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(KEYINPUT69), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(KEYINPUT69), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n495), .A2(new_n496), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n496), .A2(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(G90), .A2(new_n523), .B1(new_n524), .B2(G52), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(G301));
  INV_X1    g101(.A(G301), .ZN(G171));
  AOI22_X1  g102(.A1(new_n495), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n503), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(G81), .A2(new_n523), .B1(new_n524), .B2(G43), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n529), .A2(new_n530), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(G153));
  NAND4_X1  g111(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND4_X1  g114(.A1(G319), .A2(G483), .A3(G661), .A4(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT71), .ZN(G188));
  NAND3_X1  g116(.A1(new_n496), .A2(G53), .A3(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT9), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT9), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n496), .A2(new_n544), .A3(G53), .A4(G543), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n543), .A2(new_n545), .B1(G91), .B2(new_n523), .ZN(new_n546));
  NAND2_X1  g121(.A1(G78), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n510), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(KEYINPUT72), .B1(new_n549), .B2(G651), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n495), .A2(G65), .ZN(new_n552));
  AOI211_X1 g127(.A(new_n551), .B(new_n503), .C1(new_n552), .C2(new_n547), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n546), .B1(new_n550), .B2(new_n553), .ZN(G299));
  AND2_X1   g129(.A1(new_n515), .A2(new_n516), .ZN(G286));
  INV_X1    g130(.A(G166), .ZN(G303));
  AND2_X1   g131(.A1(new_n523), .A2(G87), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n495), .B2(G74), .ZN(new_n558));
  INV_X1    g133(.A(G49), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n499), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(G288));
  NAND2_X1  g137(.A1(new_n495), .A2(G61), .ZN(new_n563));
  NAND2_X1  g138(.A1(G73), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n503), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(G86), .A2(new_n523), .B1(new_n524), .B2(G48), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(G305));
  AOI22_X1  g144(.A1(G85), .A2(new_n523), .B1(new_n524), .B2(G47), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n495), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n503), .B2(new_n571), .ZN(G290));
  NAND2_X1  g147(.A1(G301), .A2(G868), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n523), .A2(G92), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT10), .Z(new_n575));
  NAND2_X1  g150(.A1(G79), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G66), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n510), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n524), .B2(G54), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n573), .B1(new_n581), .B2(G868), .ZN(G284));
  OAI21_X1  g157(.A(new_n573), .B1(new_n581), .B2(G868), .ZN(G321));
  NAND2_X1  g158(.A1(G286), .A2(G868), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT74), .ZN(new_n585));
  INV_X1    g160(.A(G299), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n584), .B(KEYINPUT74), .C1(G868), .C2(new_n586), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n585), .A2(new_n587), .ZN(G297));
  XNOR2_X1  g163(.A(G297), .B(KEYINPUT75), .ZN(G280));
  INV_X1    g164(.A(G559), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n581), .B1(new_n590), .B2(G860), .ZN(G148));
  NAND2_X1  g166(.A1(new_n581), .A2(new_n590), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G868), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(G868), .B2(new_n535), .ZN(G323));
  XNOR2_X1  g169(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g170(.A1(new_n480), .A2(G135), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT76), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n477), .A2(G123), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT77), .ZN(new_n599));
  OR2_X1    g174(.A1(G99), .A2(G2105), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n600), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n597), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT78), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(G2096), .Z(new_n604));
  NAND2_X1  g179(.A1(new_n461), .A2(new_n468), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT12), .Z(new_n606));
  XOR2_X1   g181(.A(KEYINPUT13), .B(G2100), .Z(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(G156));
  XOR2_X1   g184(.A(G2451), .B(G2454), .Z(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT16), .ZN(new_n611));
  XNOR2_X1  g186(.A(G1341), .B(G1348), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT14), .ZN(new_n614));
  XNOR2_X1  g189(.A(G2427), .B(G2438), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2430), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2435), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n617), .B2(new_n616), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n613), .B(new_n619), .Z(new_n620));
  XNOR2_X1  g195(.A(G2443), .B(G2446), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(new_n623), .A3(G14), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT79), .Z(G401));
  INV_X1    g200(.A(KEYINPUT18), .ZN(new_n626));
  XOR2_X1   g201(.A(G2084), .B(G2090), .Z(new_n627));
  XNOR2_X1  g202(.A(G2067), .B(G2678), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT17), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  XOR2_X1   g208(.A(G2072), .B(G2078), .Z(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n629), .B2(KEYINPUT18), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(G227));
  XOR2_X1   g212(.A(G1971), .B(G1976), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT19), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1956), .B(G2474), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1961), .B(G1966), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NOR3_X1   g218(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n639), .A2(new_n642), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT20), .Z(new_n646));
  AOI211_X1 g221(.A(new_n644), .B(new_n646), .C1(new_n639), .C2(new_n643), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1991), .B(G1996), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1981), .B(G1986), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G229));
  MUX2_X1   g229(.A(G6), .B(G305), .S(G16), .Z(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT32), .B(G1981), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT81), .Z(new_n657));
  XOR2_X1   g232(.A(new_n655), .B(new_n657), .Z(new_n658));
  INV_X1    g233(.A(G16), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G23), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n561), .B2(new_n659), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT82), .Z(new_n662));
  XOR2_X1   g237(.A(KEYINPUT33), .B(G1976), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n662), .A2(new_n664), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(G22), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(G166), .B2(new_n659), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1971), .ZN(new_n669));
  NOR4_X1   g244(.A1(new_n658), .A2(new_n665), .A3(new_n666), .A4(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT34), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n480), .A2(G131), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n477), .A2(G119), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n460), .A2(G107), .ZN(new_n676));
  OAI21_X1  g251(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n674), .B(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  MUX2_X1   g253(.A(G25), .B(new_n678), .S(G29), .Z(new_n679));
  XOR2_X1   g254(.A(KEYINPUT35), .B(G1991), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  MUX2_X1   g256(.A(G24), .B(G290), .S(G16), .Z(new_n682));
  XOR2_X1   g257(.A(KEYINPUT80), .B(G1986), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND4_X1  g259(.A1(new_n672), .A2(new_n673), .A3(new_n681), .A4(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT36), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n659), .A2(G5), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G171), .B2(new_n659), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT91), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1961), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G32), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT87), .Z(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT26), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n480), .A2(G141), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n477), .A2(G129), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT86), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n692), .B1(new_n701), .B2(new_n691), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT27), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1996), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n691), .A2(G27), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G164), .B2(new_n691), .ZN(new_n706));
  INV_X1    g281(.A(G2078), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(KEYINPUT92), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(KEYINPUT92), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n603), .B2(new_n691), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n659), .A2(G21), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G168), .B2(new_n659), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n709), .B(new_n711), .C1(G1966), .C2(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n690), .A2(new_n704), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT31), .B(G11), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT88), .B(G28), .ZN(new_n717));
  AOI21_X1  g292(.A(G29), .B1(new_n717), .B2(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(KEYINPUT89), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(KEYINPUT30), .B2(new_n717), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(KEYINPUT89), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n716), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n723));
  NAND2_X1  g298(.A1(G103), .A2(G2104), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G2105), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n460), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n480), .A2(G139), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n460), .B2(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G33), .B(new_n729), .S(G29), .Z(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G2072), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(KEYINPUT83), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n722), .B(new_n732), .C1(G2072), .C2(new_n730), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n659), .A2(G20), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT23), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n586), .B2(new_n659), .ZN(new_n736));
  INV_X1    g311(.A(G1956), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n731), .A2(KEYINPUT83), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n691), .A2(G26), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT28), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n480), .A2(G140), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n477), .A2(G128), .ZN(new_n743));
  OR2_X1    g318(.A1(G104), .A2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(new_n691), .ZN(new_n748));
  INV_X1    g323(.A(G2067), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n733), .A2(new_n738), .A3(new_n739), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n691), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n691), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT29), .B(G2090), .Z(new_n754));
  XOR2_X1   g329(.A(new_n753), .B(new_n754), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n659), .A2(G4), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n581), .B2(new_n659), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1348), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT84), .B(KEYINPUT24), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n760), .B2(G34), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G34), .B2(new_n760), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n691), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT85), .ZN(new_n764));
  INV_X1    g339(.A(G2084), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n751), .A2(new_n755), .A3(new_n758), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n713), .A2(G1966), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT90), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n659), .A2(G19), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n535), .B2(new_n659), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1341), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(KEYINPUT90), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n767), .A2(new_n770), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n686), .A2(new_n715), .A3(new_n775), .ZN(G311));
  INV_X1    g351(.A(G311), .ZN(G150));
  AOI22_X1  g352(.A1(G93), .A2(new_n523), .B1(new_n524), .B2(G55), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n495), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(new_n503), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT93), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n533), .A2(new_n534), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n535), .A2(new_n781), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT38), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n581), .A2(G559), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n789), .A2(KEYINPUT39), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(KEYINPUT39), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n790), .A2(new_n791), .A3(G860), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n782), .A2(G860), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT37), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n792), .A2(new_n794), .ZN(G145));
  XNOR2_X1  g370(.A(new_n701), .B(new_n729), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n477), .A2(G130), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n460), .A2(G118), .ZN(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G142), .B2(new_n480), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(new_n606), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n796), .B(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(G164), .B(new_n746), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(new_n678), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n603), .B(G160), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G162), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n806), .B(new_n808), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT94), .B(G37), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT95), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g388(.A(G868), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n782), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n784), .A2(new_n785), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(new_n592), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n580), .B(G299), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n580), .B(new_n586), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT41), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n818), .A2(KEYINPUT41), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n819), .B1(new_n824), .B2(new_n817), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT42), .Z(new_n826));
  NAND3_X1  g401(.A1(new_n567), .A2(G166), .A3(new_n568), .ZN(new_n827));
  NAND2_X1  g402(.A1(G305), .A2(G303), .ZN(new_n828));
  XNOR2_X1  g403(.A(G290), .B(new_n561), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(KEYINPUT96), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(KEYINPUT96), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n826), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n815), .B1(new_n833), .B2(new_n814), .ZN(G295));
  OAI21_X1  g409(.A(new_n815), .B1(new_n833), .B2(new_n814), .ZN(G331));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n836));
  NAND2_X1  g411(.A1(G286), .A2(KEYINPUT97), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n838));
  AOI21_X1  g413(.A(G301), .B1(G168), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n839), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n786), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n816), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n836), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT98), .B1(new_n842), .B2(new_n786), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n824), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n843), .A2(new_n844), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n849), .A3(new_n820), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n843), .A2(new_n820), .A3(new_n844), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT99), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n847), .A2(new_n850), .A3(new_n832), .A4(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n832), .B(KEYINPUT100), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n851), .B(new_n849), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(new_n847), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT43), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n832), .B(KEYINPUT100), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n845), .A2(new_n846), .A3(new_n818), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n820), .A2(KEYINPUT101), .A3(new_n821), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n824), .B2(KEYINPUT101), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n848), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n862), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  AND4_X1   g442(.A1(KEYINPUT43), .A2(new_n867), .A3(new_n810), .A4(new_n853), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT44), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n867), .A2(new_n853), .A3(new_n870), .A4(new_n810), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT43), .B1(new_n855), .B2(new_n859), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n871), .A2(new_n872), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n869), .B1(new_n877), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g453(.A(new_n701), .B(G1996), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n746), .B(new_n749), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n678), .B(new_n680), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G1384), .ZN(new_n885));
  INV_X1    g460(.A(new_n493), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n492), .B1(new_n461), .B2(new_n489), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n885), .B1(new_n888), .B2(new_n487), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT45), .ZN(new_n890));
  INV_X1    g465(.A(G40), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n464), .A2(new_n891), .A3(new_n470), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n884), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT126), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n897), .A2(G1986), .A3(G290), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G1996), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT46), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(KEYINPUT46), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n701), .A2(new_n880), .A3(new_n910), .ZN(new_n911));
  OAI22_X1  g486(.A1(new_n908), .A2(new_n909), .B1(new_n897), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT47), .Z(new_n913));
  INV_X1    g488(.A(new_n680), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n678), .A2(new_n914), .ZN(new_n915));
  OAI22_X1  g490(.A1(new_n881), .A2(new_n915), .B1(G2067), .B2(new_n746), .ZN(new_n916));
  AOI211_X1 g491(.A(new_n904), .B(new_n913), .C1(new_n898), .C2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT114), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT50), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(new_n885), .C1(new_n888), .C2(new_n487), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT104), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n491), .A2(new_n493), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n482), .A2(new_n486), .ZN(new_n923));
  AOI21_X1  g498(.A(G1384), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n892), .B1(new_n924), .B2(new_n919), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT112), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n927), .A3(new_n765), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n465), .A2(new_n466), .ZN(new_n929));
  INV_X1    g504(.A(G125), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n463), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(G2105), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n932), .A2(G40), .A3(new_n469), .A4(new_n467), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n889), .B2(new_n890), .ZN(new_n934));
  OAI211_X1 g509(.A(KEYINPUT45), .B(new_n885), .C1(new_n888), .C2(new_n487), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n928), .B1(G1966), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n927), .B1(new_n926), .B2(new_n765), .ZN(new_n938));
  OAI211_X1 g513(.A(G8), .B(G168), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G8), .ZN(new_n940));
  XNOR2_X1  g515(.A(KEYINPUT105), .B(G2090), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n926), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n936), .A2(G1971), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n940), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(G166), .A2(new_n940), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT106), .B(KEYINPUT55), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n949), .B2(KEYINPUT55), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(KEYINPUT113), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n945), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT63), .B1(new_n945), .B2(new_n953), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n939), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT107), .B(G1976), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT52), .B1(G288), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n892), .A2(new_n924), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G8), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(G1976), .B2(new_n561), .ZN(new_n961));
  MUX2_X1   g536(.A(KEYINPUT52), .B(new_n958), .S(new_n961), .Z(new_n962));
  INV_X1    g537(.A(G1981), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n567), .A2(new_n963), .A3(new_n568), .ZN(new_n964));
  INV_X1    g539(.A(new_n568), .ZN(new_n965));
  OAI21_X1  g540(.A(G1981), .B1(new_n965), .B2(new_n565), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT49), .ZN(new_n968));
  OR3_X1    g543(.A1(new_n967), .A2(KEYINPUT109), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT109), .B1(new_n967), .B2(new_n968), .ZN(new_n970));
  INV_X1    g545(.A(new_n960), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT49), .B1(new_n967), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n964), .A2(KEYINPUT108), .A3(new_n966), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT110), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n970), .A2(new_n971), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n976), .A3(new_n980), .A4(new_n969), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n962), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n918), .B1(new_n956), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n954), .A2(new_n955), .ZN(new_n984));
  INV_X1    g559(.A(new_n939), .ZN(new_n985));
  AND4_X1   g560(.A1(new_n918), .A2(new_n984), .A3(new_n985), .A4(new_n982), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n920), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n924), .A2(KEYINPUT111), .A3(new_n919), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n925), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n943), .B1(new_n990), .B2(new_n941), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n948), .B(new_n950), .C1(new_n991), .C2(new_n940), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n945), .A2(new_n951), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n982), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n939), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n983), .A2(new_n986), .B1(new_n996), .B2(KEYINPUT63), .ZN(new_n997));
  OAI21_X1  g572(.A(G8), .B1(new_n937), .B2(new_n938), .ZN(new_n998));
  NOR2_X1   g573(.A1(G168), .A2(new_n940), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT123), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n998), .B(new_n1000), .C1(new_n1001), .C2(KEYINPUT51), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT51), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1003));
  INV_X1    g578(.A(new_n938), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n928), .C1(G1966), .C2(new_n936), .ZN(new_n1005));
  OAI211_X1 g580(.A(G8), .B(new_n1003), .C1(new_n1005), .C2(G286), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n999), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1002), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1009));
  INV_X1    g584(.A(new_n995), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n936), .A2(new_n707), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n936), .A2(KEYINPUT53), .A3(new_n707), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1013), .B(new_n1014), .C1(G1961), .C2(new_n926), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1015), .A2(G171), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT62), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1002), .A2(new_n1006), .A3(new_n1017), .A4(new_n1007), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1009), .A2(new_n1010), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n978), .A2(new_n981), .ZN(new_n1020));
  OR2_X1    g595(.A1(G288), .A2(G1976), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n964), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n993), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1022), .A2(new_n971), .B1(new_n982), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n997), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1015), .B(G301), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(G171), .B2(KEYINPUT124), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1010), .A2(new_n1008), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n926), .A2(G1348), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n959), .A2(G2067), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT118), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT60), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n581), .A2(KEYINPUT121), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n581), .A2(KEYINPUT121), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1041), .B(new_n1042), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n934), .A2(new_n905), .A3(new_n935), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT58), .B(G1341), .Z(new_n1045));
  NAND2_X1  g620(.A1(new_n959), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n783), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT59), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT56), .B(G2072), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n934), .A2(KEYINPUT116), .A3(new_n935), .A4(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n890), .B1(G164), .B2(G1384), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1051), .A2(new_n935), .A3(new_n892), .A4(new_n1049), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n990), .A2(KEYINPUT115), .A3(G1956), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n933), .B1(new_n889), .B2(KEYINPUT50), .ZN(new_n1058));
  NOR4_X1   g633(.A1(G164), .A2(new_n987), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT111), .B1(new_n924), .B2(new_n919), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1057), .B1(new_n1061), .B2(new_n737), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1055), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n546), .B(new_n1065), .C1(new_n550), .C2(new_n553), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT61), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT115), .B1(new_n990), .B2(G1956), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1061), .A2(new_n1057), .A3(new_n737), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1067), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1048), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1073), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT117), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n1073), .C1(new_n1056), .C2(new_n1062), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1077), .A2(new_n1079), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1075), .B(KEYINPUT120), .C1(new_n1080), .C2(KEYINPUT61), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1079), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1078), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1068), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1069), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT120), .B1(new_n1086), .B2(new_n1075), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1043), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1068), .B1(new_n1035), .B2(new_n580), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1084), .B2(new_n1083), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1031), .B1(new_n1093), .B2(KEYINPUT122), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1088), .A2(new_n1095), .A3(new_n1092), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1025), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n884), .ZN(new_n1098));
  XOR2_X1   g673(.A(G290), .B(G1986), .Z(new_n1099));
  AOI21_X1  g674(.A(new_n897), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n917), .B1(new_n1097), .B2(new_n1100), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g676(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1103));
  AND2_X1   g677(.A1(new_n653), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g678(.A1(new_n812), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g679(.A1(new_n877), .A2(new_n1105), .ZN(G308));
  OR2_X1    g680(.A1(new_n877), .A2(new_n1105), .ZN(G225));
endmodule


