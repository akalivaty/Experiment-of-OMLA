//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  XNOR2_X1  g000(.A(KEYINPUT81), .B(G101), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT80), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  AOI22_X1  g004(.A1(new_n188), .A2(new_n189), .B1(new_n190), .B2(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n192), .A2(new_n190), .A3(G107), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n194), .A2(G104), .B1(KEYINPUT80), .B2(KEYINPUT3), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n187), .B(new_n191), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  OAI22_X1  g011(.A1(new_n194), .A2(G104), .B1(KEYINPUT80), .B2(KEYINPUT3), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n192), .B1(new_n190), .B2(G107), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n194), .A2(KEYINPUT80), .A3(KEYINPUT3), .A4(G104), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n196), .B(KEYINPUT4), .C1(new_n197), .C2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G113), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G113), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G116), .B(G119), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n207), .B(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n191), .B1(new_n193), .B2(new_n195), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(G101), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n202), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT83), .B1(new_n194), .B2(G104), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT83), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n190), .A3(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n194), .A2(G104), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n196), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n207), .A2(new_n208), .ZN(new_n221));
  INV_X1    g035(.A(G116), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G119), .ZN(new_n223));
  INV_X1    g037(.A(G119), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G116), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT5), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(G116), .ZN(new_n228));
  OAI21_X1  g042(.A(G113), .B1(new_n228), .B2(KEYINPUT5), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n221), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT85), .B1(new_n220), .B2(new_n230), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n201), .A2(new_n187), .B1(new_n218), .B2(G101), .ZN(new_n232));
  INV_X1    g046(.A(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n208), .A2(KEYINPUT5), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n233), .A2(new_n234), .B1(new_n208), .B2(new_n207), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT85), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n213), .A2(new_n231), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n213), .A2(new_n231), .A3(new_n239), .A4(new_n237), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(KEYINPUT6), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n246));
  OAI21_X1  g060(.A(G128), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(KEYINPUT64), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G143), .ZN(new_n250));
  AOI21_X1  g064(.A(G146), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n247), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G125), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n250), .A3(G146), .ZN(new_n256));
  INV_X1    g070(.A(new_n245), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n254), .A2(new_n255), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n251), .B2(new_n253), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n256), .A2(new_n263), .A3(new_n257), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n255), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G224), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n270), .B(KEYINPUT86), .Z(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n262), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n267), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G125), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n271), .B1(new_n275), .B2(new_n261), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n238), .A2(new_n278), .A3(new_n240), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n243), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(G210), .B1(G237), .B2(G902), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n239), .B(KEYINPUT8), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n232), .A2(new_n235), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n220), .A2(new_n230), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n270), .A2(KEYINPUT7), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n262), .B2(new_n268), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n261), .A4(new_n270), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n289), .B2(new_n242), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n280), .A2(new_n281), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n281), .B1(new_n280), .B2(new_n290), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G214), .B1(G237), .B2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G952), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(G953), .ZN(new_n297));
  NAND2_X1  g111(.A1(G234), .A2(G237), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(G902), .A3(G953), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT21), .B(G898), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n293), .A2(new_n295), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT9), .B(G234), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT79), .ZN(new_n307));
  OAI21_X1  g121(.A(G221), .B1(new_n307), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G469), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(G110), .B(G140), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n269), .A2(G227), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n316));
  INV_X1    g130(.A(G137), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT11), .A2(G134), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT65), .A2(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT11), .A2(G134), .ZN(new_n322));
  NOR2_X1   g136(.A1(KEYINPUT11), .A2(G134), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(G137), .ZN(new_n324));
  AND2_X1   g138(.A1(KEYINPUT66), .A2(G131), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT66), .A2(G131), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT67), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n321), .A2(new_n324), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G131), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n329), .B1(new_n321), .B2(new_n324), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n212), .A2(new_n267), .A3(new_n266), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT10), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n254), .B2(new_n260), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n335), .A2(new_n202), .B1(new_n232), .B2(new_n337), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n256), .A2(new_n257), .ZN(new_n340));
  OAI21_X1  g154(.A(G128), .B1(new_n251), .B2(new_n246), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n336), .B1(new_n342), .B2(new_n220), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n334), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n274), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n202), .A3(new_n212), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n337), .A2(new_n232), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n343), .A2(new_n334), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n315), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n315), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n341), .A2(new_n340), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n220), .B1(new_n352), .B2(new_n260), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n254), .A2(new_n260), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(new_n232), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT12), .B(new_n333), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n220), .A2(new_n254), .A3(new_n260), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n342), .B2(new_n220), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT12), .B1(new_n359), .B2(new_n333), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n351), .B(new_n348), .C1(new_n357), .C2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(G902), .B1(new_n350), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n312), .B1(new_n362), .B2(new_n310), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n348), .B1(new_n357), .B2(new_n360), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n315), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n346), .A2(new_n347), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n353), .A2(KEYINPUT10), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n333), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n348), .A2(new_n351), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT84), .B1(new_n348), .B2(new_n351), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n365), .B(G469), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n309), .B1(new_n363), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n305), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G217), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n307), .A2(new_n376), .A3(G953), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(KEYINPUT89), .A2(G122), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(KEYINPUT89), .A2(G122), .ZN(new_n381));
  OAI21_X1  g195(.A(G116), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n222), .A2(G122), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n194), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n248), .A2(new_n250), .A3(G128), .ZN(new_n385));
  INV_X1    g199(.A(G134), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n258), .A2(G143), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n386), .B1(new_n385), .B2(new_n387), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n384), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT90), .ZN(new_n392));
  INV_X1    g206(.A(G122), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n392), .B(KEYINPUT14), .C1(new_n393), .C2(G116), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n392), .B1(new_n383), .B2(KEYINPUT14), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n382), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT91), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n393), .A2(G116), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(KEYINPUT91), .B(new_n382), .C1(new_n395), .C2(new_n396), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n391), .B1(new_n404), .B2(G107), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n385), .A2(KEYINPUT13), .A3(new_n387), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n406), .B(G134), .C1(KEYINPUT13), .C2(new_n385), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n393), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n222), .B1(new_n409), .B2(new_n379), .ZN(new_n410));
  OAI21_X1  g224(.A(G107), .B1(new_n410), .B2(new_n400), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n384), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n407), .A2(new_n412), .A3(new_n388), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n378), .B1(new_n405), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n403), .A2(new_n402), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n194), .B1(new_n416), .B2(new_n399), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n413), .B(new_n377), .C1(new_n417), .C2(new_n391), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n415), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(KEYINPUT92), .B(new_n378), .C1(new_n405), .C2(new_n414), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n311), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT93), .ZN(new_n423));
  INV_X1    g237(.A(G478), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT93), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n420), .A2(new_n426), .A3(new_n311), .A4(new_n421), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n422), .B2(new_n425), .ZN(new_n429));
  XNOR2_X1  g243(.A(G113), .B(G122), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(new_n190), .ZN(new_n431));
  XNOR2_X1  g245(.A(G125), .B(G140), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT75), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n432), .A2(new_n434), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n252), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n432), .A2(KEYINPUT16), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n255), .A2(G140), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n438), .B(G146), .C1(KEYINPUT16), .C2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G237), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n441), .A2(new_n269), .A3(G143), .A4(G214), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n248), .A2(new_n250), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n441), .A2(new_n269), .A3(G214), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n327), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n437), .A2(new_n440), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n433), .A2(new_n252), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n252), .B2(new_n432), .ZN(new_n450));
  NAND2_X1  g264(.A1(KEYINPUT18), .A2(G131), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n445), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n431), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n438), .B1(KEYINPUT16), .B2(new_n439), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n252), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n445), .A2(KEYINPUT17), .A3(new_n446), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n440), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n445), .B(new_n327), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT17), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n458), .A2(KEYINPUT87), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n456), .A2(new_n457), .A3(new_n462), .A4(new_n440), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n461), .A2(new_n463), .B1(new_n450), .B2(new_n452), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n454), .B1(new_n464), .B2(new_n431), .ZN(new_n465));
  NOR2_X1   g279(.A1(G475), .A2(G902), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT20), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n461), .A2(new_n463), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n431), .A3(new_n453), .ZN(new_n470));
  INV_X1    g284(.A(new_n454), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n466), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n470), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n464), .A2(new_n431), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n311), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT88), .B(G475), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n375), .A2(new_n429), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(G472), .A2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n333), .A2(new_n345), .ZN(new_n485));
  INV_X1    g299(.A(new_n209), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n318), .A2(new_n386), .A3(new_n320), .ZN(new_n487));
  INV_X1    g301(.A(G131), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(G134), .B2(G137), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n328), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n354), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n485), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT28), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n321), .A2(new_n324), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT67), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(G131), .A3(new_n330), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n274), .B1(new_n498), .B2(new_n328), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n491), .A2(new_n354), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n209), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n493), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT69), .B1(new_n502), .B2(KEYINPUT28), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n504));
  AOI211_X1 g318(.A(new_n504), .B(new_n494), .C1(new_n501), .C2(new_n493), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n495), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n441), .A2(new_n269), .A3(G210), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT27), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(G101), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT30), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n485), .B2(new_n492), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n209), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(KEYINPUT68), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n493), .A3(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n499), .A2(new_n500), .A3(new_n209), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT30), .B1(new_n499), .B2(new_n500), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n485), .A2(new_n514), .A3(new_n492), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n520), .B1(new_n523), .B2(new_n209), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n517), .A2(KEYINPUT31), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n519), .A2(KEYINPUT31), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n484), .B1(new_n512), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT70), .B1(new_n527), .B2(KEYINPUT32), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n486), .B1(new_n485), .B2(new_n492), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT28), .B1(new_n520), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n504), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n502), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n510), .B1(new_n533), .B2(new_n495), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n519), .A2(KEYINPUT31), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n524), .A2(new_n525), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n483), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT70), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT32), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n511), .B1(new_n493), .B2(new_n494), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n531), .B2(new_n532), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT29), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n524), .B2(new_n510), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n542), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n516), .A2(new_n493), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT29), .B1(new_n549), .B2(new_n511), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n543), .B1(new_n503), .B2(new_n505), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT71), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n530), .A2(KEYINPUT29), .A3(new_n543), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT72), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT72), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n530), .A2(new_n555), .A3(KEYINPUT29), .A4(new_n543), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n548), .A2(new_n552), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G472), .ZN(new_n559));
  OAI211_X1 g373(.A(KEYINPUT32), .B(new_n483), .C1(new_n534), .C2(new_n537), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n528), .A2(new_n541), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n376), .B1(G234), .B2(new_n311), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n456), .A2(new_n440), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n224), .B2(G128), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n258), .A2(KEYINPUT73), .A3(G119), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n224), .A2(G128), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT24), .B(G110), .Z(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT23), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n224), .B2(G128), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n258), .A2(KEYINPUT23), .A3(G119), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G110), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n563), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G110), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n572), .A2(new_n573), .A3(new_n577), .A4(new_n567), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n578), .A2(KEYINPUT74), .ZN(new_n579));
  OAI22_X1  g393(.A1(new_n568), .A2(new_n569), .B1(new_n578), .B2(KEYINPUT74), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n449), .B(new_n440), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT22), .B(G137), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n576), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n576), .B2(new_n581), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT25), .B1(new_n589), .B2(new_n311), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n591));
  NOR4_X1   g405(.A1(new_n587), .A2(new_n588), .A3(new_n591), .A4(G902), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n562), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n562), .A2(G902), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n594), .B(KEYINPUT78), .Z(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n482), .A2(new_n561), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(new_n187), .Z(G3));
  INV_X1    g415(.A(new_n292), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n280), .A2(new_n290), .A3(new_n281), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n295), .B1(new_n291), .B2(KEYINPUT94), .ZN(new_n606));
  INV_X1    g420(.A(new_n304), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n420), .A2(new_n610), .A3(new_n421), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n415), .A2(new_n418), .A3(KEYINPUT33), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(G478), .A3(new_n311), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n481), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT95), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT95), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n614), .A2(new_n481), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n608), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n311), .B1(new_n534), .B2(new_n537), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n527), .B1(new_n620), .B2(G472), .ZN(new_n621));
  INV_X1    g435(.A(new_n361), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n351), .B1(new_n368), .B2(new_n348), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n310), .B(new_n311), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n312), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n373), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n308), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n598), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n619), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  AOI22_X1  g445(.A1(new_n468), .A2(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n429), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n608), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n621), .A3(new_n628), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  NAND2_X1  g451(.A1(new_n576), .A2(new_n581), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n638), .A2(KEYINPUT96), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(KEYINPUT96), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT36), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n586), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n639), .A2(new_n642), .A3(new_n586), .A4(new_n640), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n596), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n593), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n482), .A2(new_n621), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  NAND3_X1  g464(.A1(new_n626), .A2(new_n647), .A3(new_n308), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n605), .A2(new_n606), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n300), .B1(new_n302), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n633), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n528), .A2(new_n541), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n559), .A2(new_n560), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n653), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  NAND2_X1  g474(.A1(new_n549), .A2(new_n510), .ZN(new_n661));
  INV_X1    g475(.A(new_n502), .ZN(new_n662));
  AOI21_X1  g476(.A(G902), .B1(new_n662), .B2(new_n511), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n527), .A2(KEYINPUT32), .B1(G472), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n528), .A3(new_n541), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT97), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT97), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n665), .A2(new_n528), .A3(new_n541), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n293), .B(KEYINPUT38), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n429), .A2(new_n481), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n671), .A2(new_n672), .A3(new_n295), .A4(new_n647), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n670), .A2(KEYINPUT98), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n655), .B(KEYINPUT39), .Z(new_n675));
  NAND2_X1  g489(.A1(new_n374), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT40), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT98), .B1(new_n670), .B2(new_n673), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(new_n443), .Z(G45));
  INV_X1    g495(.A(new_n655), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n614), .A2(new_n481), .A3(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n683), .A2(new_n651), .A3(new_n652), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n561), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  OR2_X1    g500(.A1(new_n362), .A2(new_n310), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n308), .A3(new_n624), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n619), .A2(new_n561), .A3(new_n599), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G15));
  NAND4_X1  g506(.A1(new_n561), .A2(new_n634), .A3(new_n599), .A4(new_n689), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  INV_X1    g508(.A(new_n647), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n429), .A2(new_n695), .A3(new_n481), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n652), .A2(new_n688), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n561), .A2(new_n607), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  NAND2_X1  g513(.A1(new_n530), .A2(new_n495), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n511), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n484), .B1(new_n526), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n620), .B2(G472), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(new_n599), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n672), .A2(new_n652), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n607), .A3(new_n689), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  INV_X1    g521(.A(new_n683), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n697), .A2(new_n708), .A3(new_n647), .A4(new_n703), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  INV_X1    g524(.A(KEYINPUT101), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n560), .A2(KEYINPUT100), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n527), .A2(new_n714), .A3(KEYINPUT32), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n558), .A2(G472), .B1(new_n538), .B2(new_n540), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n598), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT99), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n293), .A2(new_n294), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n719), .B1(new_n627), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n374), .A2(KEYINPUT99), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n708), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n712), .B1(new_n718), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT99), .B1(new_n374), .B2(new_n722), .ZN(new_n727));
  AND4_X1   g541(.A1(KEYINPUT99), .A2(new_n722), .A3(new_n308), .A4(new_n626), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n683), .A2(KEYINPUT42), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n561), .A3(new_n599), .A4(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n711), .B1(new_n726), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n538), .A2(new_n540), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n713), .A2(new_n559), .A3(new_n715), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n599), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT42), .B1(new_n736), .B2(new_n724), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(KEYINPUT101), .A3(new_n731), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT102), .B(G131), .Z(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G33));
  NAND4_X1  g555(.A1(new_n729), .A2(new_n561), .A3(new_n599), .A4(new_n656), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NAND2_X1  g557(.A1(new_n614), .A2(new_n632), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n621), .A2(new_n695), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n722), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(KEYINPUT103), .B(new_n722), .C1(new_n748), .C2(new_n749), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n365), .B1(new_n371), .B2(new_n372), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n310), .B1(new_n754), .B2(new_n755), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n312), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n758), .A2(KEYINPUT46), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n624), .B1(new_n758), .B2(KEYINPUT46), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n308), .B(new_n675), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n749), .B2(new_n748), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n752), .A2(new_n753), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  OAI21_X1  g578(.A(new_n308), .B1(new_n759), .B2(new_n760), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n765), .B(new_n767), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n561), .A2(new_n599), .A3(new_n683), .A4(new_n720), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n746), .A2(new_n300), .ZN(new_n773));
  INV_X1    g587(.A(new_n704), .ZN(new_n774));
  OR4_X1    g588(.A1(KEYINPUT111), .A2(new_n773), .A3(new_n774), .A4(new_n720), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n746), .A2(new_n300), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n704), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT111), .B1(new_n777), .B2(new_n720), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n687), .A2(new_n624), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT106), .Z(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n308), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n775), .B(new_n778), .C1(new_n768), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n670), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n689), .A2(new_n722), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n598), .A3(new_n299), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n614), .A2(new_n481), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(KEYINPUT114), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(KEYINPUT114), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n782), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n689), .A2(KEYINPUT112), .A3(new_n295), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n688), .B2(new_n294), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n671), .A3(new_n793), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n773), .A2(new_n774), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n797), .B1(new_n795), .B2(new_n796), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n703), .A2(new_n647), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n773), .A2(new_n784), .ZN(new_n803));
  OAI22_X1  g617(.A1(new_n799), .A2(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n772), .B1(new_n790), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n803), .A2(new_n736), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT48), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n616), .A2(new_n618), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n783), .A2(new_n808), .A3(new_n785), .ZN(new_n809));
  INV_X1    g623(.A(new_n697), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n777), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n805), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n788), .A2(new_n789), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n803), .A2(new_n802), .ZN(new_n816));
  INV_X1    g630(.A(new_n800), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n817), .B2(new_n798), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n818), .A3(new_n782), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n814), .B1(new_n819), .B2(new_n772), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n790), .A2(new_n804), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(KEYINPUT115), .A3(KEYINPUT51), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n813), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n690), .A2(new_n693), .A3(new_n706), .A4(new_n698), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n633), .A2(new_n615), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n305), .A3(new_n621), .A4(new_n628), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n600), .A2(new_n648), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n627), .A2(new_n720), .A3(new_n655), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n696), .B(new_n830), .C1(new_n657), .C2(new_n658), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT107), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n729), .A2(new_n708), .A3(new_n801), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n561), .A2(KEYINPUT107), .A3(new_n696), .A4(new_n830), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n742), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n829), .A2(new_n836), .A3(new_n733), .A4(new_n738), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n659), .A2(new_n685), .A3(new_n709), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT108), .B1(new_n647), .B2(new_n655), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT108), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n593), .A2(new_n646), .A3(new_n841), .A4(new_n682), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n705), .A2(new_n843), .A3(new_n374), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n670), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n838), .A2(new_n839), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n659), .A2(new_n685), .A3(new_n709), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n844), .B1(new_n667), .B2(new_n669), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT52), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT53), .B1(new_n837), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n847), .A2(new_n850), .A3(KEYINPUT109), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT109), .B1(new_n847), .B2(new_n850), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n738), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT101), .B1(new_n737), .B2(new_n731), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n829), .A4(new_n836), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n852), .B(KEYINPUT54), .C1(new_n855), .C2(new_n860), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n690), .A2(new_n693), .A3(new_n698), .A4(new_n706), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n729), .A2(new_n561), .A3(new_n599), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n729), .A2(new_n599), .A3(new_n708), .A4(new_n735), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n863), .A2(new_n730), .B1(new_n864), .B2(KEYINPUT42), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT110), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n737), .A2(new_n731), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT110), .B1(new_n868), .B2(new_n825), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n828), .A2(new_n859), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n836), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n870), .B(new_n872), .C1(new_n853), .C2(new_n854), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n859), .B1(new_n837), .B2(new_n851), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n823), .A2(new_n824), .A3(new_n861), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(G953), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n823), .A2(KEYINPUT116), .A3(new_n861), .A4(new_n876), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n297), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n780), .A2(KEYINPUT49), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n780), .A2(KEYINPUT49), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n671), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT105), .ZN(new_n884));
  OR4_X1    g698(.A1(new_n598), .A2(new_n744), .A3(new_n295), .A4(new_n309), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n881), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n886), .B(new_n783), .C1(new_n884), .C2(new_n885), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n878), .A2(new_n880), .A3(new_n887), .ZN(G75));
  NAND2_X1  g702(.A1(new_n873), .A2(new_n875), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(G210), .A3(G902), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT117), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT55), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n243), .A2(new_n279), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n277), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT55), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n890), .A2(new_n898), .A3(new_n893), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n895), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n897), .B1(new_n895), .B2(new_n899), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n296), .A2(G953), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT118), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(G51));
  NAND2_X1  g719(.A1(new_n889), .A2(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n876), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n312), .B(KEYINPUT57), .Z(new_n909));
  OAI22_X1  g723(.A1(new_n908), .A2(new_n909), .B1(new_n623), .B2(new_n622), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n889), .A2(G902), .A3(new_n756), .A4(new_n757), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(G54));
  AND4_X1   g726(.A1(KEYINPUT58), .A2(new_n889), .A3(G475), .A4(G902), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n913), .A2(new_n914), .A3(new_n472), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n913), .B2(new_n472), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n904), .B1(new_n913), .B2(new_n472), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G60));
  NAND2_X1  g732(.A1(new_n861), .A2(new_n876), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n611), .A2(new_n612), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n921), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n904), .B1(new_n907), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n921), .B1(new_n861), .B2(new_n876), .ZN(new_n929));
  INV_X1    g743(.A(new_n925), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT120), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n926), .A2(new_n928), .A3(new_n931), .A4(KEYINPUT121), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT60), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT122), .B1(new_n889), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n589), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n889), .A2(KEYINPUT122), .A3(new_n939), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n945), .B(new_n938), .C1(new_n873), .C2(new_n875), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n645), .B(new_n644), .C1(new_n940), .C2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n944), .A2(new_n947), .A3(new_n903), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n944), .A2(new_n947), .A3(KEYINPUT61), .A4(new_n903), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(G66));
  INV_X1    g766(.A(G224), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n303), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n829), .B2(G953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n896), .B1(G898), .B2(new_n269), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  NAND2_X1  g771(.A1(new_n435), .A2(new_n436), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n523), .B(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n960), .A2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n838), .B1(new_n678), .B2(new_n679), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n676), .A2(new_n720), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n561), .A2(new_n964), .A3(new_n599), .A4(new_n826), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(new_n763), .A3(new_n770), .A4(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n961), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n654), .A2(new_n269), .ZN(new_n970));
  INV_X1    g784(.A(new_n761), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n705), .A3(new_n718), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n763), .A2(new_n770), .A3(new_n838), .A4(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT123), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n858), .A2(new_n974), .A3(new_n742), .ZN(new_n975));
  INV_X1    g789(.A(new_n742), .ZN(new_n976));
  OAI21_X1  g790(.A(KEYINPUT123), .B1(new_n739), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n973), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n970), .B1(new_n978), .B2(new_n269), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n968), .B(new_n969), .C1(new_n979), .C2(new_n959), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n968), .B1(new_n979), .B2(new_n959), .ZN(new_n983));
  INV_X1    g797(.A(new_n969), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT124), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n983), .A2(KEYINPUT124), .A3(new_n984), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n982), .B1(new_n985), .B2(new_n987), .ZN(G72));
  NOR2_X1   g802(.A1(new_n966), .A2(new_n967), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n829), .ZN(new_n990));
  XNOR2_X1  g804(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n991));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n661), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n524), .A2(new_n511), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT127), .Z(new_n996));
  NAND2_X1  g810(.A1(new_n978), .A2(new_n829), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(new_n993), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n852), .B1(new_n855), .B2(new_n860), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n661), .A2(new_n993), .A3(new_n995), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n903), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n994), .A2(new_n998), .A3(new_n1001), .ZN(G57));
endmodule


