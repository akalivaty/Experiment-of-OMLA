//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(G228gat), .ZN(new_n207));
  INV_X1    g006(.A(G233gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT73), .ZN(new_n213));
  INV_X1    g012(.A(G211gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n215));
  INV_X1    g014(.A(G218gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n213), .B1(new_n219), .B2(KEYINPUT22), .ZN(new_n220));
  AND2_X1   g019(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n222));
  OAI21_X1  g021(.A(G211gat), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(KEYINPUT73), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(G197gat), .B(G204gat), .Z(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n212), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n212), .ZN(new_n230));
  AOI211_X1 g029(.A(new_n227), .B(new_n230), .C1(new_n220), .C2(new_n225), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n211), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n223), .A2(KEYINPUT73), .A3(new_n224), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT73), .B1(new_n223), .B2(new_n224), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n228), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n230), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n226), .A2(new_n228), .A3(new_n212), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(KEYINPUT74), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239));
  INV_X1    g038(.A(G141gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G148gat), .ZN(new_n241));
  INV_X1    g040(.A(G148gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G141gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G155gat), .B(G162gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n240), .A2(G148gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT77), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G162gat), .ZN(new_n250));
  INV_X1    g049(.A(G155gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT78), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT78), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G155gat), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n250), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT2), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT79), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT79), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT78), .B(G155gat), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n258), .B(KEYINPUT2), .C1(new_n259), .C2(new_n250), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n249), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n242), .A2(G141gat), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT75), .B1(new_n262), .B2(new_n247), .ZN(new_n263));
  NAND2_X1  g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(KEYINPUT2), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT75), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n241), .A2(new_n243), .A3(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n263), .A2(new_n265), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n246), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n261), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n232), .A2(new_n238), .B1(new_n239), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n261), .A2(new_n273), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n239), .B1(new_n229), .B2(new_n231), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(new_n274), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n210), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT86), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n239), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n229), .A2(new_n231), .A3(new_n211), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT74), .B1(new_n236), .B2(new_n237), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n261), .A2(new_n273), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT29), .B1(new_n236), .B2(new_n237), .ZN(new_n287));
  INV_X1    g086(.A(new_n274), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT86), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(new_n210), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n281), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n261), .A2(new_n273), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n261), .B2(new_n273), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(KEYINPUT3), .B2(new_n287), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n285), .A2(new_n298), .A3(new_n209), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n206), .B1(new_n293), .B2(new_n300), .ZN(new_n301));
  AOI211_X1 g100(.A(G22gat), .B(new_n299), .C1(new_n281), .C2(new_n292), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n205), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n291), .B1(new_n290), .B2(new_n210), .ZN(new_n304));
  AOI211_X1 g103(.A(KEYINPUT86), .B(new_n209), .C1(new_n285), .C2(new_n289), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n300), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G22gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n293), .A2(new_n206), .A3(new_n300), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n204), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n286), .A2(KEYINPUT80), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n261), .A2(new_n273), .A3(new_n294), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(KEYINPUT3), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G127gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(KEYINPUT69), .ZN(new_n316));
  XNOR2_X1  g115(.A(G113gat), .B(G120gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(KEYINPUT1), .ZN(new_n318));
  INV_X1    g117(.A(G134gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  INV_X1    g119(.A(G113gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n321), .A2(G120gat), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(G113gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n320), .B(new_n315), .C1(new_n322), .C2(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n318), .A2(new_n319), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n319), .B1(new_n318), .B2(new_n325), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n314), .A2(new_n328), .A3(new_n275), .ZN(new_n329));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(KEYINPUT5), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n261), .B(new_n273), .C1(new_n326), .C2(new_n327), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT82), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n325), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G134gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n319), .A3(new_n325), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n273), .A4(new_n261), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n334), .A2(KEYINPUT4), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT83), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(new_n333), .B2(KEYINPUT4), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n277), .A2(KEYINPUT83), .A3(new_n344), .A4(new_n338), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n329), .B(new_n332), .C1(new_n341), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT84), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n340), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n343), .B(new_n345), .C1(new_n350), .C2(new_n344), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n351), .A2(KEYINPUT84), .A3(new_n329), .A4(new_n332), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n297), .A2(new_n328), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(new_n334), .A3(new_n340), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n356), .B2(new_n331), .ZN(new_n357));
  INV_X1    g156(.A(new_n333), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n331), .B1(new_n358), .B2(KEYINPUT4), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n329), .B(new_n359), .C1(new_n350), .C2(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n353), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(G57gat), .B(G85gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(KEYINPUT6), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT85), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(new_n353), .B2(new_n361), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT6), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n370), .A2(KEYINPUT6), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n349), .A2(new_n352), .B1(new_n357), .B2(new_n360), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n366), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n369), .A2(new_n372), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT66), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT26), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n382), .A2(new_n385), .B1(G183gat), .B2(G190gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(G183gat), .ZN(new_n388));
  INV_X1    g187(.A(G183gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(KEYINPUT27), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT68), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(KEYINPUT27), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT68), .ZN(new_n393));
  AOI21_X1  g192(.A(G190gat), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT28), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n387), .A2(G183gat), .ZN(new_n396));
  INV_X1    g195(.A(G190gat), .ZN(new_n397));
  AND4_X1   g196(.A1(KEYINPUT28), .A2(new_n392), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n386), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n384), .B1(KEYINPUT65), .B2(KEYINPUT23), .ZN(new_n400));
  NAND2_X1  g199(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  OAI22_X1  g201(.A1(new_n400), .A2(new_n402), .B1(G169gat), .B2(G176gat), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(G183gat), .A2(G190gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT67), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n379), .A2(KEYINPUT23), .A3(new_n381), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n403), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT25), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT25), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n406), .A2(new_n408), .ZN(new_n416));
  INV_X1    g215(.A(G169gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT64), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT64), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G169gat), .ZN(new_n420));
  INV_X1    g219(.A(G176gat), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT23), .A4(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n403), .A2(new_n415), .A3(new_n416), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n414), .A3(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(new_n424), .B2(new_n239), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(new_n283), .B2(new_n284), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n283), .A2(new_n284), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n426), .B2(new_n427), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n435), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n429), .A2(new_n431), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(KEYINPUT30), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n432), .A2(new_n440), .A3(new_n435), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n311), .B1(new_n376), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n424), .A2(new_n338), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n403), .A2(new_n415), .A3(new_n422), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n447), .A2(new_n416), .B1(new_n413), .B2(KEYINPUT25), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(new_n328), .A3(new_n399), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G227gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n208), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n445), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  AOI211_X1 g253(.A(KEYINPUT34), .B(new_n452), .C1(new_n446), .C2(new_n449), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n446), .A2(new_n449), .A3(new_n452), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT32), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(G15gat), .B(G43gat), .Z(new_n461));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n463), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n457), .B(KEYINPUT32), .C1(new_n459), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n456), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT70), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT70), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n456), .A2(new_n464), .A3(new_n469), .A4(new_n466), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n464), .A2(new_n466), .ZN(new_n472));
  INV_X1    g271(.A(new_n456), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT36), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n474), .A2(KEYINPUT71), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT71), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n472), .A2(new_n473), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n481), .A2(new_n471), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n477), .B1(new_n482), .B2(KEYINPUT36), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n369), .A2(new_n372), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n435), .B1(new_n432), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT38), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n429), .A2(new_n431), .A3(KEYINPUT37), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n488), .A2(new_n489), .B1(new_n490), .B2(new_n486), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n486), .A2(KEYINPUT87), .A3(new_n489), .A4(new_n490), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n436), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n362), .A2(new_n367), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n496), .A3(new_n375), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n484), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n301), .A2(new_n302), .A3(new_n205), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n204), .B1(new_n307), .B2(new_n308), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n355), .A2(new_n334), .A3(new_n340), .A4(new_n330), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT39), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n329), .B1(new_n341), .B2(new_n346), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(new_n331), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT39), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n507), .A3(new_n331), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n366), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n502), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(new_n331), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(KEYINPUT39), .A3(new_n503), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n512), .A2(KEYINPUT40), .A3(new_n366), .A4(new_n508), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n439), .B(new_n441), .C1(new_n374), .C2(new_n366), .ZN(new_n515));
  OAI22_X1  g314(.A1(new_n500), .A2(new_n501), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n444), .B(new_n483), .C1(new_n499), .C2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT35), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n519));
  AOI211_X1 g318(.A(new_n519), .B(new_n475), .C1(new_n309), .C2(new_n303), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT88), .B1(new_n310), .B2(new_n476), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n443), .B1(new_n484), .B2(new_n497), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n371), .B1(new_n370), .B2(KEYINPUT6), .ZN(new_n525));
  NOR4_X1   g324(.A1(new_n374), .A2(KEYINPUT85), .A3(new_n496), .A4(new_n366), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n497), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n481), .A2(new_n471), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n529));
  AND4_X1   g328(.A1(new_n527), .A2(new_n529), .A3(new_n310), .A4(new_n442), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n517), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT15), .ZN(new_n532));
  XNOR2_X1  g331(.A(G43gat), .B(G50gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n534), .B2(new_n533), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n537), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT14), .B(G29gat), .ZN(new_n539));
  INV_X1    g338(.A(G36gat), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n536), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT17), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  XNOR2_X1  g347(.A(G15gat), .B(G22gat), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n549), .A2(G1gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT16), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n551), .B2(G1gat), .ZN(new_n552));
  INV_X1    g351(.A(G8gat), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n553), .A2(KEYINPUT90), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(KEYINPUT90), .A3(new_n553), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(KEYINPUT90), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n550), .A2(new_n552), .A3(new_n557), .A4(new_n554), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT91), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n561), .A3(new_n558), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n546), .A2(new_n548), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n556), .A2(KEYINPUT92), .A3(new_n558), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n566), .A2(new_n567), .A3(new_n544), .A4(new_n542), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n545), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n568), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n564), .B(KEYINPUT13), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n563), .A2(new_n568), .A3(KEYINPUT18), .A4(new_n564), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G197gat), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT11), .B(G169gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT12), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n571), .A2(new_n576), .A3(new_n583), .A4(new_n577), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(KEYINPUT93), .A3(new_n586), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n531), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g394(.A(KEYINPUT102), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G99gat), .ZN(new_n598));
  INV_X1    g397(.A(G106gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT99), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n600), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G85gat), .A2(G92gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT7), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  INV_X1    g408(.A(G92gat), .ZN(new_n610));
  AOI22_X1  g409(.A1(KEYINPUT8), .A2(new_n601), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n606), .B(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n546), .A2(new_n548), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n545), .B2(new_n613), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n597), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n620));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n614), .B(new_n617), .C1(new_n545), .C2(new_n613), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n597), .A3(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n595), .A2(new_n596), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n623), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n623), .B2(new_n626), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(G71gat), .A2(G78gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(G71gat), .A2(G78gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G57gat), .B(G64gat), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT9), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(G57gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(G64gat), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT94), .B(G57gat), .Z(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(G64gat), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n635), .B1(KEYINPUT9), .B2(new_n636), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT21), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n572), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G183gat), .B(G211gat), .Z(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n646), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(G231gat), .A3(G233gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(G127gat), .B(G155gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT96), .Z(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G231gat), .A2(G233gat), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n646), .A2(new_n663), .A3(new_n657), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n659), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n659), .B2(new_n664), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n655), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n665), .A2(new_n666), .A3(new_n655), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n654), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n669), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n671), .A2(new_n652), .A3(new_n653), .A4(new_n667), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n646), .B1(KEYINPUT103), .B2(new_n606), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n613), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n603), .A2(new_n605), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n612), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n606), .A2(KEYINPUT103), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n646), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(G230gat), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n208), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT10), .B1(new_n675), .B2(new_n679), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT10), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n613), .A2(new_n688), .A3(new_n646), .ZN(new_n689));
  OAI22_X1  g488(.A1(new_n687), .A2(new_n689), .B1(new_n682), .B2(new_n208), .ZN(new_n690));
  XNOR2_X1  g489(.A(G120gat), .B(G148gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n691), .B(new_n692), .Z(new_n693));
  NAND3_X1  g492(.A1(new_n681), .A2(KEYINPUT104), .A3(new_n683), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n686), .A2(new_n690), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n690), .A2(new_n684), .ZN(new_n696));
  INV_X1    g495(.A(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n634), .A2(new_n673), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n592), .A2(new_n376), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g503(.A(KEYINPUT16), .B(G8gat), .Z(new_n705));
  NAND4_X1  g504(.A1(new_n592), .A2(new_n443), .A3(new_n702), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n592), .A2(new_n702), .ZN(new_n707));
  OAI21_X1  g506(.A(G8gat), .B1(new_n707), .B2(new_n442), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n706), .ZN(new_n709));
  MUX2_X1   g508(.A(new_n706), .B(new_n709), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g509(.A(G15gat), .B1(new_n707), .B2(new_n483), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n528), .A2(G15gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n707), .B2(new_n712), .ZN(G1326gat));
  NOR2_X1   g512(.A1(new_n707), .A2(new_n310), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  NOR3_X1   g515(.A1(new_n634), .A2(new_n673), .A3(new_n699), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n531), .A2(new_n591), .A3(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n718), .A2(G29gat), .A3(new_n527), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT45), .Z(new_n720));
  XOR2_X1   g519(.A(new_n699), .B(KEYINPUT105), .Z(new_n721));
  INV_X1    g520(.A(new_n673), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n587), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT106), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n476), .B1(new_n500), .B2(new_n501), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n519), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n310), .A2(KEYINPUT88), .A3(new_n476), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n523), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n530), .B1(new_n729), .B2(KEYINPUT35), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n516), .B1(new_n376), .B2(new_n494), .ZN(new_n731));
  MUX2_X1   g530(.A(new_n482), .B(new_n475), .S(KEYINPUT36), .Z(new_n732));
  AOI21_X1  g531(.A(new_n310), .B1(new_n527), .B2(new_n442), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n725), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(KEYINPUT107), .B(new_n517), .C1(new_n524), .C2(new_n530), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n632), .B2(new_n633), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n623), .A2(new_n626), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n629), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(KEYINPUT108), .A3(new_n631), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n735), .A2(new_n736), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n634), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n730), .B2(new_n734), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n724), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G29gat), .B1(new_n749), .B2(new_n527), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n720), .A2(new_n750), .ZN(G1328gat));
  NOR3_X1   g550(.A1(new_n718), .A2(G36gat), .A3(new_n442), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT46), .ZN(new_n753));
  OAI21_X1  g552(.A(G36gat), .B1(new_n749), .B2(new_n442), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1329gat));
  INV_X1    g554(.A(G43gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n748), .B2(new_n732), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n718), .A2(G43gat), .A3(new_n528), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n757), .B2(new_n759), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1330gat));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n763));
  INV_X1    g562(.A(new_n724), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(new_n311), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G50gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  INV_X1    g567(.A(G50gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n311), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n718), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(KEYINPUT109), .A2(KEYINPUT48), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n767), .A2(new_n768), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n769), .B1(new_n748), .B2(new_n311), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n774), .B(new_n775), .C1(new_n776), .C2(new_n771), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n773), .A2(new_n777), .ZN(G1331gat));
  NOR4_X1   g577(.A1(new_n721), .A2(new_n745), .A3(new_n587), .A4(new_n722), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n735), .A2(new_n736), .A3(new_n376), .A4(new_n779), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(new_n643), .ZN(G1332gat));
  NAND3_X1  g583(.A1(new_n735), .A2(new_n736), .A3(new_n779), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n785), .A2(KEYINPUT111), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(KEYINPUT111), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n443), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT49), .B(G64gat), .Z(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n788), .B2(new_n790), .ZN(G1333gat));
  NAND4_X1  g590(.A1(new_n786), .A2(G71gat), .A3(new_n732), .A4(new_n787), .ZN(new_n792));
  INV_X1    g591(.A(G71gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n785), .B2(new_n528), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n792), .A2(KEYINPUT50), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT50), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(G1334gat));
  NAND3_X1  g596(.A1(new_n786), .A2(new_n311), .A3(new_n787), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g598(.A1(new_n673), .A2(new_n587), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n699), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n744), .B2(new_n747), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n527), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  INV_X1    g604(.A(new_n800), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n746), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n531), .A2(KEYINPUT51), .A3(new_n745), .A4(new_n800), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n809), .A2(new_n609), .A3(new_n376), .A4(new_n699), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n804), .A2(new_n810), .ZN(G1336gat));
  NAND2_X1  g610(.A1(new_n802), .A2(new_n443), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G92gat), .ZN(new_n813));
  INV_X1    g612(.A(new_n721), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n610), .A3(new_n443), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT112), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(new_n809), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n816), .B(KEYINPUT113), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n812), .A2(G92gat), .B1(new_n809), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(G1337gat));
  OAI21_X1  g621(.A(G99gat), .B1(new_n803), .B2(new_n483), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n809), .A2(new_n598), .A3(new_n482), .A4(new_n699), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(G1338gat));
  AOI21_X1  g624(.A(new_n599), .B1(new_n802), .B2(new_n311), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n721), .A2(G106gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n809), .A2(new_n311), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n830), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT53), .B1(new_n832), .B2(new_n826), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1339gat));
  NAND2_X1  g633(.A1(new_n738), .A2(new_n741), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n690), .A2(KEYINPUT54), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n680), .A2(new_n688), .ZN(new_n837));
  INV_X1    g636(.A(new_n689), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n683), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n690), .A3(KEYINPUT54), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n836), .A2(new_n840), .A3(KEYINPUT55), .A4(new_n697), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n839), .A2(new_n690), .A3(KEYINPUT54), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n697), .B1(new_n690), .B2(KEYINPUT54), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n587), .A2(new_n695), .A3(new_n841), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n574), .A2(new_n575), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n564), .B1(new_n563), .B2(new_n568), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n582), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n699), .A2(new_n586), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n835), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n845), .A2(new_n695), .A3(new_n841), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n586), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n835), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n722), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n673), .A2(new_n631), .A3(new_n740), .ZN(new_n857));
  INV_X1    g656(.A(new_n587), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n857), .A2(KEYINPUT114), .A3(new_n858), .A4(new_n700), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n701), .B2(new_n587), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n376), .A2(new_n442), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n863), .A2(new_n310), .A3(new_n482), .A4(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n591), .ZN(new_n867));
  OAI21_X1  g666(.A(G113gat), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT115), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n863), .A2(new_n522), .A3(new_n865), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n587), .A2(new_n321), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(G1340gat));
  NOR3_X1   g671(.A1(new_n866), .A2(new_n323), .A3(new_n721), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n870), .A2(new_n700), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n323), .B2(new_n874), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n866), .B2(new_n722), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n673), .A2(new_n315), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n870), .B2(new_n877), .ZN(G1342gat));
  XOR2_X1   g677(.A(KEYINPUT69), .B(G134gat), .Z(new_n879));
  NOR3_X1   g678(.A1(new_n870), .A2(new_n634), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n882));
  OAI21_X1  g681(.A(G134gat), .B1(new_n866), .B2(new_n634), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G1343gat));
  NAND2_X1  g684(.A1(new_n863), .A2(new_n311), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n483), .A2(new_n376), .A3(new_n442), .ZN(new_n887));
  NOR4_X1   g686(.A1(new_n886), .A2(G141gat), .A3(new_n867), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n865), .A2(new_n483), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n835), .A2(new_n854), .ZN(new_n890));
  INV_X1    g689(.A(new_n850), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n841), .A2(new_n695), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n836), .A2(new_n697), .A3(new_n840), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT55), .B1(new_n893), .B2(KEYINPUT116), .ZN(new_n894));
  OR3_X1    g693(.A1(new_n843), .A2(KEYINPUT116), .A3(new_n844), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n891), .B1(new_n591), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n890), .B1(new_n897), .B2(new_n745), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n898), .A2(new_n722), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n859), .A2(new_n861), .ZN(new_n900));
  OAI211_X1 g699(.A(KEYINPUT57), .B(new_n311), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n889), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n587), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n888), .B1(new_n905), .B2(G141gat), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n240), .B1(new_n904), .B2(new_n591), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n888), .A2(KEYINPUT58), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n906), .A2(new_n907), .B1(new_n908), .B2(new_n909), .ZN(G1344gat));
  NOR2_X1   g709(.A1(new_n889), .A2(new_n700), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n911), .A2(new_n242), .A3(new_n311), .A4(new_n863), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT117), .Z(new_n913));
  XNOR2_X1  g712(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n854), .A2(new_n745), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n897), .B2(new_n745), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n722), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n867), .A2(new_n702), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n310), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n915), .B1(new_n920), .B2(KEYINPUT57), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n850), .B1(new_n858), .B2(new_n852), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n742), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n673), .B1(new_n923), .B2(new_n890), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT57), .B(new_n311), .C1(new_n924), .C2(new_n900), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n863), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n311), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n917), .A2(new_n722), .B1(new_n867), .B2(new_n702), .ZN(new_n930));
  OAI211_X1 g729(.A(KEYINPUT120), .B(new_n902), .C1(new_n930), .C2(new_n310), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n921), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n911), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n914), .B1(new_n933), .B2(G148gat), .ZN(new_n934));
  AOI211_X1 g733(.A(KEYINPUT59), .B(new_n242), .C1(new_n904), .C2(new_n699), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n913), .B1(new_n934), .B2(new_n935), .ZN(G1345gat));
  NOR2_X1   g735(.A1(new_n722), .A2(new_n259), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n886), .A2(new_n887), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n673), .ZN(new_n939));
  AOI22_X1  g738(.A1(new_n904), .A2(new_n937), .B1(new_n939), .B2(new_n259), .ZN(G1346gat));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n250), .A3(new_n745), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n904), .A2(new_n835), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n943), .B2(new_n250), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n944), .B(new_n945), .ZN(G1347gat));
  NOR2_X1   g745(.A1(new_n376), .A2(new_n442), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n863), .A2(new_n310), .A3(new_n482), .A4(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n867), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n376), .B1(new_n856), .B2(new_n862), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n443), .A3(new_n522), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n587), .A2(new_n418), .A3(new_n420), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1348gat));
  OAI21_X1  g752(.A(G176gat), .B1(new_n948), .B2(new_n721), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n699), .A2(new_n421), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n951), .B2(new_n955), .ZN(G1349gat));
  OAI21_X1  g755(.A(G183gat), .B1(new_n948), .B2(new_n722), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n673), .A2(new_n392), .A3(new_n396), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n951), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g759(.A(G190gat), .B1(new_n948), .B2(new_n634), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT61), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n835), .A2(new_n397), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n951), .B2(new_n963), .ZN(G1351gat));
  NAND3_X1  g763(.A1(new_n483), .A2(new_n311), .A3(new_n443), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n969), .A2(KEYINPUT123), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(KEYINPUT123), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(G197gat), .B1(new_n972), .B2(new_n587), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n947), .A2(new_n483), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n932), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n591), .A2(G197gat), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1352gat));
  NOR3_X1   g776(.A1(new_n969), .A2(G204gat), .A3(new_n700), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT62), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n932), .A2(new_n814), .A3(new_n974), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G204gat), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n980), .A2(new_n981), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(G1353gat));
  NAND3_X1  g784(.A1(new_n932), .A2(new_n673), .A3(new_n974), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(G211gat), .ZN(new_n987));
  NOR2_X1   g786(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n986), .B(G211gat), .C1(KEYINPUT126), .C2(KEYINPUT63), .ZN(new_n990));
  NAND2_X1  g789(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n722), .A2(G211gat), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n972), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(KEYINPUT125), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n972), .A2(new_n996), .A3(new_n993), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n992), .A2(new_n998), .ZN(G1354gat));
  NAND3_X1  g798(.A1(new_n970), .A2(new_n835), .A3(new_n971), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(new_n216), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n634), .B1(new_n217), .B2(new_n218), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n932), .A2(new_n974), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


