//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(G128), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n189), .B(new_n191), .C1(new_n192), .C2(KEYINPUT23), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G110), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT24), .B(G110), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT74), .B1(new_n188), .B2(G119), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n190), .A3(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n188), .A2(G119), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n194), .B1(new_n195), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(KEYINPUT75), .A3(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(KEYINPUT16), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n203), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n214), .A3(new_n211), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n201), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT77), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n200), .A2(new_n195), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n199), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G110), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n220), .A2(new_n189), .A3(new_n221), .A4(new_n191), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n203), .A2(new_n205), .A3(new_n214), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT76), .A4(new_n214), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n214), .B1(new_n209), .B2(new_n211), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n217), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n218), .A2(new_n222), .B1(new_n226), .B2(new_n227), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n213), .A2(new_n232), .A3(KEYINPUT77), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n216), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT22), .B(G137), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT68), .B(G953), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT78), .ZN(new_n238));
  INV_X1    g052(.A(G221), .ZN(new_n239));
  INV_X1    g053(.A(G234), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n238), .B1(new_n237), .B2(new_n241), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n236), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n244), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n242), .A3(new_n235), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n234), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT79), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT80), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n234), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n200), .A2(new_n195), .ZN(new_n256));
  INV_X1    g070(.A(new_n215), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n194), .B(new_n256), .C1(new_n257), .C2(new_n230), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n213), .A2(KEYINPUT77), .A3(new_n232), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT77), .B1(new_n213), .B2(new_n232), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT79), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT79), .B1(new_n245), .B2(new_n247), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT80), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n187), .B(new_n249), .C1(new_n255), .C2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT25), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n187), .A2(KEYINPUT25), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n234), .B2(new_n248), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n255), .B2(new_n265), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(KEYINPUT81), .B(new_n270), .C1(new_n255), .C2(new_n265), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n268), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G217), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(G234), .B2(new_n187), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n275), .A2(KEYINPUT82), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT82), .B1(new_n275), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n249), .B1(new_n255), .B2(new_n265), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n277), .A2(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n278), .A2(new_n279), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G214), .B1(G237), .B2(G902), .ZN(new_n285));
  OAI21_X1  g099(.A(G210), .B1(G237), .B2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n214), .A2(G143), .ZN(new_n288));
  INV_X1    g102(.A(G143), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G146), .ZN(new_n290));
  AND2_X1   g104(.A1(KEYINPUT0), .A2(G128), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G143), .B(G146), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT0), .B(G128), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G125), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n288), .A2(new_n290), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT1), .B1(new_n289), .B2(G146), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(G128), .A3(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n288), .B(new_n290), .C1(KEYINPUT1), .C2(new_n188), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n204), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G953), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G224), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n303), .B(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n308));
  INV_X1    g122(.A(G104), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G107), .ZN(new_n310));
  INV_X1    g124(.A(G101), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n309), .A2(G107), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT3), .B1(new_n314), .B2(KEYINPUT83), .ZN(new_n315));
  INV_X1    g129(.A(G107), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(KEYINPUT83), .A3(KEYINPUT3), .A4(G104), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n313), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(G104), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n311), .B1(new_n310), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT2), .A2(G113), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT66), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OR2_X1    g142(.A1(KEYINPUT2), .A2(G113), .ZN(new_n329));
  XNOR2_X1  g143(.A(G116), .B(G119), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n330), .A2(KEYINPUT5), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n190), .A2(G116), .ZN(new_n333));
  OAI21_X1  g147(.A(G113), .B1(new_n333), .B2(KEYINPUT5), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n323), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n316), .A2(G104), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n316), .A2(KEYINPUT83), .A3(G104), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n337), .B1(new_n340), .B2(new_n317), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n319), .B(KEYINPUT4), .C1(new_n341), .C2(new_n311), .ZN(new_n342));
  INV_X1    g156(.A(new_n341), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(G101), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n329), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G116), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G119), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n333), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n353), .A2(new_n331), .A3(KEYINPUT67), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT67), .B1(new_n353), .B2(new_n331), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n336), .B1(new_n346), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G110), .B(G122), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AND4_X1   g173(.A1(new_n308), .A2(new_n357), .A3(KEYINPUT6), .A4(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n342), .B(new_n345), .C1(new_n354), .C2(new_n355), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n358), .B1(new_n361), .B2(new_n336), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT6), .B1(new_n362), .B2(new_n308), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n336), .A3(new_n358), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT85), .ZN(new_n366));
  INV_X1    g180(.A(new_n362), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n361), .A2(new_n368), .A3(new_n336), .A4(new_n358), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n307), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n369), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n323), .B(new_n335), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n358), .B(KEYINPUT8), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n305), .A2(KEYINPUT7), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n297), .A2(new_n302), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n297), .A2(KEYINPUT87), .A3(new_n302), .A4(new_n376), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n303), .A2(KEYINPUT7), .A3(new_n305), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n375), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(G902), .B1(new_n372), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n287), .B1(new_n371), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n362), .A2(new_n308), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n362), .A2(new_n308), .A3(KEYINPUT6), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n370), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n306), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n384), .A3(new_n286), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT9), .B(G234), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n239), .B1(new_n396), .B2(new_n187), .ZN(new_n397));
  INV_X1    g211(.A(G469), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(new_n187), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n237), .A2(G227), .ZN(new_n400));
  XOR2_X1   g214(.A(G110), .B(G140), .Z(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n342), .A2(new_n345), .A3(new_n296), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n300), .A2(new_n301), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n340), .A2(new_n317), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n321), .B1(new_n405), .B2(new_n313), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n406), .A3(KEYINPUT10), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT84), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n406), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT10), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n404), .A2(new_n406), .A3(new_n412), .A4(KEYINPUT10), .ZN(new_n413));
  AND4_X1   g227(.A1(new_n403), .A2(new_n408), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G131), .ZN(new_n415));
  INV_X1    g229(.A(G134), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT11), .B1(new_n416), .B2(G137), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT11), .ZN(new_n418));
  INV_X1    g232(.A(G137), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(G134), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n419), .A2(G134), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n415), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n418), .B1(G134), .B2(new_n419), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n416), .A2(KEYINPUT11), .A3(G137), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n415), .B(new_n423), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n402), .B1(new_n414), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n408), .A2(new_n403), .A3(new_n411), .A4(new_n413), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n429), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n300), .A2(new_n301), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n312), .B1(new_n340), .B2(new_n317), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n321), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n409), .A2(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n437), .A2(KEYINPUT12), .A3(new_n429), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT12), .B1(new_n437), .B2(new_n429), .ZN(new_n439));
  OAI22_X1  g253(.A1(new_n432), .A2(new_n429), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n431), .A2(new_n433), .B1(new_n440), .B2(new_n402), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n399), .B1(new_n441), .B2(G469), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n432), .A2(new_n429), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n438), .A2(new_n439), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n443), .A2(new_n444), .A3(new_n402), .ZN(new_n445));
  INV_X1    g259(.A(new_n402), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n414), .A2(new_n430), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(new_n433), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n398), .B(new_n187), .C1(new_n445), .C2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n397), .B1(new_n442), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT68), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  INV_X1    g267(.A(G237), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n451), .A2(new_n453), .A3(G214), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n289), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n237), .A2(G143), .A3(G214), .A4(new_n454), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(new_n415), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT88), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n457), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G131), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n456), .A2(new_n457), .A3(new_n462), .A4(new_n415), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n207), .A2(KEYINPUT19), .A3(new_n208), .ZN(new_n466));
  XNOR2_X1  g280(.A(G125), .B(G140), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT19), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT89), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n207), .A2(KEYINPUT89), .A3(KEYINPUT19), .A4(new_n208), .ZN(new_n471));
  AOI21_X1  g285(.A(G146), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT90), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n213), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI211_X1 g288(.A(KEYINPUT90), .B(G146), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n465), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n207), .A2(G146), .A3(new_n208), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n228), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT18), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n456), .B(new_n457), .C1(new_n479), .C2(new_n415), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n479), .B(new_n415), .C1(new_n456), .C2(new_n457), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G113), .B(G122), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(new_n309), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n481), .A2(new_n482), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n459), .A2(new_n461), .A3(new_n489), .A4(new_n463), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n460), .A2(KEYINPUT17), .A3(G131), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n491), .A2(new_n213), .A3(new_n215), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI22_X1  g307(.A1(new_n476), .A2(new_n487), .B1(new_n493), .B2(new_n486), .ZN(new_n494));
  NOR2_X1   g308(.A1(G475), .A2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT20), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n474), .A2(new_n475), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n464), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n488), .A2(new_n485), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n490), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n491), .A2(new_n213), .A3(new_n215), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n483), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n485), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n501), .A2(new_n505), .A3(new_n506), .A4(new_n495), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n497), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n304), .A2(G952), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n240), .B2(new_n454), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n187), .B(new_n237), .C1(G234), .C2(G237), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT21), .B(G898), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n396), .A2(G217), .A3(new_n304), .ZN(new_n515));
  INV_X1    g329(.A(G122), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G116), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n350), .A2(G122), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT92), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT92), .ZN(new_n522));
  AOI21_X1  g336(.A(G107), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n188), .B2(G143), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n289), .A2(KEYINPUT93), .A3(G128), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(G128), .B2(new_n289), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G134), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n527), .B(new_n416), .C1(G128), .C2(new_n289), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n523), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n532));
  OAI21_X1  g346(.A(G107), .B1(new_n518), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n534), .B(KEYINPUT96), .C1(KEYINPUT14), .C2(new_n519), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT96), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n519), .A2(KEYINPUT14), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n536), .B1(new_n537), .B2(new_n533), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(KEYINPUT94), .A2(KEYINPUT13), .ZN(new_n540));
  NOR2_X1   g354(.A1(KEYINPUT94), .A2(KEYINPUT13), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n527), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n289), .A2(G128), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n527), .B2(new_n542), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI211_X1 g361(.A(KEYINPUT95), .B(new_n544), .C1(new_n527), .C2(new_n542), .ZN(new_n548));
  OAI21_X1  g362(.A(G134), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n530), .ZN(new_n550));
  INV_X1    g364(.A(new_n523), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n521), .A2(new_n522), .A3(G107), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI221_X4 g367(.A(new_n515), .B1(new_n531), .B2(new_n539), .C1(new_n549), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n515), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n549), .A2(new_n553), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n531), .A2(new_n539), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n187), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G478), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT97), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n561), .B(KEYINPUT97), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n187), .B(new_n566), .C1(new_n554), .C2(new_n558), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n514), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n485), .A2(KEYINPUT91), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n483), .B(new_n569), .C1(new_n502), .C2(new_n503), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n187), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n493), .A2(new_n569), .ZN(new_n572));
  OAI21_X1  g386(.A(G475), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n508), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  AND4_X1   g388(.A1(new_n285), .A2(new_n394), .A3(new_n450), .A4(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n237), .A2(G210), .A3(new_n454), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT27), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT27), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n237), .A2(new_n578), .A3(G210), .A4(new_n454), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT26), .B(G101), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n586));
  NAND2_X1  g400(.A1(new_n353), .A2(new_n331), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT67), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n353), .A2(new_n331), .A3(KEYINPUT67), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n428), .A2(new_n301), .A3(new_n300), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT64), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n419), .B2(G134), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n419), .A2(G134), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n416), .A2(KEYINPUT64), .A3(G137), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n597), .A2(KEYINPUT65), .A3(G131), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT65), .B1(new_n597), .B2(G131), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n592), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n295), .B1(new_n425), .B2(new_n428), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n591), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(G131), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT65), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n597), .A2(KEYINPUT65), .A3(G131), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n404), .A2(new_n605), .A3(new_n428), .A4(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n428), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n296), .B1(new_n608), .B2(new_n424), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n607), .A2(new_n609), .A3(new_n589), .A4(new_n590), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n586), .B1(new_n602), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n600), .A2(new_n601), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT28), .B1(new_n612), .B2(new_n356), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n585), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n607), .A2(KEYINPUT30), .A3(new_n609), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n591), .B(new_n615), .C1(new_n612), .C2(KEYINPUT30), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n585), .B1(new_n612), .B2(new_n356), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n609), .A2(KEYINPUT30), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n591), .B1(new_n621), .B2(new_n600), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT30), .B1(new_n607), .B2(new_n609), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n585), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n610), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT69), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT69), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n616), .A2(new_n628), .A3(new_n617), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(KEYINPUT31), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n620), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(G472), .A2(G902), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT72), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT32), .ZN(new_n635));
  INV_X1    g449(.A(new_n632), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n620), .B2(new_n630), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT72), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n634), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT28), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n602), .B2(new_n610), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT73), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n610), .A2(new_n641), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT73), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n644), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(KEYINPUT29), .A3(new_n625), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n611), .A2(new_n613), .A3(new_n585), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n616), .A2(new_n610), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n585), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT29), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n648), .B(new_n187), .C1(new_n649), .C2(new_n653), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n654), .A2(G472), .B1(new_n637), .B2(KEYINPUT32), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n640), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n284), .A2(new_n575), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G101), .ZN(G3));
  AND3_X1   g472(.A1(new_n627), .A2(KEYINPUT31), .A3(new_n629), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n614), .A2(new_n619), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n187), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G472), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n634), .A2(new_n450), .A3(new_n639), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n284), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT98), .ZN(new_n665));
  INV_X1    g479(.A(new_n514), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n371), .A2(new_n385), .A3(new_n287), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n286), .B1(new_n392), .B2(new_n384), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n285), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n508), .A2(new_n573), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n560), .A2(new_n187), .ZN(new_n671));
  INV_X1    g485(.A(new_n552), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n530), .B1(new_n672), .B2(new_n523), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n527), .A2(new_n542), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT95), .B1(new_n674), .B2(new_n544), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n545), .A2(new_n546), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n676), .A3(new_n543), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n673), .B1(new_n677), .B2(G134), .ZN(new_n678));
  INV_X1    g492(.A(new_n557), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n515), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n556), .A2(new_n557), .A3(new_n555), .ZN(new_n681));
  AOI21_X1  g495(.A(G902), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n671), .B1(new_n682), .B2(new_n560), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT33), .B1(new_n554), .B2(new_n558), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT33), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n680), .A2(new_n685), .A3(new_n681), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n684), .A2(new_n686), .A3(G478), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n670), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n669), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n665), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT34), .B(G104), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G6));
  OAI21_X1  g508(.A(new_n567), .B1(new_n682), .B2(new_n563), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n573), .A2(KEYINPUT99), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT99), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n698), .B(G475), .C1(new_n571), .C2(new_n572), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n508), .A2(new_n696), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n669), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n665), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT35), .B(G107), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G9));
  NAND2_X1  g518(.A1(new_n275), .A2(new_n277), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT82), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n275), .A2(KEYINPUT82), .A3(new_n277), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n264), .A2(KEYINPUT36), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n261), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n281), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n707), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n637), .A2(new_n638), .ZN(new_n713));
  INV_X1    g527(.A(G472), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n631), .B2(new_n187), .ZN(new_n715));
  AOI211_X1 g529(.A(KEYINPUT72), .B(new_n636), .C1(new_n620), .C2(new_n630), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n575), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT37), .B(G110), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT100), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n718), .B(new_n720), .ZN(G12));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT101), .B(G900), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n512), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n510), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n722), .B1(new_n700), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n697), .A2(new_n699), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n695), .B1(new_n497), .B2(new_n507), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(KEYINPUT102), .A3(new_n729), .A4(new_n725), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n394), .A2(new_n285), .A3(new_n450), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n731), .A2(new_n656), .A3(new_n733), .A4(new_n712), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G128), .ZN(G30));
  NOR3_X1   g549(.A1(new_n713), .A2(new_n716), .A3(KEYINPUT32), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n637), .A2(KEYINPUT32), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n627), .A2(new_n629), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n602), .A2(new_n610), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n585), .ZN(new_n740));
  AOI21_X1  g554(.A(G902), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n737), .B1(new_n741), .B2(new_n714), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT104), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n741), .A2(new_n714), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n640), .A2(new_n744), .A3(new_n737), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n394), .B(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n725), .B(KEYINPUT39), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n450), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT40), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n695), .B1(new_n508), .B2(new_n573), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n285), .B(new_n755), .C1(new_n752), .C2(KEYINPUT40), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n748), .A2(new_n754), .A3(new_n712), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n289), .ZN(G45));
  NAND3_X1  g572(.A1(new_n670), .A2(new_n689), .A3(new_n725), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n712), .A2(new_n733), .A3(new_n656), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G146), .ZN(G48));
  INV_X1    g576(.A(new_n433), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n402), .B1(new_n763), .B2(new_n443), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n447), .B(new_n446), .C1(new_n438), .C2(new_n439), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n187), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(G469), .ZN(new_n768));
  INV_X1    g582(.A(new_n397), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n769), .A3(new_n449), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n284), .A2(new_n691), .A3(new_n656), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT41), .B(G113), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G15));
  NAND4_X1  g588(.A1(new_n284), .A2(new_n701), .A3(new_n656), .A4(new_n771), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G116), .ZN(G18));
  OAI21_X1  g590(.A(new_n285), .B1(new_n667), .B2(new_n668), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n770), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n656), .A2(new_n712), .A3(new_n778), .A4(new_n574), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G119), .ZN(G21));
  INV_X1    g594(.A(KEYINPUT105), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n662), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n715), .A2(KEYINPUT105), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n630), .B(new_n619), .C1(new_n625), .C2(new_n647), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n782), .A2(new_n783), .B1(new_n632), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n394), .A2(new_n285), .A3(new_n755), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n770), .A2(new_n514), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n284), .A2(new_n785), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G122), .ZN(G24));
  NAND4_X1  g604(.A1(new_n785), .A2(new_n712), .A3(new_n778), .A4(new_n760), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G125), .ZN(G27));
  INV_X1    g606(.A(new_n450), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n386), .A2(new_n285), .A3(new_n393), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n284), .A2(new_n656), .A3(new_n760), .A4(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT42), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n654), .A2(G472), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n633), .A2(new_n635), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n737), .ZN(new_n800));
  INV_X1    g614(.A(new_n283), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n707), .A2(new_n800), .A3(new_n708), .A4(new_n801), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n793), .A2(new_n794), .A3(new_n759), .A4(new_n797), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n796), .A2(new_n797), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(new_n415), .ZN(G33));
  NAND4_X1  g619(.A1(new_n731), .A2(new_n284), .A3(new_n656), .A4(new_n795), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G134), .ZN(G36));
  INV_X1    g621(.A(KEYINPUT45), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n763), .A2(new_n443), .A3(new_n402), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n440), .A2(new_n402), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n441), .A2(KEYINPUT45), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(G469), .A3(new_n812), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT106), .Z(new_n814));
  INV_X1    g628(.A(new_n399), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(KEYINPUT46), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT107), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n815), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT46), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT107), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n814), .A2(new_n821), .A3(KEYINPUT46), .A4(new_n815), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n817), .A2(new_n820), .A3(new_n449), .A4(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n823), .A2(new_n769), .A3(new_n751), .ZN(new_n824));
  NAND2_X1  g638(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n825));
  XNOR2_X1  g639(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n670), .A2(new_n688), .ZN(new_n827));
  MUX2_X1   g641(.A(new_n825), .B(new_n826), .S(new_n827), .Z(new_n828));
  NOR2_X1   g642(.A1(new_n278), .A2(new_n279), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n717), .B1(new_n829), .B2(new_n711), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT44), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n794), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n828), .A2(new_n830), .A3(KEYINPUT44), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT109), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT109), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n833), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n824), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G137), .ZN(G39));
  NOR4_X1   g654(.A1(new_n284), .A2(new_n656), .A3(new_n759), .A4(new_n794), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n823), .A2(KEYINPUT47), .A3(new_n769), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT47), .B1(new_n823), .B2(new_n769), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(G140), .ZN(G42));
  NAND2_X1  g659(.A1(new_n768), .A2(new_n449), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n846), .A2(KEYINPUT49), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(KEYINPUT49), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n769), .A2(new_n285), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n847), .A2(new_n827), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n750), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n284), .A3(new_n748), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n770), .A2(new_n794), .A3(new_n510), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n748), .A2(new_n854), .A3(new_n284), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n855), .A2(new_n670), .A3(new_n689), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT117), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n284), .A2(new_n828), .A3(new_n511), .A4(new_n785), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n750), .A2(new_n285), .A3(new_n770), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(KEYINPUT50), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(KEYINPUT50), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n828), .A2(new_n712), .A3(new_n785), .A4(new_n854), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT116), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n857), .A2(new_n862), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n846), .A2(new_n769), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n842), .A2(new_n843), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n794), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n853), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n802), .A2(new_n828), .A3(new_n854), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT48), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n778), .B2(new_n859), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n874), .A2(KEYINPUT48), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n878), .A3(new_n875), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n879), .A2(new_n509), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n877), .B(new_n880), .C1(new_n690), .C2(new_n855), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT119), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n872), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n725), .B(KEYINPUT111), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n397), .B(new_n884), .C1(new_n442), .C2(new_n449), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n829), .A2(KEYINPUT112), .A3(new_n711), .A4(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n707), .A2(new_n885), .A3(new_n708), .A4(new_n711), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT112), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n747), .A2(new_n787), .A3(new_n886), .A4(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n734), .A2(new_n761), .A3(new_n791), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT52), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n785), .A2(new_n712), .A3(new_n760), .A4(new_n795), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n508), .A2(new_n728), .A3(new_n695), .A4(new_n725), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n712), .A2(new_n656), .A3(new_n795), .A4(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n806), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n669), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT110), .ZN(new_n898));
  INV_X1    g712(.A(new_n572), .ZN(new_n899));
  AOI21_X1  g713(.A(G902), .B1(new_n493), .B2(new_n569), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n497), .A2(new_n507), .B1(G475), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n898), .B1(new_n902), .B2(new_n688), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n670), .A2(KEYINPUT110), .A3(new_n689), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n903), .B(new_n904), .C1(new_n670), .C2(new_n695), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n284), .A2(new_n897), .A3(new_n663), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n657), .A3(new_n718), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n896), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n747), .A2(new_n886), .A3(new_n889), .A4(new_n787), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT52), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n732), .B1(new_n640), .B2(new_n655), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n912), .B(new_n712), .C1(new_n731), .C2(new_n760), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n910), .A2(new_n911), .A3(new_n791), .A4(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n772), .A2(new_n775), .A3(new_n789), .A4(new_n779), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n804), .ZN(new_n916));
  AND4_X1   g730(.A1(new_n892), .A2(new_n909), .A3(new_n914), .A4(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT114), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n896), .A2(new_n907), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n892), .A2(new_n914), .A3(new_n916), .A4(new_n919), .ZN(new_n920));
  XOR2_X1   g734(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n921));
  AOI22_X1  g735(.A1(new_n917), .A2(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n892), .A2(new_n914), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n909), .A2(new_n916), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT114), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n920), .A2(new_n908), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n920), .B2(new_n921), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT54), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n866), .A2(new_n871), .A3(new_n853), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n883), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(G952), .A2(G953), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n852), .B1(new_n933), .B2(new_n934), .ZN(G75));
  NOR2_X1   g749(.A1(new_n391), .A2(new_n306), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n371), .ZN(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n796), .A2(new_n797), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n802), .A2(new_n803), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n772), .A2(new_n789), .A3(new_n779), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n943), .A3(new_n775), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n806), .A2(new_n893), .A3(new_n895), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n906), .A2(new_n657), .A3(new_n718), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT53), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n948), .A2(new_n918), .A3(new_n892), .A4(new_n914), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n920), .A2(new_n921), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n949), .A2(new_n926), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(G902), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(G210), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT56), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT121), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n955), .A2(KEYINPUT121), .ZN(new_n957));
  AND4_X1   g771(.A1(new_n939), .A2(new_n954), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n939), .B1(new_n954), .B2(new_n955), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n237), .A2(G952), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(G51));
  NOR2_X1   g775(.A1(new_n952), .A2(new_n814), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n399), .B(KEYINPUT57), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n923), .B1(new_n922), .B2(new_n926), .ZN(new_n964));
  AND4_X1   g778(.A1(new_n923), .A2(new_n949), .A3(new_n926), .A4(new_n950), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n962), .B1(new_n966), .B2(new_n766), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT122), .B1(new_n967), .B2(new_n960), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT122), .ZN(new_n969));
  INV_X1    g783(.A(new_n960), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n951), .A2(KEYINPUT54), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n927), .ZN(new_n972));
  AOI22_X1  g786(.A1(new_n972), .A2(new_n963), .B1(new_n764), .B2(new_n765), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n969), .B(new_n970), .C1(new_n973), .C2(new_n962), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n968), .A2(new_n974), .ZN(G54));
  NAND3_X1  g789(.A1(new_n953), .A2(KEYINPUT58), .A3(G475), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n976), .A2(new_n494), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n494), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n977), .A2(new_n978), .A3(new_n960), .ZN(G60));
  NAND2_X1  g793(.A1(new_n684), .A2(new_n686), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n671), .B(KEYINPUT59), .Z(new_n981));
  AND3_X1   g795(.A1(new_n972), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n931), .B2(new_n981), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n982), .A2(new_n983), .A3(new_n960), .ZN(G63));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT60), .Z(new_n986));
  NAND2_X1  g800(.A1(new_n951), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n280), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n951), .A2(new_n710), .A3(new_n986), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT61), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n960), .B1(KEYINPUT123), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n990), .A2(KEYINPUT123), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n992), .B(new_n993), .Z(G66));
  INV_X1    g808(.A(G224), .ZN(new_n995));
  OAI21_X1  g809(.A(G953), .B1(new_n513), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n915), .A2(new_n907), .ZN(new_n997));
  INV_X1    g811(.A(new_n237), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n364), .B(new_n370), .C1(G898), .C2(new_n237), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT124), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n999), .B(new_n1001), .ZN(G69));
  AND2_X1   g816(.A1(new_n905), .A2(new_n751), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n1003), .A2(new_n656), .A3(new_n284), .A4(new_n795), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n839), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(KEYINPUT125), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  OR3_X1    g821(.A1(new_n757), .A2(new_n1007), .A3(new_n891), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1007), .B1(new_n757), .B2(new_n891), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1010), .A2(new_n844), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT125), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n839), .A2(new_n1012), .A3(new_n1004), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1006), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n237), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n615), .B1(new_n612), .B2(KEYINPUT30), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n470), .A2(new_n471), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G227), .A2(G900), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n998), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT126), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n942), .A2(new_n791), .A3(new_n806), .A4(new_n913), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n802), .A2(new_n787), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n824), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n844), .A2(new_n1026), .A3(new_n839), .ZN(new_n1027));
  OR2_X1    g841(.A1(new_n1027), .A2(new_n998), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1018), .B1(G900), .B2(new_n998), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1019), .A2(new_n1023), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1023), .B1(new_n1019), .B2(new_n1030), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1031), .A2(new_n1032), .ZN(G72));
  NAND2_X1  g847(.A1(new_n650), .A2(new_n625), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1006), .A2(new_n1011), .A3(new_n997), .A4(new_n1013), .ZN(new_n1035));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  AOI21_X1  g851(.A(new_n1034), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n997), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1037), .B1(new_n1027), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n616), .A2(new_n610), .A3(new_n585), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1037), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1044), .B1(new_n738), .B2(new_n651), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n960), .B1(new_n929), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1038), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(KEYINPUT127), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g864(.A(KEYINPUT127), .B1(new_n1038), .B2(new_n1047), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(G57));
endmodule


