

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745;

  XNOR2_X1 U372 ( .A(n581), .B(n580), .ZN(n607) );
  INV_X1 U373 ( .A(n671), .ZN(n593) );
  NOR2_X1 U374 ( .A1(G953), .A2(G237), .ZN(n504) );
  NOR2_X1 U375 ( .A1(n578), .A2(n577), .ZN(n581) );
  XNOR2_X1 U376 ( .A(n357), .B(n476), .ZN(n442) );
  INV_X1 U377 ( .A(G953), .ZN(n449) );
  BUF_X1 U378 ( .A(n645), .Z(n352) );
  XNOR2_X2 U379 ( .A(n372), .B(n719), .ZN(n626) );
  XNOR2_X2 U380 ( .A(KEYINPUT33), .B(n594), .ZN(n668) );
  XNOR2_X2 U381 ( .A(n727), .B(n463), .ZN(n476) );
  XNOR2_X1 U382 ( .A(n353), .B(n562), .ZN(n563) );
  INV_X1 U383 ( .A(n591), .ZN(n587) );
  XNOR2_X1 U384 ( .A(G902), .B(KEYINPUT15), .ZN(n623) );
  INV_X1 U385 ( .A(KEYINPUT4), .ZN(n422) );
  NOR2_X1 U386 ( .A1(n354), .A2(n430), .ZN(n374) );
  OR2_X1 U387 ( .A1(n742), .A2(n640), .ZN(n621) );
  XNOR2_X1 U388 ( .A(n416), .B(n415), .ZN(n742) );
  NOR2_X1 U389 ( .A1(n563), .A2(n671), .ZN(n564) );
  NOR2_X1 U390 ( .A1(n587), .A2(n369), .ZN(n528) );
  NAND2_X1 U391 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U392 ( .A(n499), .B(n498), .Z(n719) );
  XNOR2_X1 U393 ( .A(n521), .B(n440), .ZN(n727) );
  XNOR2_X1 U394 ( .A(n422), .B(KEYINPUT66), .ZN(n489) );
  INV_X1 U395 ( .A(n623), .ZN(n376) );
  AND2_X4 U396 ( .A1(n377), .A2(n376), .ZN(n417) );
  BUF_X2 U397 ( .A(n417), .Z(n350) );
  INV_X1 U398 ( .A(n587), .ZN(n351) );
  XNOR2_X1 U399 ( .A(n608), .B(KEYINPUT6), .ZN(n591) );
  XNOR2_X1 U400 ( .A(n396), .B(n520), .ZN(n704) );
  NOR2_X2 U401 ( .A1(G902), .A2(n442), .ZN(n443) );
  XNOR2_X1 U402 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U403 ( .A(KEYINPUT18), .B(KEYINPUT86), .Z(n491) );
  XNOR2_X1 U404 ( .A(n381), .B(KEYINPUT68), .ZN(n533) );
  XNOR2_X1 U405 ( .A(n511), .B(n726), .ZN(n701) );
  INV_X1 U406 ( .A(n486), .ZN(n412) );
  XOR2_X1 U407 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n454) );
  INV_X1 U408 ( .A(G137), .ZN(n439) );
  NAND2_X1 U409 ( .A1(n601), .A2(n600), .ZN(n430) );
  NOR2_X1 U410 ( .A1(G237), .A2(G902), .ZN(n441) );
  INV_X1 U411 ( .A(n533), .ZN(n370) );
  NAND2_X1 U412 ( .A1(n582), .A2(n659), .ZN(n665) );
  XNOR2_X1 U413 ( .A(n560), .B(n386), .ZN(n662) );
  INV_X1 U414 ( .A(KEYINPUT38), .ZN(n386) );
  XNOR2_X1 U415 ( .A(n522), .B(G478), .ZN(n555) );
  NOR2_X1 U416 ( .A1(n704), .A2(G902), .ZN(n522) );
  INV_X1 U417 ( .A(n670), .ZN(n604) );
  XNOR2_X1 U418 ( .A(n586), .B(n585), .ZN(n590) );
  INV_X1 U419 ( .A(KEYINPUT71), .ZN(n584) );
  XNOR2_X1 U420 ( .A(n393), .B(n435), .ZN(n497) );
  XNOR2_X1 U421 ( .A(n434), .B(G119), .ZN(n393) );
  INV_X1 U422 ( .A(G104), .ZN(n478) );
  INV_X1 U423 ( .A(KEYINPUT8), .ZN(n390) );
  XNOR2_X1 U424 ( .A(n535), .B(n379), .ZN(n671) );
  INV_X1 U425 ( .A(KEYINPUT1), .ZN(n379) );
  XNOR2_X1 U426 ( .A(n513), .B(n420), .ZN(n556) );
  XNOR2_X1 U427 ( .A(n512), .B(G475), .ZN(n420) );
  INV_X1 U428 ( .A(n555), .ZN(n525) );
  XNOR2_X1 U429 ( .A(KEYINPUT94), .B(G472), .ZN(n432) );
  XNOR2_X1 U430 ( .A(n473), .B(n468), .ZN(n401) );
  NAND2_X1 U431 ( .A1(n657), .A2(n409), .ZN(n408) );
  NOR2_X1 U432 ( .A1(n693), .A2(n359), .ZN(n409) );
  INV_X1 U433 ( .A(KEYINPUT118), .ZN(n407) );
  XNOR2_X1 U434 ( .A(n544), .B(n368), .ZN(n658) );
  INV_X1 U435 ( .A(KEYINPUT99), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n419), .B(KEYINPUT101), .ZN(n660) );
  AND2_X1 U437 ( .A1(n555), .A2(n556), .ZN(n419) );
  XOR2_X1 U438 ( .A(G131), .B(G140), .Z(n509) );
  XNOR2_X1 U439 ( .A(n411), .B(n410), .ZN(n496) );
  XNOR2_X1 U440 ( .A(n487), .B(n488), .ZN(n410) );
  XNOR2_X1 U441 ( .A(n412), .B(n489), .ZN(n411) );
  XOR2_X1 U442 ( .A(KEYINPUT17), .B(KEYINPUT87), .Z(n488) );
  NAND2_X1 U443 ( .A1(n466), .A2(n465), .ZN(n486) );
  XOR2_X1 U444 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n506) );
  XOR2_X1 U445 ( .A(G143), .B(G104), .Z(n503) );
  XNOR2_X1 U446 ( .A(G113), .B(G122), .ZN(n502) );
  XNOR2_X1 U447 ( .A(n510), .B(n509), .ZN(n726) );
  OR2_X1 U448 ( .A1(n694), .A2(G902), .ZN(n367) );
  XNOR2_X1 U449 ( .A(n472), .B(n471), .ZN(n473) );
  INV_X1 U450 ( .A(n743), .ZN(n426) );
  XNOR2_X1 U451 ( .A(KEYINPUT16), .B(G122), .ZN(n499) );
  XNOR2_X1 U452 ( .A(n486), .B(n421), .ZN(n510) );
  INV_X1 U453 ( .A(KEYINPUT10), .ZN(n421) );
  INV_X1 U454 ( .A(n684), .ZN(n656) );
  NAND2_X1 U455 ( .A1(n647), .A2(n370), .ZN(n369) );
  XNOR2_X1 U456 ( .A(n418), .B(n538), .ZN(n684) );
  NOR2_X1 U457 ( .A1(n665), .A2(n662), .ZN(n418) );
  AND2_X1 U458 ( .A1(n680), .A2(n605), .ZN(n682) );
  INV_X1 U459 ( .A(n532), .ZN(n560) );
  INV_X1 U460 ( .A(KEYINPUT19), .ZN(n403) );
  NOR2_X1 U461 ( .A1(n590), .A2(n593), .ZN(n602) );
  XOR2_X1 U462 ( .A(G131), .B(KEYINPUT5), .Z(n437) );
  BUF_X1 U463 ( .A(n490), .Z(n733) );
  NAND2_X1 U464 ( .A1(n479), .A2(n480), .ZN(n481) );
  XNOR2_X1 U465 ( .A(n521), .B(n371), .ZN(n396) );
  INV_X1 U466 ( .A(KEYINPUT40), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n425), .B(n595), .ZN(n424) );
  XNOR2_X1 U468 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n415) );
  NAND2_X1 U469 ( .A1(n392), .A2(n589), .ZN(n416) );
  AND2_X1 U470 ( .A1(n602), .A2(n413), .ZN(n640) );
  NOR2_X1 U471 ( .A1(n674), .A2(n680), .ZN(n413) );
  XOR2_X1 U472 ( .A(n523), .B(KEYINPUT98), .Z(n651) );
  INV_X1 U473 ( .A(KEYINPUT60), .ZN(n384) );
  INV_X1 U474 ( .A(KEYINPUT53), .ZN(n394) );
  NAND2_X1 U475 ( .A1(n406), .A2(n713), .ZN(n395) );
  XNOR2_X1 U476 ( .A(n408), .B(n407), .ZN(n406) );
  OR2_X1 U477 ( .A1(n561), .A2(n560), .ZN(n353) );
  AND2_X1 U478 ( .A1(n622), .A2(n621), .ZN(n354) );
  XNOR2_X1 U479 ( .A(n557), .B(KEYINPUT102), .ZN(n355) );
  XOR2_X1 U480 ( .A(KEYINPUT69), .B(G469), .Z(n356) );
  XNOR2_X1 U481 ( .A(n497), .B(n438), .ZN(n357) );
  XOR2_X1 U482 ( .A(n618), .B(n617), .Z(n358) );
  NOR2_X1 U483 ( .A1(n525), .A2(n556), .ZN(n647) );
  AND2_X1 U484 ( .A1(n668), .A2(n656), .ZN(n359) );
  XOR2_X1 U485 ( .A(n442), .B(KEYINPUT62), .Z(n360) );
  XOR2_X1 U486 ( .A(n701), .B(n700), .Z(n361) );
  XNOR2_X1 U487 ( .A(n628), .B(n627), .ZN(n362) );
  NOR2_X1 U488 ( .A1(n733), .A2(G952), .ZN(n711) );
  INV_X1 U489 ( .A(n711), .ZN(n387) );
  XOR2_X1 U490 ( .A(n630), .B(KEYINPUT79), .Z(n363) );
  AND2_X1 U491 ( .A1(n552), .A2(n551), .ZN(n567) );
  NAND2_X1 U492 ( .A1(n365), .A2(n364), .ZN(n372) );
  NAND2_X1 U493 ( .A1(n495), .A2(n496), .ZN(n364) );
  NAND2_X1 U494 ( .A1(n400), .A2(n399), .ZN(n365) );
  NOR2_X1 U495 ( .A1(n366), .A2(n358), .ZN(n373) );
  NAND2_X1 U496 ( .A1(n380), .A2(n616), .ZN(n366) );
  XNOR2_X2 U497 ( .A(n367), .B(n356), .ZN(n535) );
  INV_X1 U498 ( .A(n658), .ZN(n612) );
  NAND2_X1 U499 ( .A1(n658), .A2(n352), .ZN(n545) );
  NAND2_X1 U500 ( .A1(n519), .A2(G217), .ZN(n371) );
  NAND2_X1 U501 ( .A1(n374), .A2(n373), .ZN(n429) );
  NAND2_X2 U502 ( .A1(n732), .A2(n712), .ZN(n654) );
  XNOR2_X2 U503 ( .A(n654), .B(KEYINPUT2), .ZN(n377) );
  XNOR2_X1 U504 ( .A(n375), .B(n363), .ZN(G51) );
  NAND2_X1 U505 ( .A1(n378), .A2(n387), .ZN(n375) );
  INV_X1 U506 ( .A(n496), .ZN(n399) );
  XNOR2_X1 U507 ( .A(n629), .B(n362), .ZN(n378) );
  NOR2_X1 U508 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U509 ( .A(n404), .B(n403), .ZN(n578) );
  INV_X1 U510 ( .A(n495), .ZN(n400) );
  NAND2_X1 U511 ( .A1(n615), .A2(KEYINPUT65), .ZN(n380) );
  NAND2_X1 U512 ( .A1(n527), .A2(n673), .ZN(n381) );
  XNOR2_X1 U513 ( .A(n462), .B(n382), .ZN(n467) );
  XNOR2_X1 U514 ( .A(n460), .B(n383), .ZN(n382) );
  INV_X1 U515 ( .A(n461), .ZN(n383) );
  INV_X1 U516 ( .A(n590), .ZN(n392) );
  XNOR2_X1 U517 ( .A(n385), .B(n384), .ZN(G60) );
  NAND2_X1 U518 ( .A1(n388), .A2(n387), .ZN(n385) );
  NAND2_X1 U519 ( .A1(n626), .A2(n623), .ZN(n405) );
  NAND2_X1 U520 ( .A1(n424), .A2(n355), .ZN(n423) );
  XNOR2_X1 U521 ( .A(n483), .B(n475), .ZN(n402) );
  XNOR2_X1 U522 ( .A(n476), .B(n402), .ZN(n694) );
  NAND2_X1 U523 ( .A1(n485), .A2(n484), .ZN(n553) );
  NOR2_X2 U524 ( .A1(n741), .A2(n744), .ZN(n389) );
  XNOR2_X1 U525 ( .A(n702), .B(n361), .ZN(n388) );
  OR2_X2 U526 ( .A1(n540), .A2(n543), .ZN(n398) );
  XNOR2_X1 U527 ( .A(n389), .B(KEYINPUT46), .ZN(n552) );
  NOR2_X2 U528 ( .A1(n553), .A2(n662), .ZN(n501) );
  XNOR2_X2 U529 ( .A(n391), .B(n390), .ZN(n519) );
  NAND2_X1 U530 ( .A1(n490), .A2(G234), .ZN(n391) );
  INV_X1 U531 ( .A(n608), .ZN(n414) );
  XNOR2_X1 U532 ( .A(n395), .B(n394), .ZN(G75) );
  XNOR2_X2 U533 ( .A(n398), .B(n397), .ZN(n741) );
  NOR2_X1 U534 ( .A1(n684), .A2(n541), .ZN(n539) );
  XNOR2_X2 U535 ( .A(n405), .B(n433), .ZN(n532) );
  XNOR2_X1 U536 ( .A(n467), .B(n510), .ZN(n707) );
  XNOR2_X2 U537 ( .A(n469), .B(n401), .ZN(n674) );
  XNOR2_X2 U538 ( .A(n429), .B(KEYINPUT45), .ZN(n712) );
  NAND2_X1 U539 ( .A1(n532), .A2(n659), .ZN(n404) );
  XNOR2_X2 U540 ( .A(n720), .B(KEYINPUT70), .ZN(n494) );
  XNOR2_X2 U541 ( .A(n481), .B(G107), .ZN(n720) );
  NAND2_X1 U542 ( .A1(n417), .A2(G475), .ZN(n702) );
  NAND2_X1 U543 ( .A1(n417), .A2(G210), .ZN(n629) );
  NAND2_X1 U544 ( .A1(n417), .A2(G472), .ZN(n431) );
  NAND2_X1 U545 ( .A1(n417), .A2(G478), .ZN(n703) );
  NAND2_X1 U546 ( .A1(n350), .A2(G469), .ZN(n697) );
  NAND2_X1 U547 ( .A1(n350), .A2(G217), .ZN(n709) );
  XNOR2_X2 U548 ( .A(n423), .B(KEYINPUT35), .ZN(n739) );
  NAND2_X1 U549 ( .A1(n668), .A2(n607), .ZN(n425) );
  AND2_X2 U550 ( .A1(n427), .A2(n426), .ZN(n732) );
  XNOR2_X1 U551 ( .A(n428), .B(KEYINPUT78), .ZN(n427) );
  NOR2_X2 U552 ( .A1(n571), .A2(n653), .ZN(n428) );
  XNOR2_X1 U553 ( .A(n431), .B(n360), .ZN(n624) );
  XNOR2_X2 U554 ( .A(n443), .B(n432), .ZN(n608) );
  AND2_X1 U555 ( .A1(n500), .A2(G210), .ZN(n433) );
  INV_X1 U556 ( .A(n733), .ZN(n450) );
  INV_X1 U557 ( .A(KEYINPUT81), .ZN(n617) );
  XNOR2_X1 U558 ( .A(n568), .B(KEYINPUT67), .ZN(n569) );
  INV_X1 U559 ( .A(KEYINPUT30), .ZN(n444) );
  XNOR2_X1 U560 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U561 ( .A(n474), .B(KEYINPUT74), .ZN(n475) );
  XNOR2_X1 U562 ( .A(n445), .B(n444), .ZN(n485) );
  XNOR2_X1 U563 ( .A(n494), .B(n482), .ZN(n483) );
  XNOR2_X1 U564 ( .A(n584), .B(KEYINPUT22), .ZN(n585) );
  XNOR2_X1 U565 ( .A(n579), .B(KEYINPUT85), .ZN(n580) );
  AND2_X1 U566 ( .A1(n588), .A2(n593), .ZN(n589) );
  INV_X1 U567 ( .A(KEYINPUT92), .ZN(n471) );
  INV_X1 U568 ( .A(KEYINPUT121), .ZN(n706) );
  NAND2_X1 U569 ( .A1(n624), .A2(n387), .ZN(n625) );
  XNOR2_X1 U570 ( .A(n709), .B(n708), .ZN(n710) );
  XOR2_X1 U571 ( .A(KEYINPUT3), .B(G116), .Z(n435) );
  XNOR2_X1 U572 ( .A(G113), .B(G101), .ZN(n434) );
  NAND2_X1 U573 ( .A1(n504), .A2(G210), .ZN(n436) );
  XNOR2_X1 U574 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X2 U575 ( .A(G143), .B(G128), .Z(n487) );
  XNOR2_X2 U576 ( .A(n487), .B(G134), .ZN(n521) );
  XNOR2_X1 U577 ( .A(n489), .B(n439), .ZN(n440) );
  XOR2_X1 U578 ( .A(KEYINPUT72), .B(n441), .Z(n500) );
  NAND2_X1 U579 ( .A1(n500), .A2(G214), .ZN(n659) );
  INV_X1 U580 ( .A(n608), .ZN(n680) );
  NAND2_X1 U581 ( .A1(n659), .A2(n414), .ZN(n445) );
  NAND2_X1 U582 ( .A1(G234), .A2(G237), .ZN(n446) );
  XNOR2_X1 U583 ( .A(n446), .B(KEYINPUT14), .ZN(n447) );
  NAND2_X1 U584 ( .A1(n447), .A2(G952), .ZN(n691) );
  NOR2_X1 U585 ( .A1(G953), .A2(n691), .ZN(n575) );
  NAND2_X1 U586 ( .A1(n447), .A2(G902), .ZN(n448) );
  XOR2_X1 U587 ( .A(KEYINPUT88), .B(n448), .Z(n572) );
  XNOR2_X2 U588 ( .A(n449), .B(KEYINPUT64), .ZN(n490) );
  NAND2_X1 U589 ( .A1(n572), .A2(n450), .ZN(n451) );
  NOR2_X1 U590 ( .A1(G900), .A2(n451), .ZN(n452) );
  NOR2_X1 U591 ( .A1(n575), .A2(n452), .ZN(n526) );
  NAND2_X1 U592 ( .A1(G234), .A2(n623), .ZN(n453) );
  XNOR2_X1 U593 ( .A(n454), .B(n453), .ZN(n470) );
  NAND2_X1 U594 ( .A1(n470), .A2(G221), .ZN(n455) );
  XOR2_X1 U595 ( .A(KEYINPUT21), .B(n455), .Z(n456) );
  XOR2_X1 U596 ( .A(KEYINPUT93), .B(n456), .Z(n673) );
  XNOR2_X1 U597 ( .A(G119), .B(G137), .ZN(n457) );
  XNOR2_X1 U598 ( .A(n457), .B(KEYINPUT23), .ZN(n461) );
  XOR2_X1 U599 ( .A(KEYINPUT24), .B(G140), .Z(n459) );
  XNOR2_X1 U600 ( .A(G110), .B(G128), .ZN(n458) );
  XNOR2_X1 U601 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U602 ( .A1(G221), .A2(n519), .ZN(n462) );
  INV_X1 U603 ( .A(G146), .ZN(n463) );
  NAND2_X1 U604 ( .A1(G125), .A2(n463), .ZN(n466) );
  INV_X1 U605 ( .A(G125), .ZN(n464) );
  NAND2_X1 U606 ( .A1(n464), .A2(G146), .ZN(n465) );
  NOR2_X1 U607 ( .A1(n707), .A2(G902), .ZN(n469) );
  XNOR2_X1 U608 ( .A(KEYINPUT25), .B(KEYINPUT73), .ZN(n468) );
  NAND2_X1 U609 ( .A1(n470), .A2(G217), .ZN(n472) );
  NAND2_X1 U610 ( .A1(n673), .A2(n674), .ZN(n670) );
  XOR2_X1 U611 ( .A(G101), .B(n509), .Z(n474) );
  INV_X1 U612 ( .A(G110), .ZN(n477) );
  NAND2_X1 U613 ( .A1(n477), .A2(G104), .ZN(n480) );
  NAND2_X1 U614 ( .A1(n478), .A2(G110), .ZN(n479) );
  NAND2_X1 U615 ( .A1(G227), .A2(n733), .ZN(n482) );
  NAND2_X1 U616 ( .A1(n604), .A2(n535), .ZN(n610) );
  NOR2_X1 U617 ( .A1(n526), .A2(n610), .ZN(n484) );
  NAND2_X1 U618 ( .A1(G224), .A2(n490), .ZN(n492) );
  XNOR2_X1 U619 ( .A(n492), .B(n491), .ZN(n493) );
  INV_X1 U620 ( .A(n497), .ZN(n498) );
  XNOR2_X1 U621 ( .A(n501), .B(KEYINPUT39), .ZN(n540) );
  XNOR2_X1 U622 ( .A(n503), .B(n502), .ZN(n508) );
  NAND2_X1 U623 ( .A1(n504), .A2(G214), .ZN(n505) );
  XNOR2_X1 U624 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U625 ( .A(n508), .B(n507), .ZN(n511) );
  NOR2_X1 U626 ( .A1(G902), .A2(n701), .ZN(n513) );
  XNOR2_X1 U627 ( .A(KEYINPUT13), .B(KEYINPUT95), .ZN(n512) );
  XNOR2_X1 U628 ( .A(G116), .B(G122), .ZN(n514) );
  XNOR2_X1 U629 ( .A(n514), .B(KEYINPUT97), .ZN(n518) );
  XOR2_X1 U630 ( .A(KEYINPUT96), .B(KEYINPUT7), .Z(n516) );
  XNOR2_X1 U631 ( .A(G107), .B(KEYINPUT9), .ZN(n515) );
  XNOR2_X1 U632 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U633 ( .A(n518), .B(n517), .Z(n520) );
  NAND2_X1 U634 ( .A1(n556), .A2(n525), .ZN(n523) );
  INV_X1 U635 ( .A(n651), .ZN(n542) );
  NOR2_X1 U636 ( .A1(n540), .A2(n542), .ZN(n524) );
  XNOR2_X1 U637 ( .A(n524), .B(KEYINPUT108), .ZN(n743) );
  INV_X1 U638 ( .A(n647), .ZN(n543) );
  NOR2_X1 U639 ( .A1(n674), .A2(n526), .ZN(n527) );
  NAND2_X1 U640 ( .A1(n528), .A2(n659), .ZN(n561) );
  NOR2_X1 U641 ( .A1(n561), .A2(n593), .ZN(n529) );
  XNOR2_X1 U642 ( .A(n529), .B(KEYINPUT43), .ZN(n530) );
  XOR2_X1 U643 ( .A(KEYINPUT103), .B(n530), .Z(n531) );
  NOR2_X1 U644 ( .A1(n532), .A2(n531), .ZN(n653) );
  NOR2_X1 U645 ( .A1(n608), .A2(n533), .ZN(n534) );
  XNOR2_X1 U646 ( .A(KEYINPUT28), .B(n534), .ZN(n536) );
  NAND2_X1 U647 ( .A1(n536), .A2(n535), .ZN(n541) );
  INV_X1 U648 ( .A(n660), .ZN(n582) );
  XOR2_X1 U649 ( .A(KEYINPUT106), .B(KEYINPUT41), .Z(n537) );
  XNOR2_X1 U650 ( .A(KEYINPUT105), .B(n537), .ZN(n538) );
  XNOR2_X1 U651 ( .A(n539), .B(KEYINPUT42), .ZN(n744) );
  NOR2_X1 U652 ( .A1(n541), .A2(n578), .ZN(n645) );
  NAND2_X1 U653 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U654 ( .A(n545), .B(KEYINPUT47), .ZN(n547) );
  INV_X1 U655 ( .A(KEYINPUT77), .ZN(n546) );
  NAND2_X1 U656 ( .A1(n547), .A2(n546), .ZN(n550) );
  NAND2_X1 U657 ( .A1(KEYINPUT47), .A2(n658), .ZN(n548) );
  NAND2_X1 U658 ( .A1(n548), .A2(KEYINPUT77), .ZN(n549) );
  AND2_X1 U659 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U660 ( .A1(n560), .A2(n553), .ZN(n554) );
  XNOR2_X1 U661 ( .A(n554), .B(KEYINPUT104), .ZN(n558) );
  NOR2_X1 U662 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U663 ( .A1(n558), .A2(n355), .ZN(n644) );
  NAND2_X1 U664 ( .A1(n352), .A2(KEYINPUT77), .ZN(n559) );
  NAND2_X1 U665 ( .A1(n644), .A2(n559), .ZN(n565) );
  XOR2_X1 U666 ( .A(KEYINPUT36), .B(KEYINPUT83), .Z(n562) );
  XOR2_X1 U667 ( .A(KEYINPUT107), .B(n564), .Z(n737) );
  NOR2_X1 U668 ( .A1(n565), .A2(n737), .ZN(n566) );
  NAND2_X1 U669 ( .A1(n567), .A2(n566), .ZN(n570) );
  XOR2_X1 U670 ( .A(KEYINPUT80), .B(KEYINPUT48), .Z(n568) );
  INV_X1 U671 ( .A(G953), .ZN(n713) );
  NOR2_X1 U672 ( .A1(G898), .A2(n713), .ZN(n723) );
  NAND2_X1 U673 ( .A1(n723), .A2(n572), .ZN(n573) );
  XNOR2_X1 U674 ( .A(KEYINPUT89), .B(n573), .ZN(n574) );
  NOR2_X1 U675 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U676 ( .A(n576), .B(KEYINPUT90), .ZN(n577) );
  INV_X1 U677 ( .A(KEYINPUT0), .ZN(n579) );
  AND2_X1 U678 ( .A1(n673), .A2(n582), .ZN(n583) );
  NAND2_X1 U679 ( .A1(n607), .A2(n583), .ZN(n586) );
  NOR2_X1 U680 ( .A1(n591), .A2(n674), .ZN(n588) );
  INV_X1 U681 ( .A(KEYINPUT34), .ZN(n595) );
  AND2_X1 U682 ( .A1(n604), .A2(n591), .ZN(n592) );
  NOR2_X1 U683 ( .A1(n621), .A2(n739), .ZN(n598) );
  INV_X1 U684 ( .A(KEYINPUT44), .ZN(n596) );
  AND2_X1 U685 ( .A1(KEYINPUT82), .A2(n596), .ZN(n597) );
  NAND2_X1 U686 ( .A1(n598), .A2(n597), .ZN(n601) );
  INV_X1 U687 ( .A(KEYINPUT65), .ZN(n599) );
  OR2_X1 U688 ( .A1(KEYINPUT44), .A2(n599), .ZN(n600) );
  NAND2_X1 U689 ( .A1(n674), .A2(n602), .ZN(n603) );
  NOR2_X1 U690 ( .A1(n351), .A2(n603), .ZN(n631) );
  AND2_X1 U691 ( .A1(n604), .A2(n593), .ZN(n605) );
  NAND2_X1 U692 ( .A1(n607), .A2(n682), .ZN(n606) );
  XNOR2_X1 U693 ( .A(n606), .B(KEYINPUT31), .ZN(n650) );
  NAND2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U695 ( .A1(n610), .A2(n609), .ZN(n637) );
  NOR2_X1 U696 ( .A1(n650), .A2(n637), .ZN(n611) );
  XNOR2_X1 U697 ( .A(n613), .B(KEYINPUT100), .ZN(n614) );
  NOR2_X1 U698 ( .A1(n631), .A2(n614), .ZN(n616) );
  INV_X1 U699 ( .A(n621), .ZN(n615) );
  NAND2_X1 U700 ( .A1(n739), .A2(KEYINPUT44), .ZN(n618) );
  NOR2_X1 U701 ( .A1(n739), .A2(KEYINPUT82), .ZN(n619) );
  NOR2_X1 U702 ( .A1(KEYINPUT44), .A2(n619), .ZN(n620) );
  NOR2_X1 U703 ( .A1(KEYINPUT65), .A2(n620), .ZN(n622) );
  XNOR2_X1 U704 ( .A(n625), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U705 ( .A(KEYINPUT84), .B(KEYINPUT55), .Z(n628) );
  XNOR2_X1 U706 ( .A(n626), .B(KEYINPUT54), .ZN(n627) );
  INV_X1 U707 ( .A(KEYINPUT56), .ZN(n630) );
  XNOR2_X1 U708 ( .A(G101), .B(n631), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT109), .ZN(G3) );
  NAND2_X1 U710 ( .A1(n637), .A2(n647), .ZN(n633) );
  XNOR2_X1 U711 ( .A(n633), .B(G104), .ZN(G6) );
  XOR2_X1 U712 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n635) );
  XNOR2_X1 U713 ( .A(G107), .B(KEYINPUT110), .ZN(n634) );
  XNOR2_X1 U714 ( .A(n635), .B(n634), .ZN(n636) );
  XOR2_X1 U715 ( .A(KEYINPUT26), .B(n636), .Z(n639) );
  NAND2_X1 U716 ( .A1(n637), .A2(n651), .ZN(n638) );
  XNOR2_X1 U717 ( .A(n639), .B(n638), .ZN(G9) );
  XOR2_X1 U718 ( .A(G110), .B(n640), .Z(G12) );
  XOR2_X1 U719 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n642) );
  NAND2_X1 U720 ( .A1(n352), .A2(n651), .ZN(n641) );
  XNOR2_X1 U721 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U722 ( .A(G128), .B(n643), .ZN(G30) );
  XNOR2_X1 U723 ( .A(G143), .B(n644), .ZN(G45) );
  NAND2_X1 U724 ( .A1(n352), .A2(n647), .ZN(n646) );
  XNOR2_X1 U725 ( .A(n646), .B(G146), .ZN(G48) );
  XOR2_X1 U726 ( .A(G113), .B(KEYINPUT113), .Z(n649) );
  NAND2_X1 U727 ( .A1(n650), .A2(n647), .ZN(n648) );
  XNOR2_X1 U728 ( .A(n649), .B(n648), .ZN(G15) );
  NAND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n652), .B(G116), .ZN(G18) );
  XOR2_X1 U731 ( .A(G140), .B(n653), .Z(G42) );
  NAND2_X1 U732 ( .A1(KEYINPUT76), .A2(n654), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n655), .B(KEYINPUT2), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n661) );
  NAND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n664) );
  INV_X1 U736 ( .A(n662), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n666) );
  NAND2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n669), .B(KEYINPUT115), .ZN(n687) );
  NAND2_X1 U741 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U742 ( .A(KEYINPUT50), .B(n672), .ZN(n678) );
  NOR2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n676) );
  XNOR2_X1 U744 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U749 ( .A(KEYINPUT51), .B(n683), .Z(n685) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U752 ( .A(n688), .B(KEYINPUT52), .ZN(n689) );
  XNOR2_X1 U753 ( .A(KEYINPUT116), .B(n689), .ZN(n690) );
  NOR2_X1 U754 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U755 ( .A(KEYINPUT117), .B(n692), .Z(n693) );
  XNOR2_X1 U756 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n696) );
  XNOR2_X1 U757 ( .A(n694), .B(KEYINPUT57), .ZN(n695) );
  XNOR2_X1 U758 ( .A(n696), .B(n695), .ZN(n698) );
  XNOR2_X1 U759 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U760 ( .A1(n711), .A2(n699), .ZN(G54) );
  XOR2_X1 U761 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n700) );
  XNOR2_X1 U762 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U763 ( .A1(n711), .A2(n705), .ZN(G63) );
  XNOR2_X1 U764 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U765 ( .A1(n711), .A2(n710), .ZN(G66) );
  NAND2_X1 U766 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U767 ( .A1(G953), .A2(G224), .ZN(n714) );
  XNOR2_X1 U768 ( .A(KEYINPUT61), .B(n714), .ZN(n715) );
  NAND2_X1 U769 ( .A1(n715), .A2(G898), .ZN(n716) );
  NAND2_X1 U770 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U771 ( .A(n718), .B(KEYINPUT123), .ZN(n725) );
  XNOR2_X1 U772 ( .A(KEYINPUT122), .B(n719), .ZN(n721) );
  XNOR2_X1 U773 ( .A(n720), .B(n721), .ZN(n722) );
  NOR2_X1 U774 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U775 ( .A(n725), .B(n724), .Z(G69) );
  XNOR2_X1 U776 ( .A(n727), .B(n726), .ZN(n731) );
  XOR2_X1 U777 ( .A(G227), .B(n731), .Z(n728) );
  NAND2_X1 U778 ( .A1(n728), .A2(G900), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n729), .B(KEYINPUT124), .ZN(n730) );
  NAND2_X1 U780 ( .A1(n730), .A2(G953), .ZN(n736) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(n734) );
  NAND2_X1 U782 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n736), .A2(n735), .ZN(G72) );
  XNOR2_X1 U784 ( .A(n737), .B(G125), .ZN(n738) );
  XNOR2_X1 U785 ( .A(n738), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U786 ( .A(n739), .B(G122), .Z(G24) );
  XOR2_X1 U787 ( .A(G131), .B(KEYINPUT126), .Z(n740) );
  XNOR2_X1 U788 ( .A(n741), .B(n740), .ZN(G33) );
  XOR2_X1 U789 ( .A(n742), .B(G119), .Z(G21) );
  XOR2_X1 U790 ( .A(G134), .B(n743), .Z(G36) );
  XNOR2_X1 U791 ( .A(G137), .B(KEYINPUT125), .ZN(n745) );
  XNOR2_X1 U792 ( .A(n745), .B(n744), .ZN(G39) );
endmodule

