

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U324 ( .A(n414), .B(n413), .ZN(n535) );
  XNOR2_X1 U325 ( .A(n412), .B(KEYINPUT48), .ZN(n413) );
  XNOR2_X1 U326 ( .A(n352), .B(n351), .ZN(n353) );
  AND2_X1 U327 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U328 ( .A(n431), .B(KEYINPUT54), .ZN(n432) );
  XNOR2_X1 U329 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U330 ( .A(n346), .B(n292), .ZN(n347) );
  XNOR2_X1 U331 ( .A(n374), .B(n347), .ZN(n348) );
  XNOR2_X1 U332 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n456) );
  XNOR2_X1 U333 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U334 ( .A(n354), .B(n353), .ZN(n360) );
  XNOR2_X1 U335 ( .A(n380), .B(n379), .ZN(n401) );
  XOR2_X1 U336 ( .A(n310), .B(n309), .Z(n537) );
  XOR2_X1 U337 ( .A(KEYINPUT28), .B(n477), .Z(n540) );
  XNOR2_X1 U338 ( .A(n462), .B(G190GAT), .ZN(n463) );
  XNOR2_X1 U339 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT0), .B(KEYINPUT85), .Z(n314) );
  XOR2_X1 U341 ( .A(G99GAT), .B(G190GAT), .Z(n294) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(G134GAT), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U344 ( .A(n314), .B(n295), .Z(n297) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U347 ( .A(n298), .B(G120GAT), .Z(n302) );
  XOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n300) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n427) );
  XNOR2_X1 U351 ( .A(G113GAT), .B(n427), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n310) );
  XOR2_X1 U353 ( .A(KEYINPUT67), .B(G71GAT), .Z(n304) );
  XNOR2_X1 U354 ( .A(G15GAT), .B(G183GAT), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U356 ( .A(G127GAT), .B(G176GAT), .Z(n306) );
  XNOR2_X1 U357 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U359 ( .A(n308), .B(n307), .Z(n309) );
  INV_X1 U360 ( .A(n537), .ZN(n479) );
  XOR2_X1 U361 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n312) );
  NAND2_X1 U362 ( .A1(G225GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U364 ( .A(KEYINPUT4), .B(n313), .ZN(n326) );
  XOR2_X1 U365 ( .A(G1GAT), .B(G127GAT), .Z(n330) );
  XOR2_X1 U366 ( .A(G134GAT), .B(G162GAT), .Z(n346) );
  XOR2_X1 U367 ( .A(n330), .B(n346), .Z(n316) );
  XOR2_X1 U368 ( .A(G113GAT), .B(G141GAT), .Z(n384) );
  XNOR2_X1 U369 ( .A(n384), .B(n314), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U371 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n318) );
  XNOR2_X1 U372 ( .A(G29GAT), .B(G85GAT), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U374 ( .A(n320), .B(n319), .Z(n324) );
  XNOR2_X1 U375 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n321), .B(KEYINPUT3), .ZN(n441) );
  XNOR2_X1 U377 ( .A(G120GAT), .B(G148GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n322), .B(G57GAT), .ZN(n376) );
  XNOR2_X1 U379 ( .A(n441), .B(n376), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n475) );
  XNOR2_X1 U382 ( .A(KEYINPUT95), .B(n475), .ZN(n525) );
  XNOR2_X1 U383 ( .A(KEYINPUT69), .B(KEYINPUT45), .ZN(n363) );
  XNOR2_X1 U384 ( .A(G15GAT), .B(G22GAT), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n327), .B(KEYINPUT74), .ZN(n387) );
  XOR2_X1 U386 ( .A(G71GAT), .B(G78GAT), .Z(n328) );
  XNOR2_X1 U387 ( .A(KEYINPUT13), .B(n328), .ZN(n375) );
  XNOR2_X1 U388 ( .A(n387), .B(n375), .ZN(n343) );
  XNOR2_X1 U389 ( .A(G8GAT), .B(G183GAT), .ZN(n329) );
  XNOR2_X1 U390 ( .A(n329), .B(G211GAT), .ZN(n422) );
  XOR2_X1 U391 ( .A(n422), .B(n330), .Z(n332) );
  XNOR2_X1 U392 ( .A(G155GAT), .B(G57GAT), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U394 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n334) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U396 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U397 ( .A(n336), .B(n335), .Z(n341) );
  XOR2_X1 U398 ( .A(KEYINPUT83), .B(KEYINPUT12), .Z(n338) );
  XNOR2_X1 U399 ( .A(KEYINPUT14), .B(KEYINPUT81), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n339), .B(G64GAT), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U403 ( .A(n343), .B(n342), .Z(n497) );
  INV_X1 U404 ( .A(KEYINPUT80), .ZN(n361) );
  XOR2_X1 U405 ( .A(G92GAT), .B(G85GAT), .Z(n345) );
  XNOR2_X1 U406 ( .A(G99GAT), .B(G106GAT), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n374) );
  XOR2_X1 U408 ( .A(G190GAT), .B(G218GAT), .Z(n419) );
  XOR2_X1 U409 ( .A(n348), .B(n419), .Z(n354) );
  XOR2_X1 U410 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n350) );
  XNOR2_X1 U411 ( .A(KEYINPUT68), .B(KEYINPUT11), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n352) );
  XNOR2_X1 U413 ( .A(KEYINPUT10), .B(KEYINPUT79), .ZN(n351) );
  XNOR2_X1 U414 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n355), .B(G29GAT), .ZN(n356) );
  XOR2_X1 U416 ( .A(n356), .B(KEYINPUT8), .Z(n358) );
  XNOR2_X1 U417 ( .A(G43GAT), .B(G50GAT), .ZN(n357) );
  XOR2_X1 U418 ( .A(n358), .B(n357), .Z(n395) );
  INV_X1 U419 ( .A(n395), .ZN(n359) );
  XOR2_X1 U420 ( .A(n360), .B(n359), .Z(n562) );
  XNOR2_X1 U421 ( .A(n361), .B(n562), .ZN(n461) );
  XNOR2_X1 U422 ( .A(KEYINPUT36), .B(n461), .ZN(n582) );
  AND2_X1 U423 ( .A1(n497), .A2(n582), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n400) );
  XOR2_X1 U425 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n365) );
  XNOR2_X1 U426 ( .A(G204GAT), .B(KEYINPUT77), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n367) );
  INV_X1 U428 ( .A(n367), .ZN(n366) );
  XOR2_X1 U429 ( .A(G176GAT), .B(G64GAT), .Z(n417) );
  NAND2_X1 U430 ( .A1(n366), .A2(n417), .ZN(n370) );
  INV_X1 U431 ( .A(n417), .ZN(n368) );
  NAND2_X1 U432 ( .A1(n368), .A2(n367), .ZN(n369) );
  NAND2_X1 U433 ( .A1(n370), .A2(n369), .ZN(n372) );
  NAND2_X1 U434 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n373), .B(KEYINPUT78), .ZN(n380) );
  XOR2_X1 U437 ( .A(n374), .B(KEYINPUT31), .Z(n378) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U439 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n382) );
  XNOR2_X1 U440 ( .A(G1GAT), .B(G8GAT), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U442 ( .A(n383), .B(G197GAT), .Z(n386) );
  XNOR2_X1 U443 ( .A(G169GAT), .B(n384), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n391) );
  XOR2_X1 U445 ( .A(n387), .B(KEYINPUT73), .Z(n389) );
  NAND2_X1 U446 ( .A1(G229GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U448 ( .A(n391), .B(n390), .Z(n397) );
  XOR2_X1 U449 ( .A(KEYINPUT71), .B(KEYINPUT29), .Z(n393) );
  XNOR2_X1 U450 ( .A(KEYINPUT72), .B(KEYINPUT75), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U452 ( .A(n395), .B(n394), .Z(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n570) );
  XOR2_X1 U454 ( .A(KEYINPUT76), .B(n570), .Z(n564) );
  INV_X1 U455 ( .A(n564), .ZN(n398) );
  NAND2_X1 U456 ( .A1(n401), .A2(n398), .ZN(n399) );
  OR2_X1 U457 ( .A1(n400), .A2(n399), .ZN(n411) );
  XNOR2_X1 U458 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n409) );
  XOR2_X1 U459 ( .A(KEYINPUT109), .B(n497), .Z(n546) );
  XNOR2_X1 U460 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n402) );
  XOR2_X1 U461 ( .A(n402), .B(n401), .Z(n543) );
  INV_X1 U462 ( .A(n543), .ZN(n557) );
  NOR2_X1 U463 ( .A1(n557), .A2(n570), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n403), .B(KEYINPUT46), .ZN(n404) );
  NOR2_X1 U465 ( .A1(n546), .A2(n404), .ZN(n405) );
  XNOR2_X1 U466 ( .A(KEYINPUT110), .B(n405), .ZN(n406) );
  NAND2_X1 U467 ( .A1(n406), .A2(n562), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n407), .B(KEYINPUT112), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n410) );
  NAND2_X1 U470 ( .A1(n411), .A2(n410), .ZN(n414) );
  XNOR2_X1 U471 ( .A(KEYINPUT113), .B(KEYINPUT64), .ZN(n412) );
  XOR2_X1 U472 ( .A(G92GAT), .B(KEYINPUT96), .Z(n416) );
  NAND2_X1 U473 ( .A1(G226GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n418) );
  XOR2_X1 U475 ( .A(n418), .B(n417), .Z(n421) );
  XNOR2_X1 U476 ( .A(G36GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U478 ( .A(n423), .B(n422), .Z(n429) );
  XOR2_X1 U479 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n425) );
  XNOR2_X1 U480 ( .A(KEYINPUT89), .B(G204GAT), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U482 ( .A(G197GAT), .B(n426), .Z(n445) );
  XNOR2_X1 U483 ( .A(n427), .B(n445), .ZN(n428) );
  XOR2_X1 U484 ( .A(n429), .B(n428), .Z(n528) );
  INV_X1 U485 ( .A(n528), .ZN(n430) );
  NOR2_X1 U486 ( .A1(n535), .A2(n430), .ZN(n433) );
  XNOR2_X1 U487 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n431) );
  NOR2_X1 U488 ( .A1(n525), .A2(n434), .ZN(n567) );
  XOR2_X1 U489 ( .A(G148GAT), .B(G211GAT), .Z(n436) );
  XNOR2_X1 U490 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U492 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n438) );
  XNOR2_X1 U493 ( .A(G22GAT), .B(G141GAT), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n447) );
  XOR2_X1 U496 ( .A(n441), .B(G78GAT), .Z(n443) );
  NAND2_X1 U497 ( .A1(G228GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n455) );
  XOR2_X1 U501 ( .A(KEYINPUT93), .B(KEYINPUT87), .Z(n449) );
  XNOR2_X1 U502 ( .A(KEYINPUT23), .B(KEYINPUT88), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n453) );
  XOR2_X1 U504 ( .A(G106GAT), .B(G162GAT), .Z(n451) );
  XNOR2_X1 U505 ( .A(G50GAT), .B(G218GAT), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U507 ( .A(n453), .B(n452), .Z(n454) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(n477) );
  NAND2_X1 U509 ( .A1(n567), .A2(n477), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n457), .B(n456), .ZN(n458) );
  NOR2_X1 U511 ( .A1(n479), .A2(n458), .ZN(n565) );
  NAND2_X1 U512 ( .A1(n565), .A2(n546), .ZN(n460) );
  XNOR2_X1 U513 ( .A(KEYINPUT122), .B(G183GAT), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n460), .B(n459), .ZN(G1350GAT) );
  NAND2_X1 U515 ( .A1(n565), .A2(n461), .ZN(n464) );
  XOR2_X1 U516 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n462) );
  NAND2_X1 U517 ( .A1(n565), .A2(n543), .ZN(n467) );
  XOR2_X1 U518 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n465) );
  XNOR2_X1 U519 ( .A(n465), .B(G176GAT), .ZN(n466) );
  XNOR2_X1 U520 ( .A(n467), .B(n466), .ZN(G1349GAT) );
  NAND2_X1 U521 ( .A1(n564), .A2(n401), .ZN(n500) );
  NAND2_X1 U522 ( .A1(n528), .A2(n537), .ZN(n468) );
  NAND2_X1 U523 ( .A1(n468), .A2(n477), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT97), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT25), .ZN(n473) );
  XNOR2_X1 U526 ( .A(n528), .B(KEYINPUT27), .ZN(n478) );
  NOR2_X1 U527 ( .A1(n477), .A2(n537), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n471), .B(KEYINPUT26), .ZN(n568) );
  NAND2_X1 U529 ( .A1(n478), .A2(n568), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n476), .B(KEYINPUT98), .ZN(n482) );
  NAND2_X1 U533 ( .A1(n478), .A2(n525), .ZN(n534) );
  NOR2_X1 U534 ( .A1(n540), .A2(n534), .ZN(n480) );
  NAND2_X1 U535 ( .A1(n480), .A2(n479), .ZN(n481) );
  NAND2_X1 U536 ( .A1(n482), .A2(n481), .ZN(n495) );
  INV_X1 U537 ( .A(n497), .ZN(n578) );
  NOR2_X1 U538 ( .A1(n461), .A2(n578), .ZN(n484) );
  XNOR2_X1 U539 ( .A(KEYINPUT16), .B(KEYINPUT84), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U541 ( .A1(n495), .A2(n485), .ZN(n486) );
  XOR2_X1 U542 ( .A(KEYINPUT99), .B(n486), .Z(n511) );
  NOR2_X1 U543 ( .A1(n500), .A2(n511), .ZN(n493) );
  NAND2_X1 U544 ( .A1(n525), .A2(n493), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(KEYINPUT34), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NAND2_X1 U547 ( .A1(n528), .A2(n493), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n491) );
  NAND2_X1 U550 ( .A1(n493), .A2(n537), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(n492), .ZN(G1326GAT) );
  NAND2_X1 U553 ( .A1(n540), .A2(n493), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  NAND2_X1 U556 ( .A1(n582), .A2(n495), .ZN(n496) );
  NOR2_X1 U557 ( .A1(n497), .A2(n496), .ZN(n498) );
  XOR2_X1 U558 ( .A(KEYINPUT101), .B(n498), .Z(n499) );
  XNOR2_X1 U559 ( .A(KEYINPUT37), .B(n499), .ZN(n524) );
  NOR2_X1 U560 ( .A1(n524), .A2(n500), .ZN(n502) );
  XNOR2_X1 U561 ( .A(KEYINPUT38), .B(KEYINPUT102), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(n509) );
  NAND2_X1 U563 ( .A1(n509), .A2(n525), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NAND2_X1 U565 ( .A1(n528), .A2(n509), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n505), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n507) );
  NAND2_X1 U568 ( .A1(n509), .A2(n537), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NAND2_X1 U571 ( .A1(n540), .A2(n509), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n510), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n513) );
  NAND2_X1 U574 ( .A1(n570), .A2(n543), .ZN(n523) );
  NOR2_X1 U575 ( .A1(n511), .A2(n523), .ZN(n519) );
  NAND2_X1 U576 ( .A1(n519), .A2(n525), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n514), .Z(G1332GAT) );
  NAND2_X1 U579 ( .A1(n528), .A2(n519), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n517) );
  NAND2_X1 U582 ( .A1(n519), .A2(n537), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G71GAT), .B(n518), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U586 ( .A1(n519), .A2(n540), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U588 ( .A(G78GAT), .B(n522), .Z(G1335GAT) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n527) );
  NOR2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n531), .A2(n525), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n528), .A2(n531), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n531), .A2(n537), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U597 ( .A1(n540), .A2(n531), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n542) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(KEYINPUT114), .B(n536), .ZN(n553) );
  AND2_X1 U603 ( .A1(n553), .A2(n537), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(KEYINPUT115), .ZN(n539) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n564), .A2(n549), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U609 ( .A1(n549), .A2(n543), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NAND2_X1 U611 ( .A1(n549), .A2(n546), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U615 ( .A1(n549), .A2(n461), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U617 ( .A(G134GAT), .B(n552), .Z(G1343GAT) );
  NAND2_X1 U618 ( .A1(n553), .A2(n568), .ZN(n561) );
  NOR2_X1 U619 ( .A1(n570), .A2(n561), .ZN(n554) );
  XOR2_X1 U620 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n557), .A2(n561), .ZN(n558) );
  XOR2_X1 U625 ( .A(n559), .B(n558), .Z(G1345GAT) );
  NOR2_X1 U626 ( .A1(n578), .A2(n561), .ZN(n560) );
  XOR2_X1 U627 ( .A(G155GAT), .B(n560), .Z(G1346GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U633 ( .A(n569), .B(KEYINPUT124), .Z(n581) );
  INV_X1 U634 ( .A(n581), .ZN(n579) );
  NOR2_X1 U635 ( .A1(n579), .A2(n570), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U640 ( .A1(n579), .A2(n401), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

