//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n209), .B(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  OR2_X1    g0047(.A1(KEYINPUT8), .A2(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT66), .B(G58), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT8), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n214), .A2(G1), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G13), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n214), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n213), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT65), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(KEYINPUT65), .A3(new_n213), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n256), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n253), .A2(new_n262), .B1(new_n256), .B2(new_n251), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT16), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT64), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(new_n266), .B2(new_n267), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(KEYINPUT64), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT7), .B1(new_n278), .B2(new_n214), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT75), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n270), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(G20), .B1(new_n272), .B2(new_n277), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT75), .B1(new_n282), .B2(KEYINPUT7), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n218), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n210), .B1(new_n249), .B2(new_n218), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G20), .ZN(new_n286));
  INV_X1    g0086(.A(G159), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n286), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n265), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n257), .A2(KEYINPUT65), .A3(new_n213), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT65), .B1(new_n257), .B2(new_n213), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT7), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n275), .A2(new_n276), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(G20), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n218), .B1(new_n298), .B2(new_n269), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n295), .B1(new_n300), .B2(KEYINPUT16), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n264), .B1(new_n291), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G41), .ZN(new_n303));
  INV_X1    g0103(.A(G45), .ZN(new_n304));
  AOI21_X1  g0104(.A(G1), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G41), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G1), .A3(G13), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n307), .A3(G274), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n233), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G226), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G1698), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G223), .B2(G1698), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n314), .A2(new_n268), .B1(new_n274), .B2(new_n220), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT68), .B(G179), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(new_n321), .B2(new_n317), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n302), .A2(KEYINPUT18), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT18), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n266), .A2(new_n267), .A3(new_n271), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT64), .B1(new_n275), .B2(new_n276), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n214), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(new_n280), .A3(new_n296), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(new_n283), .A3(new_n269), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n290), .B1(new_n329), .B2(G68), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n301), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n263), .ZN(new_n332));
  INV_X1    g0132(.A(new_n322), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n324), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n323), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n308), .B1(new_n312), .B2(new_n310), .ZN(new_n336));
  INV_X1    g0136(.A(G1698), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n272), .A2(new_n277), .A3(G222), .A4(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n272), .A2(new_n277), .A3(G223), .A4(G1698), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n325), .A2(new_n326), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n338), .B(new_n339), .C1(new_n340), .C2(new_n224), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n336), .B1(new_n341), .B2(new_n316), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n321), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n214), .A2(G33), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n251), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n203), .A2(KEYINPUT67), .A3(G20), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT67), .ZN(new_n348));
  NOR3_X1   g0148(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n214), .ZN(new_n350));
  INV_X1    g0150(.A(G150), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n347), .B(new_n350), .C1(new_n351), .C2(new_n289), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n294), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n252), .A2(new_n202), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n262), .A2(new_n354), .B1(new_n202), .B2(new_n256), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n342), .B2(G169), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n344), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n272), .A2(new_n277), .A3(G232), .A4(new_n337), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n272), .A2(new_n277), .A3(G238), .A4(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n340), .C2(new_n226), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n316), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n307), .A2(G244), .A3(new_n309), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n308), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT69), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n308), .A2(new_n363), .A3(KEYINPUT69), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n362), .A2(new_n368), .A3(G190), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G20), .A2(G77), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT15), .B(G87), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT8), .B(G58), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n370), .B1(new_n371), .B2(new_n345), .C1(new_n289), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n294), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n262), .B(G77), .C1(G1), .C2(new_n214), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n256), .A2(new_n224), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n366), .A2(new_n367), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n316), .B2(new_n361), .ZN(new_n380));
  XOR2_X1   g0180(.A(KEYINPUT70), .B(G200), .Z(new_n381));
  OAI211_X1 g0181(.A(new_n369), .B(new_n378), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n362), .A2(new_n368), .A3(new_n320), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(new_n377), .C1(new_n380), .C2(G169), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT9), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n353), .A2(new_n386), .A3(new_n355), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n386), .B1(new_n353), .B2(new_n355), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n387), .A2(new_n388), .B1(new_n342), .B2(new_n381), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT71), .B1(new_n342), .B2(G190), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT10), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n388), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n353), .A2(new_n386), .A3(new_n355), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT10), .ZN(new_n396));
  INV_X1    g0196(.A(new_n381), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n343), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n395), .A2(new_n396), .A3(new_n390), .A4(new_n398), .ZN(new_n399));
  AOI211_X1 g0199(.A(new_n358), .B(new_n385), .C1(new_n392), .C2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G190), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n317), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(G200), .B2(new_n317), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n329), .A2(G68), .ZN(new_n404));
  INV_X1    g0204(.A(new_n290), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT16), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n300), .A2(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n294), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n263), .B(new_n403), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n331), .A2(KEYINPUT17), .A3(new_n263), .A4(new_n403), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n335), .A2(new_n400), .A3(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n224), .B2(new_n345), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n294), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT73), .B(KEYINPUT11), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT74), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  INV_X1    g0222(.A(G13), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(G1), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G20), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT12), .B1(new_n425), .B2(G68), .ZN(new_n426));
  OR3_X1    g0226(.A1(new_n425), .A2(KEYINPUT12), .A3(G68), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n252), .A2(new_n218), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n426), .A2(new_n427), .B1(new_n262), .B2(new_n428), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n421), .A2(new_n422), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT14), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n308), .B1(new_n219), .B2(new_n310), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n272), .A2(new_n277), .A3(G232), .A4(G1698), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n272), .A2(new_n277), .A3(G226), .A4(new_n337), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n437), .A2(KEYINPUT72), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(KEYINPUT72), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n433), .B1(new_n440), .B2(new_n316), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT13), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI211_X1 g0243(.A(KEYINPUT13), .B(new_n433), .C1(new_n440), .C2(new_n316), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n432), .B(G169), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n441), .A2(new_n442), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT72), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n340), .A2(new_n447), .A3(G226), .A4(new_n337), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n437), .A2(KEYINPUT72), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n307), .B1(new_n450), .B2(new_n436), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT13), .B1(new_n451), .B2(new_n433), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n446), .A2(new_n452), .A3(G179), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n445), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n446), .A2(new_n452), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n432), .B1(new_n455), .B2(G169), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n431), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G200), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n446), .B2(new_n452), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n430), .C1(new_n401), .C2(new_n455), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT76), .B1(new_n414), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n430), .B1(new_n455), .B2(new_n401), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n459), .ZN(new_n465));
  OAI21_X1  g0265(.A(G169), .B1(new_n443), .B2(new_n444), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT14), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(new_n453), .A3(new_n445), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n468), .B2(new_n431), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT18), .B1(new_n302), .B2(new_n322), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n332), .A2(new_n324), .A3(new_n333), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n411), .A4(new_n412), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n392), .A2(new_n399), .ZN(new_n473));
  INV_X1    g0273(.A(new_n358), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(new_n382), .A4(new_n384), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT76), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n469), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n463), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n256), .A2(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n254), .A2(G33), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n425), .B(new_n481), .C1(new_n292), .C2(new_n293), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n480), .B1(new_n482), .B2(G97), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT77), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g0285(.A(G97), .B(G107), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT6), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n487), .A2(new_n489), .A3(G107), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n491), .A2(new_n214), .B1(new_n224), .B2(new_n289), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n329), .B2(G107), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n485), .B1(new_n493), .B2(new_n295), .ZN(new_n494));
  OAI211_X1 g0294(.A(G244), .B(new_n337), .C1(new_n266), .C2(new_n267), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n495), .A2(new_n496), .B1(G33), .B2(G283), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n272), .A2(new_n277), .A3(G250), .A4(G1698), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n496), .A2(new_n225), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n272), .A2(new_n277), .A3(new_n337), .A4(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n501), .A2(new_n316), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n304), .A2(G1), .ZN(new_n503));
  AND2_X1   g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  NOR2_X1   g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G257), .A3(new_n307), .ZN(new_n507));
  OR2_X1    g0307(.A1(KEYINPUT5), .A2(G41), .ZN(new_n508));
  NAND2_X1  g0308(.A1(KEYINPUT5), .A2(G41), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n510), .A2(G274), .A3(new_n307), .A4(new_n503), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT78), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT78), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n507), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(G200), .B1(new_n502), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n512), .B1(new_n501), .B2(new_n316), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G190), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT79), .B1(new_n494), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n226), .B1(new_n281), .B2(new_n283), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n294), .B1(new_n522), .B2(new_n492), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n501), .A2(new_n316), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(new_n513), .A3(new_n515), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n525), .A2(G200), .B1(G190), .B2(new_n518), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT79), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n523), .A2(new_n526), .A3(new_n527), .A4(new_n485), .ZN(new_n528));
  INV_X1    g0328(.A(new_n518), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n523), .A2(new_n485), .B1(new_n318), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n516), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(KEYINPUT80), .A3(new_n320), .A4(new_n524), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n524), .A2(new_n320), .A3(new_n513), .A4(new_n515), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT80), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n521), .A2(new_n528), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n307), .A2(G274), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n503), .A2(new_n221), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n538), .A2(new_n503), .B1(new_n307), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G238), .B(new_n337), .C1(new_n266), .C2(new_n267), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n297), .A2(new_n544), .A3(G244), .A4(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(G244), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n320), .B(new_n540), .C1(new_n548), .C2(new_n307), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n214), .B1(new_n435), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n220), .A2(new_n489), .A3(new_n226), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n214), .B(G68), .C1(new_n266), .C2(new_n267), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n550), .B1(new_n345), .B2(new_n489), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n294), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n256), .A2(new_n371), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n371), .C2(new_n482), .ZN(new_n559));
  INV_X1    g0359(.A(new_n540), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n547), .A2(new_n545), .ZN(new_n561));
  INV_X1    g0361(.A(new_n543), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n563), .B2(new_n316), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n549), .B(new_n559), .C1(new_n564), .C2(G169), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n557), .A2(new_n558), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT82), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n482), .B2(new_n220), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n262), .A2(KEYINPUT82), .A3(G87), .A4(new_n481), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n307), .B1(new_n561), .B2(new_n562), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n397), .B1(new_n571), .B2(new_n560), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n572), .A3(KEYINPUT83), .ZN(new_n573));
  OAI211_X1 g0373(.A(G190), .B(new_n540), .C1(new_n548), .C2(new_n307), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT83), .B1(new_n570), .B2(new_n572), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n565), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n214), .B2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n226), .A2(KEYINPUT23), .A3(G20), .ZN(new_n581));
  INV_X1    g0381(.A(new_n542), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n580), .A2(new_n581), .B1(new_n582), .B2(new_n214), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n220), .A2(KEYINPUT22), .A3(G20), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n272), .A2(new_n277), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n214), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT22), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n585), .A2(new_n587), .A3(KEYINPUT87), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT87), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n583), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(KEYINPUT24), .B(new_n583), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n294), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n424), .A2(G20), .A3(new_n226), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT25), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n595), .B(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n226), .B2(new_n482), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT88), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT90), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n506), .A2(new_n307), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n227), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n506), .A2(KEYINPUT90), .A3(G264), .A4(new_n307), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(G250), .B(new_n337), .C1(new_n266), .C2(new_n267), .ZN(new_n606));
  NAND2_X1  g0406(.A1(G33), .A2(G294), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT89), .ZN(new_n609));
  NAND2_X1  g0409(.A1(G257), .A2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n268), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n297), .A2(KEYINPUT89), .A3(G257), .A4(G1698), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n605), .B(new_n511), .C1(new_n307), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n318), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n612), .ZN(new_n616));
  INV_X1    g0416(.A(new_n608), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n618), .A2(new_n316), .B1(new_n603), .B2(new_n604), .ZN(new_n619));
  INV_X1    g0419(.A(G179), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n620), .A3(new_n511), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n600), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n619), .A2(G190), .A3(new_n511), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n614), .A2(G200), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n594), .A2(new_n599), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n262), .A2(G116), .A3(new_n481), .ZN(new_n628));
  INV_X1    g0428(.A(G116), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n257), .A2(new_n213), .B1(G20), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(G33), .A2(G283), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n631), .B(new_n214), .C1(G33), .C2(new_n489), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT20), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(KEYINPUT20), .A3(new_n632), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n424), .A2(G20), .A3(new_n629), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n628), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(KEYINPUT84), .A2(G303), .ZN(new_n640));
  NOR2_X1   g0440(.A1(KEYINPUT84), .A2(G303), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n272), .B2(new_n277), .ZN(new_n643));
  OR2_X1    g0443(.A1(G257), .A2(G1698), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n227), .A2(G1698), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n644), .B(new_n645), .C1(new_n266), .C2(new_n267), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n316), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n316), .B1(new_n503), .B2(new_n510), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n254), .A2(G45), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n508), .B2(new_n509), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n649), .A2(G270), .B1(new_n538), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n639), .B(KEYINPUT86), .C1(new_n653), .C2(new_n458), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT86), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n458), .B1(new_n648), .B2(new_n652), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n628), .A2(new_n637), .A3(new_n638), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n652), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n654), .B(new_n658), .C1(new_n401), .C2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT21), .ZN(new_n661));
  AOI211_X1 g0461(.A(new_n661), .B(new_n318), .C1(new_n648), .C2(new_n652), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n659), .A2(new_n620), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT85), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n318), .B1(new_n648), .B2(new_n652), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n657), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n667), .B2(new_n661), .ZN(new_n668));
  AOI211_X1 g0468(.A(KEYINPUT85), .B(KEYINPUT21), .C1(new_n666), .C2(new_n657), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n660), .B(new_n664), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n627), .A2(new_n670), .ZN(new_n671));
  AND4_X1   g0471(.A1(new_n479), .A2(new_n537), .A3(new_n578), .A4(new_n671), .ZN(G372));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n323), .B2(new_n334), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n470), .A2(KEYINPUT91), .A3(new_n471), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n384), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n461), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n457), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n677), .B1(new_n413), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n473), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n474), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n529), .A2(new_n318), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n536), .A2(new_n494), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n565), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n684), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n576), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n573), .A3(new_n574), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n530), .A3(new_n536), .A4(new_n565), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n689), .B1(new_n692), .B2(new_n684), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n666), .A2(KEYINPUT21), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n653), .A2(G179), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n639), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n667), .A2(new_n661), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT85), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n667), .A2(new_n665), .A3(new_n661), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n623), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n521), .A2(new_n528), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n687), .A2(new_n565), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n626), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n701), .A2(new_n702), .A3(new_n704), .A4(new_n686), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n693), .A2(new_n705), .A3(new_n565), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n683), .B1(new_n479), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT92), .ZN(G369));
  XNOR2_X1  g0508(.A(KEYINPUT93), .B(G330), .ZN(new_n709));
  OR3_X1    g0509(.A1(new_n255), .A2(KEYINPUT27), .A3(G20), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT27), .B1(new_n255), .B2(G20), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G213), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G343), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n639), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n670), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n716), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n709), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n715), .B1(new_n594), .B2(new_n599), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n627), .A2(new_n721), .B1(new_n623), .B2(new_n715), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n627), .A2(new_n700), .A3(new_n714), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n615), .A2(new_n621), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n599), .B2(new_n594), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n724), .B1(new_n726), .B2(new_n715), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n723), .A2(new_n727), .ZN(G399));
  INV_X1    g0528(.A(new_n207), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n552), .A2(G116), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(G1), .A3(new_n732), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n733), .A2(KEYINPUT94), .B1(new_n211), .B2(new_n731), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(KEYINPUT94), .B2(new_n733), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT28), .Z(new_n736));
  NAND2_X1  g0536(.A1(new_n702), .A2(new_n686), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n626), .B(new_n703), .C1(new_n726), .C2(new_n718), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n565), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n684), .B1(new_n577), .B2(new_n686), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n530), .A2(KEYINPUT26), .A3(new_n536), .A4(new_n703), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT29), .B(new_n715), .C1(new_n739), .C2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT29), .B1(new_n706), .B2(new_n715), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n671), .A2(new_n537), .A3(new_n578), .A4(new_n715), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n619), .A2(new_n564), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n748), .A2(KEYINPUT30), .A3(new_n518), .A4(new_n663), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n663), .A2(new_n518), .A3(new_n564), .A4(new_n619), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n653), .A2(new_n321), .ZN(new_n753));
  INV_X1    g0553(.A(new_n564), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n753), .A2(new_n754), .A3(new_n525), .A4(new_n614), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n749), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n756), .A2(KEYINPUT31), .A3(new_n714), .ZN(new_n757));
  AOI21_X1  g0557(.A(KEYINPUT31), .B1(new_n756), .B2(new_n714), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n747), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n709), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n746), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n736), .B1(new_n764), .B2(G1), .ZN(G364));
  INV_X1    g0565(.A(new_n720), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n717), .A2(new_n709), .A3(new_n719), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n423), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n254), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n730), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n766), .A2(new_n767), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n214), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n397), .A2(new_n401), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(G283), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n401), .A2(G200), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n214), .B1(new_n778), .B2(new_n620), .ZN(new_n779));
  INV_X1    g0579(.A(G294), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G190), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n774), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G329), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n779), .A2(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n320), .A2(new_n214), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT95), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n778), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n777), .B(new_n784), .C1(new_n788), .C2(G322), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n786), .A2(G190), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G326), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n786), .A2(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G190), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT33), .B(G317), .Z(new_n796));
  OAI211_X1 g0596(.A(new_n789), .B(new_n792), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n786), .A2(new_n781), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n397), .A2(G190), .A3(new_n774), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n278), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n798), .A2(G311), .B1(KEYINPUT97), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(KEYINPUT97), .B2(new_n801), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n779), .B(KEYINPUT96), .Z(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G97), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n775), .A2(new_n226), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n278), .ZN(new_n807));
  INV_X1    g0607(.A(new_n799), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G87), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n782), .A2(new_n287), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT32), .ZN(new_n811));
  AND4_X1   g0611(.A1(new_n805), .A2(new_n807), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n798), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n224), .B2(new_n813), .C1(new_n249), .C2(new_n787), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n795), .A2(new_n218), .B1(new_n202), .B2(new_n790), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n797), .A2(new_n803), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n213), .B1(G20), .B2(new_n318), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G13), .A2(G33), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(G20), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n717), .A2(new_n719), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n817), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n278), .A2(new_n729), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G355), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G116), .B2(new_n207), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n729), .A2(new_n297), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(G45), .B2(new_n211), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n246), .B2(G45), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n823), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n818), .A2(new_n822), .A3(new_n771), .A4(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n773), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  INV_X1    g0633(.A(new_n817), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n820), .ZN(new_n835));
  XOR2_X1   g0635(.A(KEYINPUT98), .B(G283), .Z(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n794), .A2(new_n837), .B1(new_n791), .B2(G303), .ZN(new_n838));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n278), .B1(new_n839), .B2(new_n782), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n775), .A2(new_n220), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n840), .B(new_n841), .C1(G107), .C2(new_n808), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G294), .A2(new_n788), .B1(new_n798), .B2(G116), .ZN(new_n843));
  AND4_X1   g0643(.A1(new_n805), .A2(new_n838), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G143), .A2(new_n788), .B1(new_n798), .B2(G159), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n845), .B1(new_n846), .B2(new_n790), .C1(new_n351), .C2(new_n795), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT34), .ZN(new_n848));
  INV_X1    g0648(.A(G132), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n297), .B1(new_n782), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT99), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n776), .A2(G68), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n249), .B2(new_n779), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n851), .B(new_n853), .C1(G50), .C2(new_n808), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n844), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n771), .B1(G77), .B2(new_n835), .C1(new_n855), .C2(new_n834), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n377), .A2(new_n714), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n382), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(new_n678), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n384), .A2(new_n714), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n856), .A2(KEYINPUT100), .B1(new_n820), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n856), .A2(KEYINPUT100), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n706), .A2(new_n715), .ZN(new_n865));
  INV_X1    g0665(.A(new_n861), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n706), .A2(new_n715), .A3(new_n861), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n762), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT102), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n763), .A2(new_n867), .A3(new_n868), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT101), .B1(new_n872), .B2(new_n772), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(KEYINPUT101), .A3(new_n772), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n864), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(G384));
  OAI211_X1 g0677(.A(new_n431), .B(new_n714), .C1(new_n468), .C2(new_n465), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n431), .A2(new_n714), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n457), .A2(new_n461), .A3(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n860), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n882), .B2(new_n868), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n301), .B1(KEYINPUT16), .B2(new_n300), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n712), .B1(new_n884), .B2(new_n263), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n472), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT104), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n472), .A2(KEYINPUT104), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n332), .A2(new_n333), .ZN(new_n891));
  INV_X1    g0691(.A(new_n712), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n332), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n891), .A2(new_n893), .A3(new_n894), .A4(new_n409), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n884), .A2(new_n263), .B1(new_n322), .B2(new_n712), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n302), .B2(new_n403), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n897), .B2(new_n894), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n890), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n472), .A2(KEYINPUT104), .A3(new_n885), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT104), .B1(new_n472), .B2(new_n885), .ZN(new_n901));
  OAI211_X1 g0701(.A(KEYINPUT38), .B(new_n898), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n883), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n677), .A2(new_n712), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n409), .B1(new_n302), .B2(new_n322), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n302), .A2(new_n712), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n895), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n323), .A2(new_n334), .A3(new_n673), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT91), .B1(new_n470), .B2(new_n471), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n413), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n911), .B1(new_n914), .B2(new_n909), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n902), .B(new_n907), .C1(new_n915), .C2(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT105), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT39), .B1(new_n899), .B2(new_n903), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n893), .B1(new_n676), .B2(new_n413), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n919), .B1(new_n920), .B2(new_n911), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(new_n907), .A4(new_n902), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n917), .A2(new_n918), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n468), .A2(new_n431), .A3(new_n715), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n906), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT107), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT106), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n414), .A2(new_n462), .A3(KEYINPUT76), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n477), .B1(new_n469), .B2(new_n476), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n565), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n626), .A2(new_n703), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n623), .B2(new_n700), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n935), .B2(new_n537), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n714), .B1(new_n936), .B2(new_n693), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n743), .B1(new_n937), .B2(KEYINPUT29), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n929), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT29), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n865), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n479), .A2(new_n941), .A3(KEYINPUT106), .A4(new_n743), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n683), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n928), .B(new_n943), .Z(new_n944));
  NOR2_X1   g0744(.A1(new_n899), .A2(new_n903), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n866), .B1(new_n878), .B2(new_n880), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n947), .A3(new_n760), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n878), .A2(new_n880), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(new_n760), .A3(new_n861), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n921), .B2(new_n902), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n945), .A2(new_n948), .B1(new_n951), .B2(new_n947), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n479), .A2(new_n760), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n952), .B(new_n953), .Z(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n709), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n944), .A2(new_n955), .B1(new_n254), .B2(new_n768), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n944), .B2(new_n955), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n212), .B(G77), .C1(new_n218), .C2(new_n249), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n202), .A2(G68), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n254), .B(G13), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n491), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT35), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(KEYINPUT35), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n962), .A2(G116), .A3(new_n215), .A4(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT103), .B(KEYINPUT36), .Z(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  OR3_X1    g0766(.A1(new_n957), .A2(new_n960), .A3(new_n966), .ZN(G367));
  INV_X1    g0767(.A(KEYINPUT110), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT42), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n494), .A2(new_n714), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n537), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n530), .A2(new_n536), .A3(new_n714), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT108), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(KEYINPUT108), .A3(new_n972), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n969), .B1(new_n976), .B2(new_n724), .ZN(new_n977));
  INV_X1    g0777(.A(new_n975), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(new_n973), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n686), .B1(new_n979), .B2(new_n623), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n977), .B1(new_n980), .B2(new_n715), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n969), .B(new_n724), .C1(new_n978), .C2(new_n973), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT109), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n968), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n981), .A2(new_n984), .A3(new_n968), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n570), .A2(new_n715), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n933), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n688), .B2(new_n988), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n986), .A2(new_n987), .A3(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n990), .B(KEYINPUT43), .Z(new_n993));
  INV_X1    g0793(.A(new_n987), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(new_n985), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n979), .A2(new_n723), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT111), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n992), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(KEYINPUT111), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n730), .B(KEYINPUT41), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n727), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n979), .B(new_n1003), .C1(KEYINPUT112), .C2(KEYINPUT44), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n976), .B2(new_n727), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n979), .B2(new_n1003), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n976), .A2(KEYINPUT45), .A3(new_n727), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AND3_X1   g0812(.A1(new_n1008), .A2(new_n1012), .A3(new_n723), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n723), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n724), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n700), .A2(new_n714), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1015), .B1(new_n722), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(new_n720), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1018), .A2(new_n938), .A3(new_n762), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1013), .A2(new_n1014), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n764), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1002), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n769), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n992), .A2(new_n995), .A3(KEYINPUT111), .A4(new_n996), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1000), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AND3_X1   g0825(.A1(new_n808), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1026));
  AOI21_X1  g0826(.A(KEYINPUT46), .B1(new_n808), .B2(G116), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n775), .A2(new_n489), .ZN(new_n1028));
  INV_X1    g0828(.A(G317), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n268), .B1(new_n782), .B2(new_n1029), .C1(new_n779), .C2(new_n226), .ZN(new_n1030));
  NOR4_X1   g0830(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n642), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1032), .A2(new_n788), .B1(new_n798), .B2(new_n837), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT113), .B(G311), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n791), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n794), .A2(G294), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n804), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1038), .A2(new_n218), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n775), .A2(new_n224), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n782), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n278), .B(new_n1040), .C1(G137), .C2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n249), .B2(new_n799), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1039), .B(new_n1043), .C1(G150), .C2(new_n788), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n795), .A2(new_n287), .B1(new_n813), .B2(new_n202), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(KEYINPUT114), .ZN(new_n1046));
  INV_X1    g0846(.A(G143), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1044), .B(new_n1046), .C1(new_n1047), .C2(new_n790), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1045), .A2(KEYINPUT114), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1037), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT115), .Z(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT47), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT47), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n817), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n239), .A2(new_n827), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n371), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n817), .B(new_n821), .C1(new_n729), .C2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n772), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n821), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1054), .B(new_n1058), .C1(new_n1059), .C2(new_n990), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1025), .A2(new_n1060), .ZN(G387));
  NOR2_X1   g0861(.A1(new_n722), .A2(new_n1059), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n236), .A2(new_n304), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n732), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1063), .A2(new_n827), .B1(new_n1064), .B2(new_n824), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n372), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n202), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1067), .A2(KEYINPUT50), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1067), .A2(KEYINPUT50), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n732), .B(new_n304), .C1(new_n218), .C2(new_n224), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1065), .A2(new_n1071), .B1(G107), .B2(new_n207), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n823), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n771), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1038), .A2(new_n371), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n799), .A2(new_n224), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n297), .B1(new_n782), .B2(new_n351), .ZN(new_n1077));
  NOR4_X1   g0877(.A1(new_n1075), .A2(new_n1028), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n251), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1079), .A2(new_n794), .B1(new_n791), .B2(G159), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G50), .A2(new_n788), .B1(new_n798), .B2(G68), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G317), .A2(new_n788), .B1(new_n798), .B2(new_n1032), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n794), .A2(new_n1034), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n791), .A2(G322), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n799), .A2(new_n780), .B1(new_n779), .B2(new_n836), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(KEYINPUT49), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n297), .B1(new_n1041), .B2(G326), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(new_n629), .C2(new_n775), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT49), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1082), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1062), .B(new_n1074), .C1(new_n1095), .C2(new_n817), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n770), .B2(new_n1018), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n764), .A2(new_n1018), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1019), .A2(new_n730), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(G393));
  NAND2_X1  g0900(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n723), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1008), .A2(new_n1012), .A3(new_n723), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1103), .A2(new_n764), .A3(new_n1018), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1019), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n1106), .A3(new_n730), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n243), .A2(new_n827), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1108), .B(new_n823), .C1(new_n489), .C2(new_n207), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n340), .B1(G322), .B2(new_n1041), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n629), .B2(new_n779), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n806), .B(new_n1111), .C1(new_n808), .C2(new_n837), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n780), .B2(new_n813), .C1(new_n642), .C2(new_n795), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n790), .A2(new_n1029), .B1(new_n787), .B2(new_n839), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT116), .Z(new_n1115));
  AOI21_X1  g0915(.A(new_n1113), .B1(new_n1115), .B2(KEYINPUT52), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1115), .A2(KEYINPUT52), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n790), .A2(new_n351), .B1(new_n787), .B2(new_n287), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT51), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n297), .B1(new_n782), .B2(new_n1047), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1120), .B(new_n841), .C1(G68), .C2(new_n808), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n804), .A2(G77), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(new_n372), .C2(new_n813), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G50), .B2(new_n794), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1116), .A2(new_n1117), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n771), .B(new_n1109), .C1(new_n1125), .C2(new_n834), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT117), .Z(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n821), .B2(new_n979), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n770), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1107), .A2(new_n1130), .ZN(G390));
  OAI21_X1  g0931(.A(new_n771), .B1(new_n1079), .B2(new_n835), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT54), .B(G143), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n813), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n799), .A2(new_n351), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT53), .Z(new_n1136));
  AOI21_X1  g0936(.A(new_n278), .B1(G125), .B2(new_n1041), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n202), .B2(new_n775), .C1(new_n1038), .C2(new_n287), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n787), .A2(new_n849), .ZN(new_n1139));
  OR4_X1    g0939(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n791), .A2(G128), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n795), .B2(new_n846), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G116), .A2(new_n788), .B1(new_n798), .B2(G97), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1041), .A2(G294), .ZN(new_n1144));
  AND4_X1   g0944(.A1(new_n278), .A2(new_n809), .A3(new_n852), .A4(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1122), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n791), .A2(G283), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n795), .B2(new_n226), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1140), .A2(new_n1142), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1132), .B1(new_n1149), .B2(new_n817), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n924), .B2(new_n820), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT119), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n860), .B1(new_n937), .B2(new_n861), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n925), .B1(new_n1153), .B2(new_n881), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n917), .A2(new_n918), .A3(new_n923), .A4(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n902), .B1(new_n915), .B2(KEYINPUT38), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n715), .B1(new_n678), .B2(new_n858), .C1(new_n739), .C2(new_n742), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1157), .A2(new_n882), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1156), .B(new_n925), .C1(new_n881), .C2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n760), .A2(new_n761), .A3(new_n861), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1160), .A2(new_n881), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1155), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(G330), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n747), .B2(new_n759), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n946), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n770), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n683), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1164), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n478), .B2(new_n463), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT106), .B1(new_n746), .B2(new_n479), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n942), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1169), .B(new_n1172), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n882), .B(new_n1157), .C1(new_n1160), .C2(new_n881), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n949), .B1(new_n1164), .B2(new_n861), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1160), .A2(new_n881), .B1(new_n946), .B2(new_n1164), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1176), .A2(new_n1177), .B1(new_n1178), .B2(new_n1153), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT118), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT118), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n943), .A2(new_n1182), .A3(new_n1179), .A4(new_n1172), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n730), .B1(new_n1167), .B2(new_n1184), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n683), .B(new_n1171), .C1(new_n939), .C2(new_n942), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1182), .B1(new_n1186), .B2(new_n1179), .ZN(new_n1187));
  AND4_X1   g0987(.A1(new_n1182), .A2(new_n943), .A3(new_n1172), .A4(new_n1179), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1165), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1155), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1189), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1152), .B(new_n1168), .C1(new_n1185), .C2(new_n1195), .ZN(G378));
  NAND2_X1  g0996(.A1(new_n924), .A2(new_n926), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n906), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n473), .A2(new_n474), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n356), .A2(new_n892), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1202), .B(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n950), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n947), .B1(new_n1156), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n919), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n948), .B1(new_n1208), .B2(new_n902), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1204), .B(G330), .C1(new_n1206), .C2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1204), .B1(new_n952), .B2(G330), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1199), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(G330), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1204), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n927), .A2(new_n1216), .A3(new_n1210), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1213), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n819), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n771), .B1(new_n835), .B2(G50), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n297), .A2(G41), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G50), .B(new_n1221), .C1(new_n274), .C2(new_n303), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n775), .A2(new_n249), .ZN(new_n1223));
  INV_X1    g1023(.A(G283), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1221), .B1(new_n1224), .B2(new_n782), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1039), .A2(new_n1076), .A3(new_n1223), .A4(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G97), .A2(new_n794), .B1(new_n791), .B2(G116), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G107), .A2(new_n788), .B1(new_n798), .B2(new_n1056), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT58), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1222), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n788), .A2(G128), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1133), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n804), .A2(G150), .B1(new_n808), .B2(new_n1233), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(new_n813), .C2(new_n846), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n795), .A2(new_n849), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(G125), .C2(new_n791), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(KEYINPUT59), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(KEYINPUT120), .B(G124), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n274), .B(new_n303), .C1(new_n782), .C2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n776), .B2(G159), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT59), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1242), .B1(new_n1237), .B2(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1231), .B1(new_n1230), .B2(new_n1229), .C1(new_n1239), .C2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1220), .B1(new_n1245), .B2(new_n817), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1218), .A2(new_n770), .B1(new_n1219), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1218), .A2(KEYINPUT57), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1175), .B1(new_n1167), .B2(new_n1184), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n730), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1186), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1251), .B2(new_n1218), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1247), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT121), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(KEYINPUT121), .B(new_n1247), .C1(new_n1250), .C2(new_n1252), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(G375));
  NAND2_X1  g1058(.A1(new_n1179), .A2(new_n770), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n771), .B1(new_n835), .B2(G68), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n268), .B(new_n1223), .C1(G128), .C2(new_n1041), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n287), .B2(new_n799), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G50), .B2(new_n804), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G137), .A2(new_n788), .B1(new_n798), .B2(G150), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n795), .C2(new_n1133), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n791), .A2(G132), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT123), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1075), .B1(new_n788), .B2(G283), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT122), .Z(new_n1269));
  OAI21_X1  g1069(.A(new_n278), .B1(new_n800), .B2(new_n782), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1270), .B(new_n1040), .C1(G97), .C2(new_n808), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n798), .A2(G107), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n1273), .B1(new_n629), .B2(new_n795), .C1(new_n780), .C2(new_n790), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n1265), .A2(new_n1267), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1260), .B1(new_n1275), .B2(new_n817), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n949), .B2(new_n820), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1259), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1181), .A2(new_n1183), .A3(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1279), .B1(new_n1281), .B2(new_n1001), .ZN(G381));
  INV_X1    g1082(.A(G378), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1097), .B(new_n832), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1284));
  OR2_X1    g1084(.A1(G384), .A2(new_n1284), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(G387), .A2(new_n1285), .A3(G390), .A4(G381), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1257), .A2(new_n1283), .A3(new_n1286), .ZN(G407));
  NAND2_X1  g1087(.A1(new_n1257), .A2(new_n1283), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(new_n1288), .C2(G343), .ZN(G409));
  NAND2_X1  g1089(.A1(new_n713), .A2(G213), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT124), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n927), .A2(new_n1216), .A3(new_n1210), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n927), .B1(new_n1210), .B2(new_n1216), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1002), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1292), .B1(new_n1295), .B2(new_n1249), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1001), .B1(new_n1213), .B2(new_n1217), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1251), .A2(new_n1297), .A3(KEYINPUT124), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1247), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1283), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G378), .B(new_n1247), .C1(new_n1250), .C2(new_n1252), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1291), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1281), .A2(KEYINPUT60), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1280), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1303), .B(new_n730), .C1(KEYINPUT60), .C2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G384), .B1(new_n1305), .B2(new_n1279), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n730), .B1(new_n1304), .B2(KEYINPUT60), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(KEYINPUT60), .B2(new_n1281), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1308), .A2(new_n876), .A3(new_n1278), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1302), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1291), .A2(G2897), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1305), .A2(G384), .A3(new_n1279), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n876), .B1(new_n1308), .B2(new_n1278), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1317), .A2(new_n1318), .A3(new_n1314), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n1302), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1302), .A2(KEYINPUT63), .A3(new_n1310), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G393), .A2(G396), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1284), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1107), .A2(new_n1130), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1107), .B2(new_n1130), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1327), .A2(new_n1025), .A3(new_n1060), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1326), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1107), .A2(new_n1130), .A3(new_n1324), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1025), .A2(new_n1060), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1328), .A2(new_n1331), .A3(KEYINPUT61), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1313), .A2(new_n1321), .A3(new_n1322), .A4(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1302), .A2(new_n1334), .A3(new_n1310), .ZN(new_n1335));
  XOR2_X1   g1135(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1302), .B2(new_n1320), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1334), .B1(new_n1302), .B2(new_n1310), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1335), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT126), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1340), .B1(new_n1328), .B2(new_n1331), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1327), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(G387), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1327), .A2(new_n1025), .A3(new_n1060), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(KEYINPUT126), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1341), .A2(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1333), .B1(new_n1339), .B2(new_n1346), .ZN(G405));
  INV_X1    g1147(.A(KEYINPUT127), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1341), .A2(new_n1348), .A3(new_n1345), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1348), .B1(new_n1341), .B2(new_n1345), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1310), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1253), .A2(G378), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1352), .B1(new_n1288), .B2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(G378), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1353), .ZN(new_n1356));
  NOR3_X1   g1156(.A1(new_n1355), .A2(new_n1310), .A3(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1351), .B1(new_n1354), .B2(new_n1357), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1288), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1310), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1359), .A2(new_n1349), .A3(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1358), .A2(new_n1361), .ZN(G402));
endmodule


