

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U557 ( .A(n549), .B(KEYINPUT65), .ZN(G160) );
  NOR2_X1 U558 ( .A1(n611), .A2(n725), .ZN(n655) );
  NOR2_X1 U559 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U560 ( .A1(G8), .A2(n680), .ZN(n714) );
  NOR2_X1 U561 ( .A1(n678), .A2(n677), .ZN(n527) );
  NOR2_X1 U562 ( .A1(n677), .A2(n676), .ZN(n612) );
  INV_X1 U563 ( .A(KEYINPUT28), .ZN(n629) );
  INV_X1 U564 ( .A(KEYINPUT31), .ZN(n622) );
  XNOR2_X1 U565 ( .A(n623), .B(n622), .ZN(n685) );
  INV_X1 U566 ( .A(n984), .ZN(n716) );
  NOR2_X1 U567 ( .A1(n716), .A2(n715), .ZN(n717) );
  INV_X1 U568 ( .A(KEYINPUT105), .ZN(n719) );
  XNOR2_X1 U569 ( .A(n720), .B(n719), .ZN(n721) );
  INV_X1 U570 ( .A(KEYINPUT17), .ZN(n535) );
  NAND2_X1 U571 ( .A1(n913), .A2(G137), .ZN(n542) );
  AND2_X2 U572 ( .A1(G2104), .A2(G2105), .ZN(n916) );
  XNOR2_X1 U573 ( .A(n540), .B(n539), .ZN(G164) );
  INV_X1 U574 ( .A(KEYINPUT94), .ZN(n540) );
  INV_X1 U575 ( .A(G2105), .ZN(n528) );
  AND2_X1 U576 ( .A1(n528), .A2(G2104), .ZN(n912) );
  NAND2_X1 U577 ( .A1(G102), .A2(n912), .ZN(n531) );
  NOR2_X1 U578 ( .A1(n528), .A2(G2104), .ZN(n529) );
  XNOR2_X1 U579 ( .A(n529), .B(KEYINPUT66), .ZN(n729) );
  NAND2_X1 U580 ( .A1(n729), .A2(G126), .ZN(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n534) );
  NAND2_X1 U582 ( .A1(G114), .A2(n916), .ZN(n532) );
  XNOR2_X1 U583 ( .A(KEYINPUT93), .B(n532), .ZN(n533) );
  NOR2_X1 U584 ( .A1(n534), .A2(n533), .ZN(n538) );
  NOR2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  XNOR2_X2 U586 ( .A(n536), .B(n535), .ZN(n913) );
  NAND2_X1 U587 ( .A1(n913), .A2(G138), .ZN(n537) );
  NAND2_X1 U588 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U589 ( .A1(G125), .A2(n729), .ZN(n541) );
  NAND2_X1 U590 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U591 ( .A1(G113), .A2(n916), .ZN(n543) );
  XNOR2_X1 U592 ( .A(KEYINPUT67), .B(n543), .ZN(n544) );
  NOR2_X1 U593 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U594 ( .A1(G101), .A2(n912), .ZN(n546) );
  XOR2_X1 U595 ( .A(KEYINPUT23), .B(n546), .Z(n547) );
  NAND2_X1 U596 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U597 ( .A(KEYINPUT0), .B(G543), .Z(n598) );
  NOR2_X1 U598 ( .A1(G651), .A2(n598), .ZN(n550) );
  XNOR2_X1 U599 ( .A(KEYINPUT64), .B(n550), .ZN(n811) );
  NAND2_X1 U600 ( .A1(G51), .A2(n811), .ZN(n551) );
  XNOR2_X1 U601 ( .A(n551), .B(KEYINPUT78), .ZN(n555) );
  INV_X1 U602 ( .A(G651), .ZN(n558) );
  NOR2_X1 U603 ( .A1(G543), .A2(n558), .ZN(n552) );
  XOR2_X1 U604 ( .A(KEYINPUT68), .B(n552), .Z(n553) );
  XNOR2_X1 U605 ( .A(KEYINPUT1), .B(n553), .ZN(n812) );
  NAND2_X1 U606 ( .A1(G63), .A2(n812), .ZN(n554) );
  NAND2_X1 U607 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U608 ( .A(KEYINPUT6), .B(n556), .ZN(n564) );
  NOR2_X1 U609 ( .A1(G651), .A2(G543), .ZN(n815) );
  NAND2_X1 U610 ( .A1(n815), .A2(G89), .ZN(n557) );
  XNOR2_X1 U611 ( .A(n557), .B(KEYINPUT4), .ZN(n560) );
  NOR2_X1 U612 ( .A1(n598), .A2(n558), .ZN(n816) );
  NAND2_X1 U613 ( .A1(G76), .A2(n816), .ZN(n559) );
  NAND2_X1 U614 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U615 ( .A(KEYINPUT5), .B(n561), .ZN(n562) );
  XNOR2_X1 U616 ( .A(KEYINPUT77), .B(n562), .ZN(n563) );
  NOR2_X1 U617 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U618 ( .A(KEYINPUT7), .B(n565), .Z(G168) );
  NAND2_X1 U619 ( .A1(G52), .A2(n811), .ZN(n567) );
  NAND2_X1 U620 ( .A1(G64), .A2(n812), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U622 ( .A1(G90), .A2(n815), .ZN(n569) );
  NAND2_X1 U623 ( .A1(G77), .A2(n816), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U625 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  NOR2_X1 U626 ( .A1(n572), .A2(n571), .ZN(G171) );
  NAND2_X1 U627 ( .A1(G91), .A2(n815), .ZN(n574) );
  NAND2_X1 U628 ( .A1(G78), .A2(n816), .ZN(n573) );
  NAND2_X1 U629 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U630 ( .A(KEYINPUT69), .B(n575), .ZN(n579) );
  NAND2_X1 U631 ( .A1(n811), .A2(G53), .ZN(n577) );
  NAND2_X1 U632 ( .A1(n812), .A2(G65), .ZN(n576) );
  AND2_X1 U633 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n579), .A2(n578), .ZN(G299) );
  NAND2_X1 U635 ( .A1(n815), .A2(G88), .ZN(n580) );
  XNOR2_X1 U636 ( .A(n580), .B(KEYINPUT84), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G75), .A2(n816), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U639 ( .A(n583), .B(KEYINPUT85), .ZN(n585) );
  NAND2_X1 U640 ( .A1(G50), .A2(n811), .ZN(n584) );
  NAND2_X1 U641 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U642 ( .A1(G62), .A2(n812), .ZN(n586) );
  XNOR2_X1 U643 ( .A(KEYINPUT83), .B(n586), .ZN(n587) );
  NOR2_X1 U644 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U645 ( .A(KEYINPUT86), .B(n589), .ZN(G166) );
  INV_X1 U646 ( .A(G166), .ZN(G303) );
  XOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U648 ( .A1(n815), .A2(G86), .ZN(n591) );
  NAND2_X1 U649 ( .A1(G61), .A2(n812), .ZN(n590) );
  NAND2_X1 U650 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U651 ( .A(KEYINPUT82), .B(n592), .ZN(n595) );
  NAND2_X1 U652 ( .A1(n816), .A2(G73), .ZN(n593) );
  XOR2_X1 U653 ( .A(KEYINPUT2), .B(n593), .Z(n594) );
  NOR2_X1 U654 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U655 ( .A1(G48), .A2(n811), .ZN(n596) );
  NAND2_X1 U656 ( .A1(n597), .A2(n596), .ZN(G305) );
  NAND2_X1 U657 ( .A1(G49), .A2(n811), .ZN(n603) );
  NAND2_X1 U658 ( .A1(G87), .A2(n598), .ZN(n600) );
  NAND2_X1 U659 ( .A1(G74), .A2(G651), .ZN(n599) );
  NAND2_X1 U660 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U661 ( .A1(n812), .A2(n601), .ZN(n602) );
  NAND2_X1 U662 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U663 ( .A(KEYINPUT81), .B(n604), .Z(G288) );
  NAND2_X1 U664 ( .A1(G47), .A2(n811), .ZN(n606) );
  NAND2_X1 U665 ( .A1(G60), .A2(n812), .ZN(n605) );
  NAND2_X1 U666 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U667 ( .A1(G85), .A2(n815), .ZN(n608) );
  NAND2_X1 U668 ( .A1(G72), .A2(n816), .ZN(n607) );
  NAND2_X1 U669 ( .A1(n608), .A2(n607), .ZN(n609) );
  OR2_X1 U670 ( .A1(n610), .A2(n609), .ZN(G290) );
  NOR2_X1 U671 ( .A1(G1384), .A2(G164), .ZN(n726) );
  INV_X1 U672 ( .A(n726), .ZN(n611) );
  NAND2_X1 U673 ( .A1(G160), .A2(G40), .ZN(n725) );
  INV_X1 U674 ( .A(n655), .ZN(n680) );
  NOR2_X1 U675 ( .A1(G1966), .A2(n714), .ZN(n677) );
  NOR2_X1 U676 ( .A1(G2084), .A2(n680), .ZN(n676) );
  XOR2_X1 U677 ( .A(KEYINPUT103), .B(n612), .Z(n613) );
  NAND2_X1 U678 ( .A1(G8), .A2(n613), .ZN(n614) );
  XNOR2_X1 U679 ( .A(KEYINPUT30), .B(n614), .ZN(n615) );
  NOR2_X1 U680 ( .A1(n615), .A2(G168), .ZN(n616) );
  XNOR2_X1 U681 ( .A(n616), .B(KEYINPUT104), .ZN(n621) );
  NOR2_X1 U682 ( .A1(n655), .A2(G1961), .ZN(n617) );
  XNOR2_X1 U683 ( .A(n617), .B(KEYINPUT99), .ZN(n619) );
  XOR2_X1 U684 ( .A(n680), .B(KEYINPUT100), .Z(n662) );
  XNOR2_X1 U685 ( .A(G2078), .B(KEYINPUT25), .ZN(n966) );
  NAND2_X1 U686 ( .A1(n662), .A2(n966), .ZN(n618) );
  NAND2_X1 U687 ( .A1(n619), .A2(n618), .ZN(n624) );
  NOR2_X1 U688 ( .A1(n624), .A2(G171), .ZN(n620) );
  AND2_X1 U689 ( .A1(n624), .A2(G171), .ZN(n625) );
  XNOR2_X1 U690 ( .A(n625), .B(KEYINPUT101), .ZN(n675) );
  INV_X1 U691 ( .A(G299), .ZN(n632) );
  NAND2_X1 U692 ( .A1(G2072), .A2(n662), .ZN(n626) );
  XNOR2_X1 U693 ( .A(n626), .B(KEYINPUT27), .ZN(n628) );
  INV_X1 U694 ( .A(G1956), .ZN(n1011) );
  NOR2_X1 U695 ( .A1(n662), .A2(n1011), .ZN(n627) );
  NOR2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n631) );
  NOR2_X1 U697 ( .A1(n632), .A2(n631), .ZN(n630) );
  XNOR2_X1 U698 ( .A(n630), .B(n629), .ZN(n672) );
  NAND2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n670) );
  NAND2_X1 U700 ( .A1(G79), .A2(n816), .ZN(n633) );
  XNOR2_X1 U701 ( .A(n633), .B(KEYINPUT76), .ZN(n640) );
  NAND2_X1 U702 ( .A1(G54), .A2(n811), .ZN(n635) );
  NAND2_X1 U703 ( .A1(G66), .A2(n812), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U705 ( .A1(G92), .A2(n815), .ZN(n636) );
  XNOR2_X1 U706 ( .A(KEYINPUT75), .B(n636), .ZN(n637) );
  NOR2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U709 ( .A(KEYINPUT15), .B(n641), .Z(n884) );
  INV_X1 U710 ( .A(n884), .ZN(n987) );
  XOR2_X1 U711 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n643) );
  NAND2_X1 U712 ( .A1(G56), .A2(n812), .ZN(n642) );
  XNOR2_X1 U713 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n644), .B(KEYINPUT70), .ZN(n651) );
  XNOR2_X1 U715 ( .A(KEYINPUT72), .B(KEYINPUT13), .ZN(n649) );
  NAND2_X1 U716 ( .A1(n815), .A2(G81), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(KEYINPUT12), .ZN(n647) );
  NAND2_X1 U718 ( .A1(G68), .A2(n816), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n652), .B(KEYINPUT73), .ZN(n654) );
  NAND2_X1 U723 ( .A1(G43), .A2(n811), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n1001) );
  NAND2_X1 U725 ( .A1(G1996), .A2(n655), .ZN(n656) );
  XNOR2_X1 U726 ( .A(KEYINPUT26), .B(n656), .ZN(n659) );
  NAND2_X1 U727 ( .A1(n680), .A2(G1341), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n657), .B(KEYINPUT102), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U730 ( .A1(n1001), .A2(n660), .ZN(n661) );
  OR2_X1 U731 ( .A1(n987), .A2(n661), .ZN(n668) );
  NAND2_X1 U732 ( .A1(n987), .A2(n661), .ZN(n666) );
  NAND2_X1 U733 ( .A1(G2067), .A2(n662), .ZN(n664) );
  NAND2_X1 U734 ( .A1(G1348), .A2(n680), .ZN(n663) );
  NAND2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U740 ( .A(n673), .B(KEYINPUT29), .Z(n674) );
  NAND2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n684) );
  NAND2_X1 U742 ( .A1(n685), .A2(n684), .ZN(n679) );
  AND2_X1 U743 ( .A1(G8), .A2(n676), .ZN(n678) );
  NAND2_X1 U744 ( .A1(n679), .A2(n527), .ZN(n703) );
  NOR2_X1 U745 ( .A1(G1971), .A2(n714), .ZN(n682) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n680), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n683), .A2(G303), .ZN(n687) );
  AND2_X1 U749 ( .A1(n684), .A2(n687), .ZN(n686) );
  NAND2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n691) );
  INV_X1 U751 ( .A(n687), .ZN(n688) );
  OR2_X1 U752 ( .A1(n688), .A2(G286), .ZN(n689) );
  AND2_X1 U753 ( .A1(G8), .A2(n689), .ZN(n690) );
  NAND2_X1 U754 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U755 ( .A(n692), .B(KEYINPUT32), .ZN(n705) );
  NAND2_X1 U756 ( .A1(n703), .A2(n705), .ZN(n695) );
  NOR2_X1 U757 ( .A1(G2090), .A2(G303), .ZN(n693) );
  NAND2_X1 U758 ( .A1(G8), .A2(n693), .ZN(n694) );
  NAND2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U760 ( .A(n696), .B(KEYINPUT106), .ZN(n697) );
  AND2_X1 U761 ( .A1(n697), .A2(n714), .ZN(n701) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n698) );
  XOR2_X1 U763 ( .A(n698), .B(KEYINPUT24), .Z(n699) );
  NOR2_X1 U764 ( .A1(n714), .A2(n699), .ZN(n700) );
  NOR2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n722) );
  AND2_X1 U766 ( .A1(G1976), .A2(G288), .ZN(n994) );
  OR2_X1 U767 ( .A1(n994), .A2(n714), .ZN(n707) );
  INV_X1 U768 ( .A(n707), .ZN(n702) );
  AND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  AND2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n711) );
  NOR2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n712) );
  NOR2_X1 U772 ( .A1(G303), .A2(G1971), .ZN(n706) );
  NOR2_X1 U773 ( .A1(n712), .A2(n706), .ZN(n996) );
  OR2_X1 U774 ( .A1(n707), .A2(n996), .ZN(n709) );
  INV_X1 U775 ( .A(KEYINPUT33), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n710) );
  OR2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n718) );
  XOR2_X1 U778 ( .A(G1981), .B(G305), .Z(n984) );
  NAND2_X1 U779 ( .A1(n712), .A2(KEYINPUT33), .ZN(n713) );
  NOR2_X1 U780 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n720) );
  NAND2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n724) );
  INV_X1 U783 ( .A(KEYINPUT107), .ZN(n723) );
  XNOR2_X1 U784 ( .A(n724), .B(n723), .ZN(n760) );
  XNOR2_X1 U785 ( .A(G1986), .B(G290), .ZN(n993) );
  NOR2_X1 U786 ( .A1(n726), .A2(n725), .ZN(n773) );
  NAND2_X1 U787 ( .A1(n993), .A2(n773), .ZN(n758) );
  NAND2_X1 U788 ( .A1(G107), .A2(n916), .ZN(n728) );
  NAND2_X1 U789 ( .A1(G95), .A2(n912), .ZN(n727) );
  NAND2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n734) );
  BUF_X1 U791 ( .A(n729), .Z(n917) );
  NAND2_X1 U792 ( .A1(G119), .A2(n917), .ZN(n730) );
  XNOR2_X1 U793 ( .A(n730), .B(KEYINPUT96), .ZN(n732) );
  NAND2_X1 U794 ( .A1(G131), .A2(n913), .ZN(n731) );
  NAND2_X1 U795 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U796 ( .A1(n734), .A2(n733), .ZN(n895) );
  INV_X1 U797 ( .A(G1991), .ZN(n762) );
  NOR2_X1 U798 ( .A1(n895), .A2(n762), .ZN(n744) );
  NAND2_X1 U799 ( .A1(n913), .A2(G141), .ZN(n741) );
  NAND2_X1 U800 ( .A1(G117), .A2(n916), .ZN(n736) );
  NAND2_X1 U801 ( .A1(G129), .A2(n917), .ZN(n735) );
  NAND2_X1 U802 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U803 ( .A1(n912), .A2(G105), .ZN(n737) );
  XOR2_X1 U804 ( .A(KEYINPUT38), .B(n737), .Z(n738) );
  NOR2_X1 U805 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U806 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U807 ( .A(KEYINPUT97), .B(n742), .ZN(n896) );
  INV_X1 U808 ( .A(G1996), .ZN(n860) );
  NOR2_X1 U809 ( .A1(n896), .A2(n860), .ZN(n743) );
  NOR2_X1 U810 ( .A1(n744), .A2(n743), .ZN(n943) );
  INV_X1 U811 ( .A(n943), .ZN(n745) );
  NAND2_X1 U812 ( .A1(n745), .A2(n773), .ZN(n761) );
  NAND2_X1 U813 ( .A1(G104), .A2(n912), .ZN(n747) );
  NAND2_X1 U814 ( .A1(G140), .A2(n913), .ZN(n746) );
  NAND2_X1 U815 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U816 ( .A(KEYINPUT34), .B(n748), .ZN(n753) );
  NAND2_X1 U817 ( .A1(G116), .A2(n916), .ZN(n750) );
  NAND2_X1 U818 ( .A1(G128), .A2(n917), .ZN(n749) );
  NAND2_X1 U819 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U820 ( .A(n751), .B(KEYINPUT35), .Z(n752) );
  NOR2_X1 U821 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U822 ( .A(KEYINPUT36), .B(n754), .Z(n755) );
  XNOR2_X1 U823 ( .A(KEYINPUT95), .B(n755), .ZN(n925) );
  XNOR2_X1 U824 ( .A(KEYINPUT37), .B(G2067), .ZN(n771) );
  NOR2_X1 U825 ( .A1(n925), .A2(n771), .ZN(n957) );
  NAND2_X1 U826 ( .A1(n773), .A2(n957), .ZN(n769) );
  NAND2_X1 U827 ( .A1(n761), .A2(n769), .ZN(n756) );
  XOR2_X1 U828 ( .A(n756), .B(KEYINPUT98), .Z(n757) );
  AND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U830 ( .A1(n760), .A2(n759), .ZN(n776) );
  AND2_X1 U831 ( .A1(n860), .A2(n896), .ZN(n949) );
  INV_X1 U832 ( .A(n761), .ZN(n765) );
  AND2_X1 U833 ( .A1(n762), .A2(n895), .ZN(n945) );
  NOR2_X1 U834 ( .A1(G1986), .A2(G290), .ZN(n763) );
  NOR2_X1 U835 ( .A1(n945), .A2(n763), .ZN(n764) );
  NOR2_X1 U836 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U837 ( .A(n766), .B(KEYINPUT108), .ZN(n767) );
  NOR2_X1 U838 ( .A1(n949), .A2(n767), .ZN(n768) );
  XNOR2_X1 U839 ( .A(n768), .B(KEYINPUT39), .ZN(n770) );
  NAND2_X1 U840 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U841 ( .A1(n925), .A2(n771), .ZN(n954) );
  NAND2_X1 U842 ( .A1(n772), .A2(n954), .ZN(n774) );
  NAND2_X1 U843 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U844 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U845 ( .A(n777), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U846 ( .A(G2443), .B(G2446), .Z(n779) );
  XNOR2_X1 U847 ( .A(G2427), .B(G2451), .ZN(n778) );
  XNOR2_X1 U848 ( .A(n779), .B(n778), .ZN(n785) );
  XOR2_X1 U849 ( .A(G2430), .B(G2454), .Z(n781) );
  XNOR2_X1 U850 ( .A(G1341), .B(G1348), .ZN(n780) );
  XNOR2_X1 U851 ( .A(n781), .B(n780), .ZN(n783) );
  XOR2_X1 U852 ( .A(G2435), .B(G2438), .Z(n782) );
  XNOR2_X1 U853 ( .A(n783), .B(n782), .ZN(n784) );
  XOR2_X1 U854 ( .A(n785), .B(n784), .Z(n786) );
  AND2_X1 U855 ( .A1(G14), .A2(n786), .ZN(G401) );
  AND2_X1 U856 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U857 ( .A(G132), .ZN(G219) );
  INV_X1 U858 ( .A(G82), .ZN(G220) );
  INV_X1 U859 ( .A(G57), .ZN(G237) );
  INV_X1 U860 ( .A(G120), .ZN(G236) );
  NAND2_X1 U861 ( .A1(G7), .A2(G661), .ZN(n787) );
  XOR2_X1 U862 ( .A(n787), .B(KEYINPUT10), .Z(n851) );
  NAND2_X1 U863 ( .A1(n851), .A2(G567), .ZN(n788) );
  XOR2_X1 U864 ( .A(KEYINPUT11), .B(n788), .Z(G234) );
  XOR2_X1 U865 ( .A(G860), .B(KEYINPUT74), .Z(n793) );
  OR2_X1 U866 ( .A1(n793), .A2(n1001), .ZN(G153) );
  INV_X1 U867 ( .A(G171), .ZN(G301) );
  NAND2_X1 U868 ( .A1(G868), .A2(G301), .ZN(n790) );
  INV_X1 U869 ( .A(G868), .ZN(n797) );
  NAND2_X1 U870 ( .A1(n884), .A2(n797), .ZN(n789) );
  NAND2_X1 U871 ( .A1(n790), .A2(n789), .ZN(G284) );
  NOR2_X1 U872 ( .A1(G286), .A2(n797), .ZN(n792) );
  NOR2_X1 U873 ( .A1(G868), .A2(G299), .ZN(n791) );
  NOR2_X1 U874 ( .A1(n792), .A2(n791), .ZN(G297) );
  NAND2_X1 U875 ( .A1(n793), .A2(G559), .ZN(n794) );
  NAND2_X1 U876 ( .A1(n794), .A2(n987), .ZN(n795) );
  XNOR2_X1 U877 ( .A(n795), .B(KEYINPUT79), .ZN(n796) );
  XOR2_X1 U878 ( .A(KEYINPUT16), .B(n796), .Z(G148) );
  NOR2_X1 U879 ( .A1(n884), .A2(n797), .ZN(n798) );
  XOR2_X1 U880 ( .A(KEYINPUT80), .B(n798), .Z(n799) );
  NOR2_X1 U881 ( .A1(G559), .A2(n799), .ZN(n801) );
  NOR2_X1 U882 ( .A1(G868), .A2(n1001), .ZN(n800) );
  NOR2_X1 U883 ( .A1(n801), .A2(n800), .ZN(G282) );
  NAND2_X1 U884 ( .A1(G111), .A2(n916), .ZN(n803) );
  NAND2_X1 U885 ( .A1(G99), .A2(n912), .ZN(n802) );
  NAND2_X1 U886 ( .A1(n803), .A2(n802), .ZN(n808) );
  NAND2_X1 U887 ( .A1(G123), .A2(n917), .ZN(n804) );
  XNOR2_X1 U888 ( .A(n804), .B(KEYINPUT18), .ZN(n806) );
  NAND2_X1 U889 ( .A1(G135), .A2(n913), .ZN(n805) );
  NAND2_X1 U890 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U891 ( .A1(n808), .A2(n807), .ZN(n941) );
  XNOR2_X1 U892 ( .A(G2096), .B(n941), .ZN(n809) );
  INV_X1 U893 ( .A(G2100), .ZN(n874) );
  NAND2_X1 U894 ( .A1(n809), .A2(n874), .ZN(G156) );
  NAND2_X1 U895 ( .A1(n987), .A2(G559), .ZN(n833) );
  XNOR2_X1 U896 ( .A(n1001), .B(n833), .ZN(n810) );
  NOR2_X1 U897 ( .A1(n810), .A2(G860), .ZN(n821) );
  NAND2_X1 U898 ( .A1(G55), .A2(n811), .ZN(n814) );
  NAND2_X1 U899 ( .A1(G67), .A2(n812), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n814), .A2(n813), .ZN(n820) );
  NAND2_X1 U901 ( .A1(G93), .A2(n815), .ZN(n818) );
  NAND2_X1 U902 ( .A1(G80), .A2(n816), .ZN(n817) );
  NAND2_X1 U903 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U904 ( .A1(n820), .A2(n819), .ZN(n826) );
  XNOR2_X1 U905 ( .A(n821), .B(n826), .ZN(G145) );
  NOR2_X1 U906 ( .A1(G868), .A2(n826), .ZN(n822) );
  XOR2_X1 U907 ( .A(n822), .B(KEYINPUT90), .Z(n836) );
  XOR2_X1 U908 ( .A(G166), .B(n1001), .Z(n832) );
  XOR2_X1 U909 ( .A(KEYINPUT89), .B(KEYINPUT19), .Z(n824) );
  XNOR2_X1 U910 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n823) );
  XNOR2_X1 U911 ( .A(n824), .B(n823), .ZN(n825) );
  XNOR2_X1 U912 ( .A(n826), .B(n825), .ZN(n828) );
  XOR2_X1 U913 ( .A(G290), .B(G299), .Z(n827) );
  XNOR2_X1 U914 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U915 ( .A(n829), .B(G305), .Z(n830) );
  XNOR2_X1 U916 ( .A(G288), .B(n830), .ZN(n831) );
  XNOR2_X1 U917 ( .A(n832), .B(n831), .ZN(n881) );
  XOR2_X1 U918 ( .A(n881), .B(n833), .Z(n834) );
  NAND2_X1 U919 ( .A1(G868), .A2(n834), .ZN(n835) );
  NAND2_X1 U920 ( .A1(n836), .A2(n835), .ZN(G295) );
  NAND2_X1 U921 ( .A1(G2078), .A2(G2084), .ZN(n837) );
  XOR2_X1 U922 ( .A(KEYINPUT20), .B(n837), .Z(n838) );
  NAND2_X1 U923 ( .A1(G2090), .A2(n838), .ZN(n839) );
  XNOR2_X1 U924 ( .A(KEYINPUT21), .B(n839), .ZN(n840) );
  NAND2_X1 U925 ( .A1(n840), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U926 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U927 ( .A1(G236), .A2(G237), .ZN(n841) );
  NAND2_X1 U928 ( .A1(G69), .A2(n841), .ZN(n842) );
  XNOR2_X1 U929 ( .A(KEYINPUT91), .B(n842), .ZN(n843) );
  NAND2_X1 U930 ( .A1(n843), .A2(G108), .ZN(n855) );
  NAND2_X1 U931 ( .A1(G567), .A2(n855), .ZN(n848) );
  NOR2_X1 U932 ( .A1(G220), .A2(G219), .ZN(n844) );
  XOR2_X1 U933 ( .A(KEYINPUT22), .B(n844), .Z(n845) );
  NOR2_X1 U934 ( .A1(G218), .A2(n845), .ZN(n846) );
  NAND2_X1 U935 ( .A1(G96), .A2(n846), .ZN(n856) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n856), .ZN(n847) );
  NAND2_X1 U937 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U938 ( .A(KEYINPUT92), .B(n849), .ZN(n929) );
  NAND2_X1 U939 ( .A1(G661), .A2(G483), .ZN(n850) );
  NOR2_X1 U940 ( .A1(n929), .A2(n850), .ZN(n854) );
  NAND2_X1 U941 ( .A1(n854), .A2(G36), .ZN(G176) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n851), .ZN(G217) );
  INV_X1 U943 ( .A(n851), .ZN(G223) );
  AND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n852) );
  NAND2_X1 U945 ( .A1(G661), .A2(n852), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n853) );
  NAND2_X1 U947 ( .A1(n854), .A2(n853), .ZN(G188) );
  INV_X1 U949 ( .A(G108), .ZN(G238) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  NOR2_X1 U951 ( .A1(n856), .A2(n855), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  XOR2_X1 U953 ( .A(KEYINPUT114), .B(G1981), .Z(n858) );
  XOR2_X1 U954 ( .A(G1986), .B(n1011), .Z(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U956 ( .A(n859), .B(KEYINPUT113), .Z(n862) );
  XOR2_X1 U957 ( .A(n860), .B(G1991), .Z(n861) );
  XNOR2_X1 U958 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U959 ( .A(G1976), .B(G1971), .Z(n864) );
  XNOR2_X1 U960 ( .A(G1966), .B(G1961), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U962 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U963 ( .A(G2474), .B(KEYINPUT41), .ZN(n867) );
  XNOR2_X1 U964 ( .A(n868), .B(n867), .ZN(G229) );
  XOR2_X1 U965 ( .A(KEYINPUT42), .B(KEYINPUT112), .Z(n870) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(G2096), .ZN(n869) );
  XNOR2_X1 U967 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U968 ( .A(n871), .B(KEYINPUT111), .Z(n873) );
  XNOR2_X1 U969 ( .A(G2072), .B(G2090), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n878) );
  XNOR2_X1 U971 ( .A(n874), .B(G2084), .ZN(n876) );
  XNOR2_X1 U972 ( .A(G2067), .B(G2078), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U974 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U975 ( .A(G2678), .B(KEYINPUT43), .ZN(n879) );
  XNOR2_X1 U976 ( .A(n880), .B(n879), .ZN(G227) );
  XOR2_X1 U977 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n883) );
  XOR2_X1 U978 ( .A(G301), .B(n881), .Z(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n886) );
  XOR2_X1 U980 ( .A(G286), .B(n884), .Z(n885) );
  XNOR2_X1 U981 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U982 ( .A1(G37), .A2(n887), .ZN(G397) );
  NAND2_X1 U983 ( .A1(G112), .A2(n916), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G100), .A2(n912), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n894) );
  NAND2_X1 U986 ( .A1(G124), .A2(n917), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n890), .B(KEYINPUT44), .ZN(n892) );
  NAND2_X1 U988 ( .A1(G136), .A2(n913), .ZN(n891) );
  NAND2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n893) );
  NOR2_X1 U990 ( .A1(n894), .A2(n893), .ZN(G162) );
  XNOR2_X1 U991 ( .A(n895), .B(n941), .ZN(n898) );
  XNOR2_X1 U992 ( .A(G164), .B(n896), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n911) );
  XOR2_X1 U994 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n909) );
  NAND2_X1 U995 ( .A1(G106), .A2(n912), .ZN(n900) );
  NAND2_X1 U996 ( .A1(G142), .A2(n913), .ZN(n899) );
  NAND2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n901), .B(KEYINPUT45), .ZN(n903) );
  NAND2_X1 U999 ( .A1(G130), .A2(n917), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n906) );
  NAND2_X1 U1001 ( .A1(G118), .A2(n916), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(KEYINPUT115), .B(n904), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(G162), .B(n907), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(n911), .B(n910), .Z(n924) );
  NAND2_X1 U1007 ( .A1(G103), .A2(n912), .ZN(n915) );
  NAND2_X1 U1008 ( .A1(G139), .A2(n913), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(n915), .A2(n914), .ZN(n922) );
  NAND2_X1 U1010 ( .A1(G115), .A2(n916), .ZN(n919) );
  NAND2_X1 U1011 ( .A1(G127), .A2(n917), .ZN(n918) );
  NAND2_X1 U1012 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1013 ( .A(KEYINPUT47), .B(n920), .Z(n921) );
  NOR2_X1 U1014 ( .A1(n922), .A2(n921), .ZN(n935) );
  XNOR2_X1 U1015 ( .A(G160), .B(n935), .ZN(n923) );
  XNOR2_X1 U1016 ( .A(n924), .B(n923), .ZN(n926) );
  XNOR2_X1 U1017 ( .A(n926), .B(n925), .ZN(n927) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n927), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(KEYINPUT116), .B(n928), .ZN(G395) );
  XNOR2_X1 U1020 ( .A(KEYINPUT109), .B(n929), .ZN(G319) );
  NOR2_X1 U1021 ( .A1(G229), .A2(G227), .ZN(n930) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n930), .ZN(n931) );
  NOR2_X1 U1023 ( .A1(G401), .A2(n931), .ZN(n933) );
  NOR2_X1 U1024 ( .A1(G397), .A2(G395), .ZN(n932) );
  AND2_X1 U1025 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1026 ( .A1(n934), .A2(G319), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(KEYINPUT121), .ZN(n959) );
  XOR2_X1 U1030 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1031 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(KEYINPUT50), .B(n938), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(n939), .B(KEYINPUT120), .ZN(n947) );
  XOR2_X1 U1035 ( .A(G2084), .B(G160), .Z(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n953) );
  XOR2_X1 U1040 ( .A(G2090), .B(G162), .Z(n948) );
  NOR2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1042 ( .A(KEYINPUT119), .B(n950), .Z(n951) );
  XNOR2_X1 U1043 ( .A(n951), .B(KEYINPUT51), .ZN(n952) );
  NOR2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1045 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1046 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1047 ( .A(n959), .B(n958), .ZN(n960) );
  OR2_X1 U1048 ( .A1(KEYINPUT55), .A2(n960), .ZN(n961) );
  NAND2_X1 U1049 ( .A1(n961), .A2(G29), .ZN(n962) );
  XNOR2_X1 U1050 ( .A(n962), .B(KEYINPUT122), .ZN(n1039) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G26), .ZN(n964) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n963) );
  NOR2_X1 U1053 ( .A1(n964), .A2(n963), .ZN(n972) );
  XOR2_X1 U1054 ( .A(G25), .B(G1991), .Z(n965) );
  NAND2_X1 U1055 ( .A1(n965), .A2(G28), .ZN(n970) );
  XNOR2_X1 U1056 ( .A(n966), .B(G27), .ZN(n968) );
  XOR2_X1 U1057 ( .A(G1996), .B(G32), .Z(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1059 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1060 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(n973), .B(KEYINPUT53), .ZN(n976) );
  XOR2_X1 U1062 ( .A(G2084), .B(G34), .Z(n974) );
  XNOR2_X1 U1063 ( .A(KEYINPUT54), .B(n974), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(n976), .A2(n975), .ZN(n979) );
  XOR2_X1 U1065 ( .A(KEYINPUT123), .B(G2090), .Z(n977) );
  XNOR2_X1 U1066 ( .A(G35), .B(n977), .ZN(n978) );
  NOR2_X1 U1067 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(KEYINPUT55), .B(n980), .ZN(n982) );
  INV_X1 U1069 ( .A(G29), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1071 ( .A1(n983), .A2(G11), .ZN(n1037) );
  INV_X1 U1072 ( .A(G16), .ZN(n1033) );
  XOR2_X1 U1073 ( .A(n1033), .B(KEYINPUT56), .Z(n1007) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G168), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(n986), .B(KEYINPUT57), .ZN(n1005) );
  XOR2_X1 U1077 ( .A(G171), .B(G1961), .Z(n989) );
  XOR2_X1 U1078 ( .A(n987), .B(G1348), .Z(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(KEYINPUT124), .B(n990), .ZN(n1000) );
  XOR2_X1 U1081 ( .A(G299), .B(G1956), .Z(n992) );
  NAND2_X1 U1082 ( .A1(G1971), .A2(G303), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n998) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XNOR2_X1 U1088 ( .A(G1341), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1090 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1091 ( .A1(n1007), .A2(n1006), .ZN(n1035) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1009) );
  XNOR2_X1 U1093 ( .A(G5), .B(G1961), .ZN(n1008) );
  NOR2_X1 U1094 ( .A1(n1009), .A2(n1008), .ZN(n1021) );
  XNOR2_X1 U1095 ( .A(KEYINPUT59), .B(G1348), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(n1010), .B(G4), .ZN(n1018) );
  XOR2_X1 U1097 ( .A(n1011), .B(G20), .Z(n1016) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(G6), .B(G1981), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT125), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1019), .Z(n1020) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1030) );
  XOR2_X1 U1106 ( .A(G1986), .B(G24), .Z(n1026) );
  XNOR2_X1 U1107 ( .A(G1971), .B(G22), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(G1976), .B(G23), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(n1024), .B(KEYINPUT126), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1027), .Z(n1028) );
  XNOR2_X1 U1113 ( .A(KEYINPUT58), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(KEYINPUT61), .B(n1031), .ZN(n1032) );
  NAND2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1117 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1118 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1119 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1040), .ZN(G150) );
  INV_X1 U1121 ( .A(G150), .ZN(G311) );
endmodule

