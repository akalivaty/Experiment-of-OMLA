//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT65), .Z(new_n214));
  AOI22_X1  g0014(.A1(new_n208), .A2(new_n209), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n215), .B1(new_n209), .B2(new_n208), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT66), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(KEYINPUT66), .B1(new_n217), .B2(new_n218), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n216), .A2(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XNOR2_X1  g0034(.A(G50), .B(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G58), .B(G77), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(G97), .B(G107), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  INV_X1    g0041(.A(G33), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G232), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G226), .A3(new_n247), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G97), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT13), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G274), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n254), .A2(new_n259), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(G238), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n255), .A2(new_n256), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n256), .B1(new_n255), .B2(new_n263), .ZN(new_n265));
  OAI21_X1  g0065(.A(G200), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n255), .A2(new_n263), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT13), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n255), .A2(new_n256), .A3(new_n263), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G190), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G68), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT12), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n211), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n278), .A2(G77), .B1(G20), .B2(new_n274), .ZN(new_n279));
  INV_X1    g0079(.A(G50), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n210), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n285), .B1(new_n271), .B2(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n276), .B(new_n286), .C1(new_n274), .C2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT11), .B1(new_n283), .B2(new_n285), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n266), .A2(new_n270), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(G169), .B1(new_n264), .B2(new_n265), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT14), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT14), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(G169), .C1(new_n264), .C2(new_n265), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n264), .A2(new_n265), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G179), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n294), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n291), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n292), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT73), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G1), .A3(G13), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(G232), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n260), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n243), .A2(new_n245), .A3(G226), .A4(G1698), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n243), .A2(new_n245), .A3(G223), .A4(new_n247), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G87), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI211_X1 g0112(.A(G190), .B(new_n308), .C1(new_n254), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n254), .ZN(new_n314));
  INV_X1    g0114(.A(new_n308), .ZN(new_n315));
  AOI21_X1  g0115(.A(G200), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n303), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT8), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT68), .B1(new_n318), .B2(G58), .ZN(new_n319));
  INV_X1    g0119(.A(G58), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(KEYINPUT8), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(KEYINPUT68), .A3(G58), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n288), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n323), .B2(new_n273), .ZN(new_n325));
  INV_X1    g0125(.A(G190), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n314), .A2(new_n326), .A3(new_n315), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n308), .B1(new_n312), .B2(new_n254), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n327), .B(KEYINPUT73), .C1(G200), .C2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT7), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n250), .A2(new_n330), .A3(G20), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT7), .B1(new_n246), .B2(new_n211), .ZN(new_n332));
  OAI21_X1  g0132(.A(G68), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n320), .A2(new_n274), .ZN(new_n334));
  NOR2_X1   g0134(.A1(G58), .A2(G68), .ZN(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n281), .A2(G159), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n333), .A2(KEYINPUT16), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT16), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n330), .B1(new_n250), .B2(G20), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n246), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n274), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n341), .B1(new_n344), .B2(new_n338), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(new_n345), .A3(new_n285), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n317), .A2(new_n325), .A3(new_n329), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT17), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n346), .A2(new_n325), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT17), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(new_n329), .A4(new_n317), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n346), .A2(new_n325), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n328), .A2(G179), .ZN(new_n353));
  INV_X1    g0153(.A(G169), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(new_n328), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT18), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(KEYINPUT18), .A3(new_n355), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n348), .A2(new_n351), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n362));
  OR2_X1    g0162(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n272), .A2(G50), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n287), .B2(G50), .ZN(new_n365));
  INV_X1    g0165(.A(G150), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n366), .A2(new_n282), .B1(new_n201), .B2(new_n211), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n323), .B2(new_n278), .ZN(new_n368));
  INV_X1    g0168(.A(new_n285), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT9), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT9), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n365), .C1(new_n368), .C2(new_n369), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n261), .B1(new_n262), .B2(G226), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n250), .A2(G222), .A3(new_n247), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n250), .A2(G223), .A3(G1698), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n246), .A2(G77), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT67), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n305), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT67), .A4(new_n379), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n376), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G190), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n374), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G200), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n362), .B(new_n363), .C1(new_n386), .C2(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n371), .A2(new_n373), .B1(new_n384), .B2(G190), .ZN(new_n390));
  INV_X1    g0190(.A(new_n388), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT72), .A4(KEYINPUT10), .ZN(new_n392));
  INV_X1    g0192(.A(G179), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n384), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(new_n370), .C1(G169), .C2(new_n384), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n389), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n248), .A2(G238), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n250), .A2(G232), .A3(new_n247), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n246), .A2(G107), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n254), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n261), .B1(new_n262), .B2(G244), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n393), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT71), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT71), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n401), .A2(new_n405), .A3(new_n393), .A4(new_n402), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n402), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n354), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT8), .B(G58), .ZN(new_n410));
  XOR2_X1   g0210(.A(new_n410), .B(KEYINPUT69), .Z(new_n411));
  OAI22_X1  g0211(.A1(new_n411), .A2(new_n282), .B1(new_n211), .B2(new_n202), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT70), .ZN(new_n413));
  XOR2_X1   g0213(.A(KEYINPUT15), .B(G87), .Z(new_n414));
  AOI22_X1  g0214(.A1(new_n412), .A2(new_n413), .B1(new_n278), .B2(new_n414), .ZN(new_n415));
  OAI221_X1 g0215(.A(KEYINPUT70), .B1(new_n211), .B2(new_n202), .C1(new_n411), .C2(new_n282), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n369), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n272), .A2(G77), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n287), .B2(G77), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n407), .B(new_n409), .C1(new_n417), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n412), .A2(new_n413), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n414), .A2(new_n278), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n416), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n285), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n408), .A2(G200), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n401), .A2(G190), .A3(new_n402), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n425), .A2(new_n419), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  NOR4_X1   g0229(.A1(new_n302), .A2(new_n361), .A3(new_n396), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT21), .ZN(new_n431));
  INV_X1    g0231(.A(G116), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n273), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n271), .A2(G33), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n272), .A2(new_n434), .A3(new_n210), .A4(new_n284), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n433), .B1(new_n435), .B2(new_n432), .ZN(new_n436));
  AOI21_X1  g0236(.A(G20), .B1(G33), .B2(G283), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n242), .A2(G97), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n432), .A2(G20), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n285), .A2(KEYINPUT79), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT79), .B1(new_n285), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT20), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT80), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(KEYINPUT20), .B(new_n439), .C1(new_n441), .C2(new_n442), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(KEYINPUT80), .A3(new_n444), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n436), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT76), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT5), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(G41), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n257), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n258), .A2(G1), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n452), .A2(G41), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(G274), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n271), .B(G45), .C1(new_n257), .C2(KEYINPUT5), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n452), .A2(G41), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n305), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n459), .B1(new_n463), .B2(G270), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n243), .A2(new_n245), .A3(G264), .A4(G1698), .ZN(new_n465));
  INV_X1    g0265(.A(G303), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(new_n250), .ZN(new_n467));
  INV_X1    g0267(.A(G257), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n246), .A2(new_n468), .A3(G1698), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n254), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G169), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n431), .B1(new_n450), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(G200), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n450), .B(new_n474), .C1(new_n326), .C2(new_n471), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT80), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n285), .A2(new_n440), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n285), .A2(KEYINPUT79), .A3(new_n440), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n479), .A2(new_n480), .B1(new_n438), .B2(new_n437), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n476), .B1(new_n481), .B2(KEYINPUT20), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n449), .A3(new_n446), .ZN(new_n483));
  INV_X1    g0283(.A(new_n436), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n471), .A2(KEYINPUT21), .A3(G169), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n464), .A2(new_n470), .A3(G179), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n485), .B2(new_n488), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n473), .B(new_n475), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n243), .A2(new_n245), .A3(G250), .A4(new_n247), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n243), .A2(new_n245), .A3(G257), .A4(G1698), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G294), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n254), .ZN(new_n498));
  OAI211_X1 g0298(.A(G264), .B(new_n305), .C1(new_n460), .C2(new_n461), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT84), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT84), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n498), .A2(new_n502), .A3(new_n499), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n459), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n459), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n498), .A2(new_n505), .A3(new_n499), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n504), .A2(G200), .B1(G190), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n273), .A2(KEYINPUT25), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT25), .B1(new_n273), .B2(new_n508), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n510), .A2(new_n511), .B1(new_n508), .B2(new_n435), .ZN(new_n512));
  AND2_X1   g0312(.A1(KEYINPUT82), .A2(G87), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n250), .A2(new_n211), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT22), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT22), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n250), .A2(new_n516), .A3(new_n211), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT83), .B1(new_n508), .B2(G20), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT23), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI211_X1 g0321(.A(KEYINPUT83), .B(KEYINPUT23), .C1(new_n508), .C2(G20), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n521), .A2(new_n522), .B1(new_n432), .B2(new_n277), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT24), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n369), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n518), .A2(new_n524), .A3(KEYINPUT24), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n512), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n507), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n529), .ZN(new_n531));
  INV_X1    g0331(.A(new_n503), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n502), .B1(new_n498), .B2(new_n499), .ZN(new_n533));
  OAI211_X1 g0333(.A(G179), .B(new_n505), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n506), .A2(G169), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n243), .A2(new_n245), .A3(G244), .A4(G1698), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n243), .A2(new_n245), .A3(G238), .A4(new_n247), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G116), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n254), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n456), .A2(G274), .ZN(new_n543));
  OAI21_X1  g0343(.A(G250), .B1(new_n258), .B2(G1), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n254), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(G190), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT78), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n541), .B2(new_n254), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT78), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(G190), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n549), .A2(new_n387), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n414), .A2(new_n272), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n211), .B1(new_n252), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(G87), .ZN(new_n557));
  INV_X1    g0357(.A(G97), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(new_n508), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n243), .A2(new_n245), .A3(new_n211), .A4(G68), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n555), .B1(new_n277), .B2(new_n558), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n554), .B1(new_n563), .B2(new_n285), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n435), .A2(new_n557), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n553), .A2(new_n567), .ZN(new_n568));
  AOI211_X1 g0368(.A(G179), .B(new_n545), .C1(new_n541), .C2(new_n254), .ZN(new_n569));
  AOI21_X1  g0369(.A(G169), .B1(new_n542), .B2(new_n546), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n414), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n564), .B1(new_n572), .B2(new_n435), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n552), .A2(new_n568), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n530), .A2(new_n537), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT75), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT6), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n239), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n577), .A2(new_n558), .A3(G107), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(G20), .B1(G77), .B2(new_n281), .ZN(new_n582));
  OAI21_X1  g0382(.A(G107), .B1(new_n331), .B2(new_n332), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n369), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n435), .A2(G97), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT74), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n272), .A2(new_n558), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n586), .B1(new_n585), .B2(new_n587), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n576), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n590), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n588), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n579), .B1(new_n577), .B2(new_n239), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n595), .A2(new_n211), .B1(new_n202), .B2(new_n282), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n508), .B1(new_n342), .B2(new_n343), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n285), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n598), .A3(KEYINPUT75), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n462), .A2(new_n468), .B1(new_n458), .B2(new_n455), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n243), .A2(new_n245), .A3(G244), .A4(new_n247), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT4), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n247), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G283), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n250), .A2(G250), .A3(G1698), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n604), .A2(new_n605), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  AOI211_X1 g0408(.A(KEYINPUT77), .B(new_n601), .C1(new_n254), .C2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT77), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n254), .ZN(new_n611));
  INV_X1    g0411(.A(new_n601), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(G190), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n611), .A2(new_n612), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n600), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(KEYINPUT77), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n601), .B1(new_n608), .B2(new_n254), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n610), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n354), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n594), .A2(new_n598), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n619), .A2(new_n393), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n575), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n430), .A2(new_n493), .A3(new_n626), .ZN(G372));
  INV_X1    g0427(.A(KEYINPUT89), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n574), .A2(new_n622), .A3(new_n621), .A4(new_n623), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n624), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(KEYINPUT89), .A3(KEYINPUT26), .A4(new_n574), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT88), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n621), .A2(new_n623), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(new_n600), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n571), .A2(new_n573), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n542), .A2(new_n546), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT85), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(G200), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT85), .B1(new_n549), .B2(new_n387), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n554), .B(new_n565), .C1(new_n285), .C2(new_n563), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT86), .A4(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n552), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT86), .ZN(new_n647));
  INV_X1    g0447(.A(new_n642), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n644), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n639), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n592), .A2(new_n599), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n652), .A2(KEYINPUT88), .A3(new_n621), .A4(new_n623), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n637), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n630), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n634), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n530), .A2(new_n617), .A3(new_n624), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n646), .A2(new_n650), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n638), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT87), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n617), .A2(new_n624), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT87), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(new_n530), .A4(new_n651), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n485), .A2(new_n488), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n473), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n537), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n660), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n656), .A2(new_n667), .A3(new_n638), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n430), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT90), .Z(new_n670));
  NAND2_X1  g0470(.A1(new_n299), .A2(new_n300), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n421), .A2(KEYINPUT91), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n425), .A2(new_n419), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT91), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(new_n407), .A4(new_n409), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n671), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n292), .B1(new_n348), .B2(new_n351), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n676), .A2(new_n677), .B1(new_n358), .B2(new_n359), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n389), .A2(new_n392), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n395), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n670), .A2(new_n682), .ZN(G369));
  INV_X1    g0483(.A(new_n665), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n211), .A2(G13), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n271), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n450), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n684), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n492), .B2(new_n694), .ZN(new_n696));
  XNOR2_X1  g0496(.A(KEYINPUT92), .B(G330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n537), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n507), .A2(new_n529), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n529), .B2(new_n693), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n537), .B2(new_n693), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n473), .B1(new_n490), .B2(new_n491), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n706), .A2(new_n693), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n707), .A2(new_n702), .B1(new_n700), .B2(new_n693), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n705), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n207), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n559), .A2(G116), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n214), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n712), .ZN(new_n716));
  XOR2_X1   g0516(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n717));
  XNOR2_X1  g0517(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n668), .A2(new_n693), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT96), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n639), .B1(new_n634), .B2(new_n655), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n692), .B1(new_n723), .B2(new_n667), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT96), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n657), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n727), .B(new_n651), .C1(new_n706), .C2(new_n700), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n638), .B1(new_n629), .B2(KEYINPUT26), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n654), .B2(KEYINPUT26), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n728), .B1(new_n730), .B2(KEYINPUT97), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT97), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n732), .B(new_n729), .C1(KEYINPUT26), .C2(new_n654), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n693), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT98), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT98), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n736), .B(new_n693), .C1(new_n731), .C2(new_n733), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n735), .A2(KEYINPUT29), .A3(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT95), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n501), .A2(new_n503), .ZN(new_n740));
  AND4_X1   g0540(.A1(G179), .A2(new_n464), .A3(new_n549), .A4(new_n470), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n740), .B(new_n741), .C1(new_n609), .C2(new_n613), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n618), .A2(new_n620), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n464), .A2(new_n549), .A3(new_n470), .A4(G179), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n501), .B2(new_n503), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n745), .A2(new_n747), .A3(KEYINPUT95), .A4(KEYINPUT30), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  AND4_X1   g0549(.A1(new_n393), .A2(new_n615), .A3(new_n471), .A4(new_n640), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n505), .B1(new_n532), .B2(new_n533), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n742), .A2(new_n743), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n693), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n626), .A2(new_n493), .A3(new_n693), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(KEYINPUT31), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n742), .A2(new_n743), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n750), .A2(new_n751), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n759), .A2(KEYINPUT94), .B1(new_n744), .B2(new_n748), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n756), .B(new_n693), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n755), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n697), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n726), .A2(new_n738), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n718), .B1(new_n767), .B2(G1), .ZN(G364));
  AOI21_X1  g0568(.A(new_n271), .B1(new_n685), .B2(G45), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n712), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n699), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n697), .B2(new_n696), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n710), .A2(new_n246), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G355), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G116), .B2(new_n207), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n710), .A2(new_n250), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n258), .B2(new_n214), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n237), .A2(new_n258), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n211), .B1(KEYINPUT99), .B2(new_n354), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n354), .A2(KEYINPUT99), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n210), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n771), .B1(new_n781), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n211), .A2(new_n326), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n393), .A2(new_n387), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT100), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G179), .A2(G200), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n211), .B1(new_n800), .B2(G190), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n799), .A2(G326), .B1(G294), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n803), .A2(KEYINPUT102), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n211), .A2(G190), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n792), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(KEYINPUT33), .A2(G317), .ZN(new_n808));
  AND2_X1   g0608(.A1(KEYINPUT33), .A2(G317), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n393), .A2(G200), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n791), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G322), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n387), .A2(G179), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n805), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n810), .B(new_n814), .C1(new_n815), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n791), .A2(new_n816), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n805), .A2(new_n800), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G303), .A2(new_n820), .B1(new_n822), .B2(G329), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n811), .A2(new_n805), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n823), .B(new_n246), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n804), .A2(new_n818), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(KEYINPUT102), .B2(new_n803), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n801), .A2(new_n558), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G68), .B2(new_n807), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT101), .Z(new_n831));
  INV_X1    g0631(.A(new_n825), .ZN(new_n832));
  INV_X1    g0632(.A(new_n817), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G77), .A2(new_n832), .B1(new_n833), .B2(G107), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n834), .B1(new_n320), .B2(new_n812), .C1(new_n798), .C2(new_n280), .ZN(new_n835));
  INV_X1    g0635(.A(G159), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n821), .A2(KEYINPUT32), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n820), .A2(G87), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT32), .B1(new_n821), .B2(new_n836), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n838), .A2(new_n250), .A3(new_n839), .ZN(new_n840));
  OR3_X1    g0640(.A1(new_n835), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n828), .B1(new_n831), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n790), .B1(new_n842), .B2(new_n784), .ZN(new_n843));
  INV_X1    g0643(.A(new_n787), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n696), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n773), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G396));
  NAND2_X1  g0647(.A1(new_n721), .A2(new_n725), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n421), .A2(new_n428), .A3(KEYINPUT106), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n417), .A2(new_n420), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n693), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n849), .A2(new_n672), .A3(new_n675), .A4(new_n851), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n429), .A2(KEYINPUT106), .B1(new_n850), .B2(new_n693), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n692), .B(new_n854), .C1(new_n723), .C2(new_n667), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n771), .B1(new_n858), .B2(new_n766), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n766), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n784), .A2(new_n785), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(G77), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT104), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n246), .B1(new_n819), .B2(new_n508), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n799), .A2(G303), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(G294), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n812), .A2(new_n867), .B1(new_n825), .B2(new_n432), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(G311), .B2(new_n822), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n817), .A2(new_n557), .ZN(new_n870));
  XOR2_X1   g0670(.A(KEYINPUT103), .B(G283), .Z(new_n871));
  AOI211_X1 g0671(.A(new_n829), .B(new_n870), .C1(new_n807), .C2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n865), .A2(new_n864), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n866), .A2(new_n869), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  XOR2_X1   g0674(.A(KEYINPUT105), .B(G143), .Z(new_n875));
  AOI22_X1  g0675(.A1(new_n813), .A2(new_n875), .B1(new_n832), .B2(G159), .ZN(new_n876));
  INV_X1    g0676(.A(G137), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n876), .B1(new_n366), .B2(new_n806), .C1(new_n798), .C2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT34), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n250), .B1(new_n819), .B2(new_n280), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n833), .A2(G68), .ZN(new_n882));
  INV_X1    g0682(.A(G132), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(new_n821), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n881), .B(new_n884), .C1(G58), .C2(new_n802), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n878), .A2(new_n879), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n874), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n770), .B(new_n863), .C1(new_n888), .C2(new_n784), .ZN(new_n889));
  INV_X1    g0689(.A(new_n854), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n889), .B1(new_n890), .B2(new_n786), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n860), .A2(new_n891), .ZN(G384));
  OAI211_X1 g0692(.A(G116), .B(new_n212), .C1(new_n581), .C2(KEYINPUT35), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(KEYINPUT35), .B2(new_n581), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n214), .B(G77), .C1(new_n320), .C2(new_n274), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n280), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n271), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n352), .A2(new_n689), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n351), .A2(new_n348), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n358), .A2(new_n359), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n352), .B1(new_n355), .B2(new_n689), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n905), .A2(new_n906), .A3(new_n347), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(new_n905), .B2(new_n347), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n900), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n347), .ZN(new_n911));
  INV_X1    g0711(.A(new_n355), .ZN(new_n912));
  OAI211_X1 g0712(.A(KEYINPUT108), .B(new_n341), .C1(new_n344), .C2(new_n338), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n341), .A2(KEYINPUT108), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n333), .A2(new_n339), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n915), .A3(new_n285), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n912), .A2(new_n690), .B1(new_n325), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT37), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n905), .A2(new_n906), .A3(new_n347), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n325), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n689), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n920), .B(KEYINPUT38), .C1(new_n360), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n910), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n291), .A2(new_n693), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n293), .A2(KEYINPUT14), .B1(new_n297), .B2(G179), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n291), .B1(new_n927), .B2(new_n296), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n301), .A2(new_n926), .B1(new_n928), .B2(new_n692), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n854), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n749), .A2(new_n752), .ZN(new_n931));
  AND4_X1   g0731(.A1(KEYINPUT111), .A2(new_n931), .A3(KEYINPUT31), .A4(new_n692), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT111), .B1(new_n753), .B2(KEYINPUT31), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n924), .B(new_n930), .C1(new_n934), .C2(new_n755), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n928), .A2(new_n292), .A3(new_n925), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n671), .A2(new_n693), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n853), .B(new_n852), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT111), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n931), .A2(new_n692), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(new_n756), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n753), .A2(KEYINPUT111), .A3(KEYINPUT31), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR4_X1   g0743(.A1(new_n492), .A2(new_n575), .A3(new_n625), .A4(new_n692), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n940), .B1(new_n944), .B2(new_n756), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n938), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n922), .B1(new_n902), .B2(new_n903), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n921), .B1(new_n355), .B2(new_n689), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n906), .B1(new_n948), .B2(new_n347), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n907), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n900), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT40), .B1(new_n951), .B2(new_n923), .ZN(new_n952));
  AOI22_X1  g0752(.A1(KEYINPUT40), .A2(new_n935), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n430), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n945), .B2(new_n943), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n953), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n697), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n954), .B1(new_n726), .B2(new_n738), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n681), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n957), .B(new_n959), .Z(new_n960));
  INV_X1    g0760(.A(new_n929), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n951), .A2(new_n923), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n421), .A2(new_n692), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT107), .Z(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n961), .B(new_n962), .C1(new_n856), .C2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n671), .A2(new_n692), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT109), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n962), .A2(KEYINPUT39), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT39), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n910), .A2(new_n923), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n968), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n968), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n967), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n903), .A2(new_n689), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n966), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT110), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n960), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n271), .B2(new_n685), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n960), .A2(new_n979), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n899), .B1(new_n981), .B2(new_n982), .ZN(G367));
  XNOR2_X1  g0783(.A(new_n711), .B(KEYINPUT41), .ZN(new_n984));
  INV_X1    g0784(.A(new_n705), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n707), .A2(new_n702), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n704), .B2(new_n707), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n985), .B1(new_n987), .B2(new_n698), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n767), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n661), .B1(new_n600), .B2(new_n693), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n652), .A2(new_n621), .A3(new_n623), .A4(new_n692), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n708), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT45), .Z(new_n994));
  NOR2_X1   g0794(.A1(new_n708), .A2(new_n992), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT44), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n989), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n767), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n984), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n769), .B(KEYINPUT114), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n986), .A2(new_n990), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n992), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n624), .B1(new_n1007), .B2(new_n537), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n693), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n692), .A2(new_n567), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n639), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n659), .B2(new_n1012), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT112), .Z(new_n1015));
  INV_X1    g0815(.A(KEYINPUT43), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT113), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT113), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1011), .A2(new_n1020), .A3(new_n1017), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n705), .A2(new_n1007), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1019), .A2(new_n1016), .A3(new_n1015), .A4(new_n1021), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n705), .B2(new_n1007), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1004), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1015), .A2(new_n787), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n778), .A2(new_n233), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n789), .B1(new_n710), .B2(new_n414), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n770), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n812), .A2(new_n466), .B1(new_n817), .B2(new_n558), .ZN(new_n1035));
  INV_X1    g0835(.A(G317), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n806), .A2(new_n867), .B1(new_n821), .B2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1035), .B(new_n1037), .C1(new_n799), .C2(G311), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT46), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n819), .B2(new_n432), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n250), .B1(new_n832), .B2(new_n871), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n819), .A2(new_n1039), .A3(new_n432), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G107), .B2(new_n802), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n799), .A2(new_n875), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n802), .A2(G68), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n366), .A2(new_n812), .B1(new_n806), .B2(new_n836), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n817), .A2(new_n202), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1047), .A2(new_n246), .A3(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n825), .A2(new_n280), .B1(new_n821), .B2(new_n877), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G58), .B2(new_n820), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1045), .A2(new_n1046), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1044), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1054), .A2(KEYINPUT47), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n784), .B1(new_n1054), .B2(KEYINPUT47), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1031), .B(new_n1034), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1030), .A2(new_n1057), .ZN(G387));
  NOR2_X1   g0858(.A1(new_n704), .A2(new_n844), .ZN(new_n1059));
  AOI21_X1  g0859(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n411), .A2(G50), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n713), .B(new_n1060), .C1(new_n1061), .C2(KEYINPUT50), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(KEYINPUT50), .B2(new_n1061), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n778), .B1(new_n230), .B2(G45), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n713), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n774), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n508), .B2(new_n710), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n771), .B1(new_n1068), .B2(new_n789), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n799), .A2(G159), .B1(new_n323), .B2(new_n807), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n819), .A2(new_n202), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n812), .A2(new_n280), .B1(new_n821), .B2(new_n366), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G68), .C2(new_n832), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n572), .A2(new_n801), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n246), .B(new_n1074), .C1(G97), .C2(new_n833), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1070), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n822), .A2(G326), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n250), .B1(new_n833), .B2(G116), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n819), .A2(new_n867), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G317), .A2(new_n813), .B1(new_n832), .B2(G303), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n799), .A2(G322), .B1(G311), .B2(new_n807), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1082), .A2(KEYINPUT115), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(KEYINPUT115), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT48), .Z(new_n1086));
  AOI211_X1 g0886(.A(new_n1079), .B(new_n1086), .C1(new_n802), .C2(new_n871), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n1088));
  OAI211_X1 g0888(.A(new_n1077), .B(new_n1078), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1076), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1059), .B(new_n1069), .C1(new_n1091), .C2(new_n784), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n988), .B2(new_n1002), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n712), .B1(new_n767), .B2(new_n988), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n767), .B2(new_n988), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(G393));
  NOR2_X1   g0896(.A1(new_n999), .A2(new_n712), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n997), .B(new_n985), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n989), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n778), .A2(new_n240), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n788), .B1(new_n207), .B2(new_n558), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n771), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n798), .A2(new_n366), .B1(new_n836), .B2(new_n812), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT51), .Z(new_n1105));
  AOI22_X1  g0905(.A1(G68), .A2(new_n820), .B1(new_n822), .B2(new_n875), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n280), .B2(new_n806), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n801), .A2(new_n202), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1107), .A2(new_n246), .A3(new_n870), .A4(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n411), .B2(new_n825), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n798), .A2(new_n1036), .B1(new_n824), .B2(new_n812), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT52), .Z(new_n1112));
  AOI22_X1  g0912(.A1(new_n820), .A2(new_n871), .B1(new_n822), .B2(G322), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n246), .C1(new_n508), .C2(new_n817), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G303), .A2(new_n807), .B1(new_n832), .B2(G294), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n432), .B2(new_n801), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1114), .B1(KEYINPUT117), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(KEYINPUT117), .B2(new_n1116), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1105), .A2(new_n1110), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1103), .B1(new_n1119), .B2(new_n784), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n992), .B2(new_n844), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n1098), .B2(new_n1003), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1100), .A2(new_n1122), .ZN(G390));
  OAI21_X1  g0923(.A(new_n961), .B1(new_n856), .B2(new_n965), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n967), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n971), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n970), .B1(new_n951), .B2(new_n923), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT109), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n973), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1126), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n697), .B(new_n890), .C1(new_n755), .C2(new_n762), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1133), .A2(new_n929), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n943), .A2(new_n945), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(KEYINPUT118), .A3(G330), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n729), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n732), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n730), .A2(KEYINPUT97), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n728), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n736), .B1(new_n1143), .B2(new_n693), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n737), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n890), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n929), .B1(new_n1146), .B2(new_n964), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n924), .A2(new_n1125), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1132), .B(new_n1137), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n946), .A2(G330), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1150), .A2(KEYINPUT118), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1130), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n854), .B1(new_n735), .B2(new_n737), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n961), .B1(new_n1153), .B2(new_n965), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1148), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1149), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n955), .A2(G330), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n726), .A2(new_n738), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n682), .B(new_n1158), .C1(new_n1159), .C2(new_n954), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1153), .A2(new_n965), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1135), .A2(G330), .A3(new_n890), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1134), .B1(new_n1162), .B2(new_n929), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n857), .A2(new_n964), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1133), .A2(new_n929), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1150), .A2(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1161), .A2(new_n1163), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1160), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n712), .B1(new_n1157), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n1157), .B2(new_n1168), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n323), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n770), .B1(new_n1171), .B2(new_n861), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n784), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n822), .A2(G294), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n838), .A2(new_n882), .A3(new_n1174), .A4(new_n246), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(new_n1108), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G107), .A2(new_n807), .B1(new_n813), .B2(G116), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n558), .B2(new_n825), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G283), .B2(new_n799), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n250), .B1(new_n817), .B2(new_n280), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n819), .A2(new_n366), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT53), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1181), .A2(new_n1182), .B1(new_n836), .B2(new_n801), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1180), .B(new_n1183), .C1(new_n1182), .C2(new_n1181), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT54), .B(G143), .Z(new_n1185));
  AOI22_X1  g0985(.A1(new_n807), .A2(G137), .B1(new_n832), .B2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G132), .A2(new_n813), .B1(new_n822), .B2(G125), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n799), .B2(G128), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1176), .A2(new_n1179), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1172), .B1(new_n1173), .B2(new_n1190), .C1(new_n1130), .C2(new_n786), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1157), .B2(new_n1002), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1170), .A2(new_n1193), .ZN(G378));
  INV_X1    g0994(.A(new_n1149), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1151), .B1(new_n1196), .B2(new_n1132), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1168), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1158), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n958), .A2(new_n1199), .A3(new_n681), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT121), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT119), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n396), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n370), .A2(new_n689), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n389), .A2(new_n392), .A3(KEYINPUT119), .A4(new_n395), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1208), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1205), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1208), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1204), .A3(new_n1216), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1212), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n935), .A2(KEYINPUT40), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1135), .A2(new_n930), .A3(new_n952), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1219), .B1(new_n1222), .B2(G330), .ZN(new_n1223));
  INV_X1    g1023(.A(G330), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1224), .B(new_n1218), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n966), .A2(new_n975), .A3(new_n977), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1223), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1218), .B1(new_n953), .B2(new_n1224), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1222), .A2(G330), .A3(new_n1219), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n976), .B1(new_n1130), .B2(new_n967), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1228), .A2(new_n1229), .B1(new_n1230), .B2(new_n966), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1203), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1226), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT121), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1202), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1201), .A2(KEYINPUT122), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT122), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1160), .B1(new_n1157), .B2(new_n1168), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n978), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT121), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1231), .A2(new_n1203), .ZN(new_n1241));
  OAI21_X1  g1041(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1237), .B1(new_n1238), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1236), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT120), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1233), .A2(new_n1239), .A3(KEYINPUT120), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1202), .B1(new_n1238), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n711), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1244), .A2(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1248), .A2(new_n1003), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1218), .A2(new_n785), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n771), .B1(G50), .B2(new_n862), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n250), .A2(G41), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n815), .B2(new_n821), .C1(new_n572), .C2(new_n825), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1071), .B1(G58), .B2(new_n833), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G97), .A2(new_n807), .B1(new_n813), .B2(G107), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1046), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1256), .B(new_n1259), .C1(G116), .C2(new_n799), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT58), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1255), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1262), .B(new_n280), .C1(G33), .C2(G41), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n799), .A2(G125), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n802), .A2(G150), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n820), .A2(new_n1185), .B1(new_n832), .B2(G137), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(G128), .A2(new_n813), .B1(new_n807), .B2(G132), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(KEYINPUT59), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(KEYINPUT59), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n833), .A2(G159), .ZN(new_n1272));
  AOI211_X1 g1072(.A(G33), .B(G41), .C1(new_n822), .C2(G124), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n1264), .B1(KEYINPUT58), .B2(new_n1260), .C1(new_n1270), .C2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1254), .B1(new_n1275), .B2(new_n784), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1252), .B1(new_n1253), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1251), .A2(new_n1277), .ZN(G375));
  OAI221_X1 g1078(.A(new_n250), .B1(new_n801), .B2(new_n280), .C1(new_n320), .C2(new_n817), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(G137), .A2(new_n813), .B1(new_n807), .B2(new_n1185), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n366), .B2(new_n825), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1279), .B(new_n1281), .C1(G132), .C2(new_n799), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G159), .A2(new_n820), .B1(new_n822), .B2(G128), .ZN(new_n1283));
  XOR2_X1   g1083(.A(new_n1283), .B(KEYINPUT123), .Z(new_n1284));
  OAI22_X1  g1084(.A1(new_n432), .A2(new_n806), .B1(new_n812), .B2(new_n815), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(new_n1074), .A2(new_n1285), .A3(new_n250), .A4(new_n1048), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(G97), .A2(new_n820), .B1(new_n832), .B2(G107), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n466), .B2(new_n821), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(G294), .B2(new_n799), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1282), .A2(new_n1284), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1290));
  OAI221_X1 g1090(.A(new_n771), .B1(G68), .B2(new_n862), .C1(new_n1290), .C2(new_n1173), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n929), .B2(new_n785), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1166), .A2(new_n1164), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1292), .B1(new_n1295), .B2(new_n1002), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1200), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n984), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1295), .A2(new_n1200), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1296), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  XOR2_X1   g1100(.A(new_n1300), .B(KEYINPUT124), .Z(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(G381));
  NAND4_X1  g1102(.A1(new_n1251), .A2(new_n1170), .A3(new_n1193), .A4(new_n1277), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1100), .A2(new_n1122), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n1057), .A3(new_n1030), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(G384), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(G393), .A2(G396), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1306), .A2(new_n1301), .A3(new_n1307), .A4(new_n1308), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1303), .A2(new_n1309), .ZN(G407));
  OAI211_X1 g1110(.A(G407), .B(G213), .C1(G343), .C2(new_n1303), .ZN(G409));
  INV_X1    g1111(.A(KEYINPUT60), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1295), .B2(new_n1200), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1160), .A2(KEYINPUT60), .A3(new_n1167), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1313), .A2(new_n711), .A3(new_n1297), .A4(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G384), .B1(new_n1315), .B2(new_n1296), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(G213), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1318), .A2(G343), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1315), .A2(G384), .A3(new_n1296), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1317), .A2(G2897), .A3(new_n1319), .A4(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(G2897), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1320), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1322), .B1(new_n1323), .B2(new_n1316), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1321), .A2(KEYINPUT125), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT125), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(G378), .B(new_n1277), .C1(new_n1244), .C2(new_n1250), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n984), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1238), .A2(new_n1248), .A3(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1002), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1253), .A2(new_n1276), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1170), .B(new_n1193), .C1(new_n1330), .C2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1319), .B1(new_n1328), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1327), .A2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n846), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1308), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1304), .B1(new_n1030), .B2(new_n1057), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1339), .B1(new_n1306), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(G387), .A2(G390), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1342), .B(new_n1305), .C1(new_n1308), .C2(new_n1338), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1344), .A2(KEYINPUT61), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT63), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1323), .A2(new_n1316), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1335), .A2(new_n1346), .A3(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1346), .B1(new_n1335), .B2(new_n1347), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1337), .B(new_n1345), .C1(new_n1348), .C2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT62), .ZN(new_n1351));
  AND3_X1   g1151(.A1(new_n1335), .A2(new_n1351), .A3(new_n1347), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT61), .ZN(new_n1353));
  AND2_X1   g1153(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1353), .B1(new_n1335), .B2(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1351), .B1(new_n1335), .B2(new_n1347), .ZN(new_n1356));
  NOR3_X1   g1156(.A1(new_n1352), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1357));
  AND2_X1   g1157(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1350), .B1(new_n1357), .B2(new_n1358), .ZN(G405));
  INV_X1    g1159(.A(KEYINPUT126), .ZN(new_n1360));
  OR3_X1    g1160(.A1(new_n1347), .A2(new_n1360), .A3(KEYINPUT127), .ZN(new_n1361));
  OAI21_X1  g1161(.A(KEYINPUT127), .B1(new_n1347), .B2(new_n1360), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1358), .A2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1344), .A2(new_n1362), .A3(new_n1361), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1364), .A2(new_n1365), .ZN(new_n1366));
  AOI21_X1  g1166(.A(G378), .B1(new_n1251), .B2(new_n1277), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1347), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1328), .B1(KEYINPUT126), .B2(new_n1368), .ZN(new_n1369));
  OAI21_X1  g1169(.A(new_n1366), .B1(new_n1367), .B2(new_n1369), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1367), .A2(new_n1369), .ZN(new_n1371));
  NAND3_X1  g1171(.A1(new_n1364), .A2(new_n1371), .A3(new_n1365), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1370), .A2(new_n1372), .ZN(G402));
endmodule


