//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n194), .B1(new_n191), .B2(new_n193), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n189), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(new_n193), .ZN(new_n198));
  OR2_X1    g012(.A1(new_n198), .A2(new_n189), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(new_n201), .B2(G107), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  XOR2_X1   g021(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(G101), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n202), .A2(new_n205), .A3(new_n210), .A4(new_n206), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT74), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(G101), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT4), .B1(new_n214), .B2(KEYINPUT74), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n200), .B(new_n209), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n201), .A2(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n204), .A2(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n211), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT5), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n195), .A2(new_n196), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(G113), .B1(new_n191), .B2(KEYINPUT5), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n199), .B(new_n221), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g040(.A(G110), .B(G122), .Z(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n227), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n217), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(KEYINPUT6), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  INV_X1    g047(.A(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G143), .ZN(new_n235));
  INV_X1    g049(.A(G143), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G146), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n233), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n236), .A2(KEYINPUT64), .A3(G146), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT64), .B1(new_n236), .B2(G146), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n235), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n236), .A2(G146), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n243));
  OAI21_X1  g057(.A(G128), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n238), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G125), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n235), .A2(new_n237), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(new_n234), .B2(G143), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n236), .A2(KEYINPUT64), .A3(G146), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n242), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n250), .B1(new_n256), .B2(new_n249), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n247), .B1(new_n257), .B2(new_n246), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G224), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n258), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT79), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n264));
  AND4_X1   g078(.A1(new_n263), .A2(new_n226), .A3(new_n264), .A4(new_n227), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n229), .B1(new_n217), .B2(new_n225), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n263), .B1(new_n266), .B2(new_n264), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n231), .B(new_n262), .C1(new_n265), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n226), .A2(new_n264), .A3(new_n227), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT79), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(new_n263), .A3(new_n264), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n274), .A2(KEYINPUT80), .A3(new_n231), .A4(new_n262), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT7), .ZN(new_n277));
  OR4_X1    g091(.A1(KEYINPUT82), .A2(new_n258), .A3(new_n277), .A4(new_n261), .ZN(new_n278));
  AND2_X1   g092(.A1(KEYINPUT82), .A2(KEYINPUT7), .ZN(new_n279));
  OAI22_X1  g093(.A1(new_n258), .A2(new_n279), .B1(new_n277), .B2(new_n261), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n198), .A2(new_n222), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n199), .B1(new_n281), .B2(new_n224), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n227), .B(KEYINPUT81), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT8), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n221), .A2(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n199), .B1(new_n223), .B2(new_n224), .ZN(new_n286));
  OAI221_X1 g100(.A(new_n285), .B1(new_n284), .B2(new_n283), .C1(new_n221), .C2(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n278), .A2(new_n280), .A3(new_n230), .A4(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n188), .B1(new_n276), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n188), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n293), .B(new_n290), .C1(new_n270), .C2(new_n275), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n187), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT83), .ZN(new_n296));
  NOR2_X1   g110(.A1(G475), .A2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G237), .A2(G953), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n299), .A2(G143), .A3(G214), .ZN(new_n300));
  AOI21_X1  g114(.A(G143), .B1(new_n299), .B2(G214), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n300), .A2(new_n301), .A3(G131), .ZN(new_n302));
  INV_X1    g116(.A(G131), .ZN(new_n303));
  INV_X1    g117(.A(G237), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n259), .A3(G214), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n236), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n299), .A2(G143), .A3(G214), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT85), .B1(new_n302), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G125), .B(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT16), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G125), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n311), .B(G146), .C1(KEYINPUT16), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT19), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(new_n315), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n234), .ZN(new_n318));
  OAI21_X1  g132(.A(G131), .B1(new_n300), .B2(new_n301), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n306), .A2(new_n303), .A3(new_n307), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n309), .A2(new_n314), .A3(new_n318), .A4(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(new_n310), .B2(new_n234), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n246), .A2(G140), .ZN(new_n326));
  AND4_X1   g140(.A1(new_n324), .A2(new_n313), .A3(new_n326), .A4(new_n234), .ZN(new_n327));
  OAI22_X1  g141(.A1(new_n325), .A2(new_n327), .B1(new_n234), .B2(new_n310), .ZN(new_n328));
  NAND2_X1  g142(.A1(KEYINPUT18), .A2(G131), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n300), .B2(new_n301), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n306), .A2(KEYINPUT18), .A3(G131), .A4(new_n307), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT84), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n328), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n328), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n323), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G113), .B(G122), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(new_n201), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n311), .B1(KEYINPUT16), .B2(new_n313), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n234), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT17), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n319), .A2(new_n343), .A3(new_n321), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n308), .A2(KEYINPUT17), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n342), .A2(new_n344), .A3(new_n314), .A4(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n338), .B(new_n346), .C1(new_n334), .C2(new_n335), .ZN(new_n347));
  AOI211_X1 g161(.A(KEYINPUT20), .B(new_n298), .C1(new_n340), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n328), .A2(new_n332), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT84), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n328), .A2(new_n332), .A3(new_n333), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n338), .B1(new_n353), .B2(new_n323), .ZN(new_n354));
  INV_X1    g168(.A(new_n347), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT86), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT86), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n340), .A2(new_n357), .A3(new_n347), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n298), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n349), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n338), .B1(new_n353), .B2(new_n346), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n362), .A2(new_n355), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n289), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G475), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT9), .B(G234), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n367), .A2(new_n368), .A3(G953), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n236), .A2(G128), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n232), .A2(G143), .ZN(new_n372));
  INV_X1    g186(.A(G134), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G122), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G116), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n192), .A2(G122), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n378), .A3(new_n204), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT13), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT87), .B1(new_n371), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n384), .A2(new_n236), .A3(KEYINPUT13), .A4(G128), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n371), .A2(new_n382), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n383), .A2(new_n372), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  AOI221_X4 g201(.A(new_n375), .B1(new_n380), .B2(new_n381), .C1(new_n387), .C2(G134), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n371), .A2(new_n372), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G134), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n374), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n192), .A2(KEYINPUT14), .A3(G122), .ZN(new_n392));
  OAI211_X1 g206(.A(G107), .B(new_n392), .C1(new_n379), .C2(KEYINPUT14), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n381), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n370), .B1(new_n388), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n387), .A2(G134), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n380), .A2(new_n381), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n374), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n394), .A3(new_n369), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(KEYINPUT88), .B(new_n370), .C1(new_n388), .C2(new_n395), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n289), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G478), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(KEYINPUT15), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n406), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n402), .A2(new_n289), .A3(new_n403), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT89), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n407), .A2(KEYINPUT89), .A3(new_n409), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n366), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G469), .ZN(new_n416));
  XNOR2_X1  g230(.A(G110), .B(G140), .ZN(new_n417));
  INV_X1    g231(.A(G227), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G953), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n417), .B(new_n419), .Z(new_n420));
  OAI211_X1 g234(.A(new_n257), .B(new_n209), .C1(new_n215), .C2(new_n216), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT76), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n211), .A2(new_n220), .A3(KEYINPUT10), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n422), .B1(new_n245), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n233), .A2(new_n235), .A3(new_n237), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n232), .B1(new_n235), .B2(KEYINPUT1), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n425), .B1(new_n254), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n221), .A2(new_n427), .A3(KEYINPUT76), .A4(KEYINPUT10), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n244), .A2(new_n248), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n425), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n221), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT10), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n421), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(KEYINPUT65), .A2(G137), .ZN(new_n436));
  NOR2_X1   g250(.A1(KEYINPUT65), .A2(G137), .ZN(new_n437));
  OAI211_X1 g251(.A(KEYINPUT11), .B(G134), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G137), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT66), .B1(new_n439), .B2(G134), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT66), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n373), .A3(G137), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT11), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n373), .B2(G137), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G131), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n438), .A2(new_n443), .A3(new_n303), .A4(new_n445), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n435), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT78), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n435), .A2(new_n452), .A3(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n449), .B(KEYINPUT77), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n435), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n420), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n420), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT12), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n432), .B1(new_n427), .B2(new_n221), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n460), .B1(new_n461), .B2(new_n449), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n461), .A2(new_n460), .A3(new_n449), .ZN(new_n463));
  NOR4_X1   g277(.A1(new_n456), .A2(new_n459), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n416), .B(new_n289), .C1(new_n458), .C2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n416), .A2(new_n289), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n435), .A2(new_n452), .A3(new_n449), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n452), .B1(new_n435), .B2(new_n449), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n457), .B(new_n420), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n463), .A2(new_n462), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n459), .B1(new_n471), .B2(new_n456), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n472), .A3(G469), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(new_n467), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n415), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n259), .A2(G952), .ZN(new_n477));
  INV_X1    g291(.A(G234), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(new_n304), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI211_X1 g294(.A(new_n289), .B(new_n259), .C1(G234), .C2(G237), .ZN(new_n481));
  XOR2_X1   g295(.A(KEYINPUT21), .B(G898), .Z(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(new_n187), .C1(new_n292), .C2(new_n294), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n296), .A2(new_n476), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT32), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT31), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n449), .A2(new_n257), .ZN(new_n491));
  INV_X1    g305(.A(new_n200), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n436), .A2(new_n437), .A3(G134), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n373), .A2(G137), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n427), .A2(new_n448), .A3(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n491), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(KEYINPUT67), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(KEYINPUT67), .ZN(new_n501));
  INV_X1    g315(.A(new_n255), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n241), .A2(new_n249), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n250), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(new_n447), .B2(new_n448), .ZN(new_n506));
  INV_X1    g320(.A(new_n496), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n500), .B(new_n501), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n491), .A2(KEYINPUT67), .A3(new_n498), .A4(new_n496), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n497), .B1(new_n510), .B2(new_n200), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n299), .A2(G210), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(G101), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n490), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n492), .B1(new_n508), .B2(new_n509), .ZN(new_n517));
  INV_X1    g331(.A(new_n515), .ZN(new_n518));
  NOR4_X1   g332(.A1(new_n517), .A2(KEYINPUT31), .A3(new_n497), .A4(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n515), .B(KEYINPUT69), .Z(new_n520));
  AOI21_X1  g334(.A(new_n492), .B1(new_n491), .B2(new_n496), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT28), .B1(new_n497), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n491), .A2(new_n492), .A3(new_n496), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n520), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n516), .A2(new_n519), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(G472), .A2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n489), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n501), .ZN(new_n531));
  AOI211_X1 g345(.A(new_n499), .B(new_n531), .C1(new_n491), .C2(new_n496), .ZN(new_n532));
  INV_X1    g346(.A(new_n509), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n200), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n523), .A3(new_n515), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT31), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n511), .A2(new_n490), .A3(new_n515), .ZN(new_n537));
  INV_X1    g351(.A(new_n526), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(KEYINPUT32), .A3(new_n528), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n511), .A2(new_n515), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n522), .A2(new_n525), .A3(new_n520), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT29), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n522), .A2(KEYINPUT29), .A3(new_n525), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n289), .B1(new_n544), .B2(new_n518), .ZN(new_n545));
  OAI21_X1  g359(.A(G472), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n530), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n368), .B1(G234), .B2(new_n289), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n325), .A2(new_n327), .ZN(new_n549));
  XOR2_X1   g363(.A(G119), .B(G128), .Z(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT70), .ZN(new_n551));
  XOR2_X1   g365(.A(KEYINPUT24), .B(G110), .Z(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT23), .B1(new_n232), .B2(G119), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT71), .B1(new_n232), .B2(G119), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(G110), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n314), .B(new_n549), .C1(new_n553), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n342), .A2(new_n314), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(G110), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n551), .A2(new_n552), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT22), .B(G137), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n563), .B(new_n564), .Z(new_n565));
  AND3_X1   g379(.A1(new_n558), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n565), .B1(new_n558), .B2(new_n562), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT25), .B1(new_n568), .B2(new_n289), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT25), .ZN(new_n570));
  NOR4_X1   g384(.A1(new_n566), .A2(new_n567), .A3(new_n570), .A4(G902), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n548), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n548), .A2(G902), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT73), .ZN(new_n574));
  INV_X1    g388(.A(new_n568), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n547), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n488), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT90), .B(G101), .Z(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(G3));
  AOI21_X1  g395(.A(new_n526), .B1(new_n535), .B2(KEYINPUT31), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n582), .B2(new_n537), .ZN(new_n583));
  INV_X1    g397(.A(G472), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT91), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n586), .B(G472), .C1(new_n527), .C2(G902), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n539), .A2(new_n528), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n475), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n457), .B1(new_n468), .B2(new_n469), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n459), .ZN(new_n592));
  INV_X1    g406(.A(new_n464), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n466), .B1(new_n594), .B2(new_n416), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n590), .B1(new_n595), .B2(new_n473), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n589), .A2(new_n577), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n485), .B(new_n187), .C1(new_n292), .C2(new_n294), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n402), .A2(new_n599), .A3(new_n403), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n396), .A2(KEYINPUT33), .A3(new_n401), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n600), .A2(G478), .A3(new_n289), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n404), .A2(new_n405), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n366), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n597), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT34), .B(G104), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  INV_X1    g423(.A(new_n187), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n276), .A2(new_n291), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n293), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n276), .A2(new_n188), .A3(new_n291), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT92), .B1(new_n359), .B2(new_n360), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n340), .A2(new_n357), .A3(new_n347), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n357), .B1(new_n340), .B2(new_n347), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n297), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT92), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n619), .A3(KEYINPUT20), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n360), .B(new_n297), .C1(new_n616), .C2(new_n617), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT93), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n359), .A2(new_n623), .A3(new_n360), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n615), .A2(new_n620), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n625), .A2(new_n365), .A3(new_n414), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n614), .A2(new_n626), .A3(KEYINPUT94), .A4(new_n485), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n625), .A2(new_n365), .A3(new_n414), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n628), .B1(new_n598), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n597), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND3_X1  g448(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n558), .A2(new_n562), .ZN(new_n636));
  INV_X1    g450(.A(new_n565), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(KEYINPUT36), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n636), .B(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n574), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n572), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n488), .A2(new_n635), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT37), .B(G110), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  OAI211_X1 g460(.A(new_n187), .B(new_n642), .C1(new_n292), .C2(new_n294), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n481), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n479), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n629), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n648), .A2(new_n653), .A3(new_n547), .A4(new_n596), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  XNOR2_X1  g469(.A(new_n651), .B(KEYINPUT39), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n596), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT40), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n612), .A2(new_n613), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT38), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n292), .A2(new_n294), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT38), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n348), .B1(new_n618), .B2(KEYINPUT20), .ZN(new_n664));
  INV_X1    g478(.A(new_n365), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n414), .B(new_n187), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n661), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT95), .ZN(new_n669));
  INV_X1    g483(.A(new_n535), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n497), .A2(new_n521), .ZN(new_n671));
  INV_X1    g485(.A(new_n520), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n673), .B2(G902), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n530), .A2(new_n674), .A3(new_n540), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n643), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n668), .A2(new_n669), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n669), .B1(new_n668), .B2(new_n676), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n658), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n236), .ZN(G45));
  NAND3_X1  g495(.A1(new_n366), .A2(new_n604), .A3(new_n651), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n648), .A2(new_n547), .A3(new_n596), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  AOI211_X1 g499(.A(new_n489), .B(new_n529), .C1(new_n582), .C2(new_n537), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT32), .B1(new_n539), .B2(new_n528), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n576), .B1(new_n688), .B2(new_n546), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n464), .B1(new_n459), .B2(new_n591), .ZN(new_n690));
  OAI21_X1  g504(.A(G469), .B1(new_n690), .B2(G902), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n691), .A2(new_n475), .A3(new_n465), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n606), .A2(new_n689), .A3(KEYINPUT96), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT96), .ZN(new_n694));
  INV_X1    g508(.A(new_n605), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n659), .A2(new_n485), .A3(new_n187), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n547), .A2(new_n577), .A3(new_n692), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  INV_X1    g515(.A(new_n697), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n631), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  INV_X1    g518(.A(new_n692), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n705), .A2(new_n295), .A3(new_n484), .A4(new_n643), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n547), .A2(new_n415), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  INV_X1    g523(.A(KEYINPUT97), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n519), .B1(new_n582), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT97), .B1(new_n516), .B2(new_n526), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n529), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n584), .B1(new_n539), .B2(new_n289), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n576), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n666), .B1(new_n612), .B2(new_n613), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n715), .A2(new_n485), .A3(new_n716), .A4(new_n692), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  NOR3_X1   g532(.A1(new_n713), .A2(new_n682), .A3(new_n714), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n614), .A3(new_n642), .A4(new_n692), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  NAND2_X1  g535(.A1(new_n470), .A2(KEYINPUT98), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT98), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n454), .A2(new_n723), .A3(new_n420), .A4(new_n457), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(new_n724), .A3(G469), .A4(new_n472), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n590), .B1(new_n595), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n547), .A3(new_n577), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n683), .A2(new_n662), .A3(new_n187), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT42), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n727), .B2(new_n728), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT99), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT99), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n730), .A2(new_n735), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT100), .B(G131), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G33));
  NAND2_X1  g553(.A1(new_n662), .A2(new_n187), .ZN(new_n740));
  NOR4_X1   g554(.A1(new_n727), .A2(new_n740), .A3(new_n629), .A4(new_n652), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n373), .ZN(G36));
  NAND3_X1  g556(.A1(new_n361), .A2(new_n365), .A3(new_n604), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(new_n635), .A3(KEYINPUT44), .A4(new_n642), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(KEYINPUT101), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n740), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n722), .A2(new_n724), .A3(KEYINPUT45), .A4(new_n472), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n470), .A2(new_n472), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(G469), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n467), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n465), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT46), .B1(new_n753), .B2(new_n467), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n475), .B(new_n656), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(KEYINPUT101), .B2(new_n746), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n745), .A2(new_n635), .A3(new_n642), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT102), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(KEYINPUT102), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n748), .B(new_n758), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  INV_X1    g579(.A(KEYINPUT103), .ZN(new_n766));
  OR4_X1    g580(.A1(new_n766), .A2(new_n728), .A3(new_n577), .A4(new_n547), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n659), .A2(new_n610), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n576), .A3(new_n683), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n766), .B1(new_n769), .B2(new_n547), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n475), .B1(new_n755), .B2(new_n756), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n740), .A2(new_n705), .A3(KEYINPUT114), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT114), .B1(new_n740), .B2(new_n705), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n713), .A2(new_n714), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n745), .A2(new_n480), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n642), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n675), .A2(new_n479), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n366), .A2(new_n604), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n780), .A2(new_n577), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n715), .A2(new_n480), .A3(new_n745), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n661), .A2(new_n663), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n610), .A3(new_n788), .A4(new_n692), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(KEYINPUT113), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n790), .B1(new_n789), .B2(KEYINPUT113), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n783), .B(new_n786), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n772), .B(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n691), .A2(new_n465), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT104), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n590), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n787), .A2(new_n768), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n777), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n780), .A2(new_n689), .A3(new_n782), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT48), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n780), .A2(new_n577), .A3(new_n695), .A4(new_n784), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n787), .A2(new_n614), .A3(new_n692), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n477), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n806), .A2(KEYINPUT116), .A3(new_n477), .A4(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n803), .A2(new_n805), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n794), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n799), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n795), .A2(KEYINPUT115), .A3(new_n798), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n800), .A3(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n814), .A2(new_n818), .A3(KEYINPUT51), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT117), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT108), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n651), .B(KEYINPUT107), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n642), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n572), .A2(KEYINPUT108), .A3(new_n641), .A4(new_n822), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n716), .A2(new_n826), .A3(new_n675), .A4(new_n726), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT109), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n654), .A2(new_n684), .A3(new_n720), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT52), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT109), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n827), .B(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n654), .A2(new_n684), .A3(new_n720), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n644), .A2(new_n579), .ZN(new_n837));
  INV_X1    g651(.A(new_n717), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n698), .B2(new_n693), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n631), .A2(new_n702), .B1(new_n706), .B2(new_n707), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n361), .A2(new_n365), .A3(new_n410), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n605), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n589), .A2(new_n577), .A3(new_n596), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n296), .A2(new_n485), .A3(new_n487), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n837), .A2(new_n839), .A3(new_n840), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n410), .A2(new_n652), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n625), .A2(new_n365), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT106), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n625), .A2(KEYINPUT106), .A3(new_n365), .A4(new_n847), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n596), .A3(new_n547), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n781), .A2(new_n726), .A3(new_n683), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n643), .B(new_n740), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n836), .A2(new_n846), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n741), .B1(new_n734), .B2(new_n736), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT53), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n699), .A2(new_n703), .A3(new_n708), .A4(new_n717), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n843), .A2(new_n844), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n644), .A2(new_n579), .A3(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n859), .A2(new_n830), .A3(new_n861), .A4(new_n835), .ZN(new_n862));
  INV_X1    g676(.A(new_n741), .ZN(new_n863));
  INV_X1    g677(.A(new_n736), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n735), .B1(new_n730), .B2(new_n732), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n862), .A2(new_n866), .A3(new_n867), .A4(new_n854), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n857), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n783), .A2(new_n786), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n870), .B(new_n801), .C1(new_n793), .C2(new_n792), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n871), .A2(new_n777), .B1(new_n810), .B2(new_n811), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n814), .A2(new_n818), .A3(KEYINPUT51), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n805), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT111), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n858), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT111), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n733), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT112), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT110), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n854), .A2(new_n741), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n861), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n836), .ZN(new_n884));
  INV_X1    g698(.A(new_n488), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n589), .A3(new_n642), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n689), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n845), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n852), .A2(new_n853), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(new_n642), .A3(new_n768), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n863), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n867), .B1(new_n892), .B2(new_n881), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT112), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n877), .A2(new_n878), .A3(new_n894), .A4(new_n733), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n880), .A2(new_n884), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n830), .A2(new_n835), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n888), .A2(new_n858), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n856), .A3(new_n898), .A4(new_n890), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n867), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n896), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n820), .A2(new_n869), .A3(new_n875), .A4(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(G952), .B2(G953), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT49), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n590), .B1(new_n797), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n576), .A2(new_n610), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n906), .B(new_n907), .C1(new_n905), .C2(new_n797), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n788), .A2(new_n688), .A3(new_n674), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n743), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT105), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n904), .A2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n266), .A2(new_n264), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n272), .A2(new_n273), .B1(new_n913), .B2(new_n230), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n262), .ZN(new_n915));
  XOR2_X1   g729(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(KEYINPUT119), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(G210), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n921), .B(new_n289), .C1(new_n896), .C2(new_n900), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n922), .B2(KEYINPUT56), .ZN(new_n923));
  INV_X1    g737(.A(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n896), .A2(new_n900), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(G902), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n919), .B(new_n924), .C1(new_n926), .C2(new_n921), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n259), .A2(G952), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n923), .A2(new_n927), .A3(new_n929), .ZN(G51));
  XNOR2_X1  g744(.A(new_n466), .B(KEYINPUT57), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n896), .A2(new_n901), .A3(new_n900), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n901), .B1(new_n896), .B2(new_n900), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n690), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n926), .A2(new_n753), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n928), .B1(new_n936), .B2(new_n937), .ZN(G54));
  AOI21_X1  g752(.A(new_n289), .B1(new_n896), .B2(new_n900), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(KEYINPUT58), .A3(G475), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n356), .A2(new_n358), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(KEYINPUT58), .A3(G475), .A4(new_n941), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n943), .A2(new_n929), .A3(new_n944), .ZN(G60));
  XNOR2_X1  g759(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n405), .A2(new_n289), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n946), .B(new_n947), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n869), .B2(new_n902), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n600), .A2(new_n601), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n929), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n951), .B(new_n948), .C1(new_n932), .C2(new_n933), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n952), .A2(new_n954), .ZN(G63));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT60), .Z(new_n958));
  NAND3_X1  g772(.A1(new_n925), .A2(new_n639), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n929), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n568), .B1(new_n925), .B2(new_n958), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n925), .A2(new_n958), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n575), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n964), .A2(KEYINPUT61), .A3(new_n929), .A4(new_n959), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(G66));
  AOI21_X1  g780(.A(new_n259), .B1(new_n482), .B2(G224), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n846), .B(KEYINPUT121), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n259), .ZN(new_n969));
  INV_X1    g783(.A(G898), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n914), .B1(new_n970), .B2(G953), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT122), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n969), .B(new_n972), .ZN(G69));
  INV_X1    g787(.A(new_n757), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n689), .A3(new_n716), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n775), .A2(new_n764), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n866), .A2(KEYINPUT124), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n737), .A2(new_n978), .A3(new_n863), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n976), .A2(new_n977), .A3(new_n979), .A4(new_n833), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n259), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n316), .A2(new_n317), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n510), .B(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(G953), .B1(new_n418), .B2(new_n649), .ZN(new_n985));
  XOR2_X1   g799(.A(KEYINPUT125), .B(G900), .Z(new_n986));
  OAI211_X1 g800(.A(new_n981), .B(new_n984), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n775), .A2(new_n764), .ZN(new_n988));
  NAND2_X1  g802(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n989));
  INV_X1    g803(.A(new_n679), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(new_n677), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n833), .B(new_n989), .C1(new_n991), .C2(new_n658), .ZN(new_n992));
  XNOR2_X1  g806(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n680), .B2(new_n829), .ZN(new_n994));
  INV_X1    g808(.A(new_n842), .ZN(new_n995));
  OR4_X1    g809(.A1(new_n578), .A2(new_n657), .A3(new_n740), .A4(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n988), .A2(new_n992), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n259), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n985), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n983), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n987), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  OAI21_X1  g819(.A(new_n1005), .B1(new_n980), .B2(new_n968), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n511), .A3(new_n518), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1007), .A2(KEYINPUT127), .A3(new_n929), .ZN(new_n1008));
  AOI21_X1  g822(.A(KEYINPUT127), .B1(new_n1007), .B2(new_n929), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1005), .B1(new_n968), .B2(new_n997), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n1010), .B(new_n515), .C1(new_n497), .C2(new_n517), .ZN(new_n1011));
  OAI221_X1 g825(.A(new_n1005), .B1(new_n670), .B2(new_n541), .C1(new_n857), .C2(new_n868), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1008), .A2(new_n1009), .A3(new_n1013), .ZN(G57));
endmodule


