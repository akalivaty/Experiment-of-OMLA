//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1219,
    new_n1220, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OR2_X1    g0008(.A1(new_n208), .A2(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n212), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n208), .A2(KEYINPUT0), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n209), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  AOI22_X1  g0022(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  INV_X1    g0030(.A(G68), .ZN(new_n231));
  INV_X1    g0031(.A(G238), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n205), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n222), .A2(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n215), .A2(new_n253), .A3(KEYINPUT67), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G20), .B2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G50), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT73), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n215), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n261), .A2(G77), .B1(G20), .B2(new_n231), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n205), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n214), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(KEYINPUT11), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(new_n215), .A3(G1), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT74), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n270), .A2(G68), .B1(new_n271), .B2(KEYINPUT12), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT12), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(KEYINPUT74), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n271), .B(KEYINPUT12), .C1(new_n270), .C2(G68), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n266), .A2(new_n269), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n215), .A2(G1), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(new_n231), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n267), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT11), .B1(new_n263), .B2(new_n266), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT13), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n253), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n230), .A2(G1698), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n289), .B(new_n290), .C1(G226), .C2(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G97), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT72), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n211), .A2(new_n213), .A3(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n291), .A2(KEYINPUT72), .A3(new_n292), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G274), .ZN(new_n300));
  AND2_X1   g0100(.A1(G1), .A2(G13), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n294), .ZN(new_n302));
  INV_X1    g0102(.A(G1), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(G41), .B2(G45), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n294), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n304), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n306), .B1(new_n232), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n285), .B1(new_n299), .B2(new_n310), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n297), .A2(new_n293), .A3(new_n295), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n312), .A2(KEYINPUT13), .A3(new_n309), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n284), .B(G169), .C1(new_n311), .C2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT13), .B1(new_n312), .B2(new_n309), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n299), .A2(new_n285), .A3(new_n310), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(G179), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n316), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n284), .B1(new_n319), .B2(G169), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n283), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(G200), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n322), .B(new_n282), .C1(new_n323), .C2(new_n319), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G200), .ZN(new_n326));
  INV_X1    g0126(.A(new_n306), .ZN(new_n327));
  INV_X1    g0127(.A(new_n308), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n327), .B1(G226), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n295), .ZN(new_n330));
  INV_X1    g0130(.A(G1698), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G222), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G223), .A2(G1698), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n289), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n330), .B(new_n334), .C1(G77), .C2(new_n289), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n326), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n329), .A2(new_n335), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(G190), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT70), .B(KEYINPUT10), .ZN(new_n339));
  INV_X1    g0139(.A(new_n277), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n276), .A2(G50), .A3(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n254), .A2(new_n256), .ZN(new_n342));
  INV_X1    g0142(.A(G150), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT8), .B(G58), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n345), .A2(new_n260), .B1(new_n215), .B2(new_n201), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n266), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n341), .B(new_n347), .C1(G50), .C2(new_n270), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n348), .A2(KEYINPUT9), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(KEYINPUT9), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n338), .B(new_n339), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT71), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n338), .B1(new_n349), .B2(new_n350), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n351), .A2(new_n352), .B1(new_n353), .B2(KEYINPUT10), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n352), .B2(new_n351), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n337), .A2(G169), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT68), .B(G179), .Z(new_n357));
  NAND2_X1  g0157(.A1(new_n337), .A2(new_n357), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n356), .A2(new_n348), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n327), .B1(G244), .B2(new_n328), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G238), .A2(G1698), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n289), .B(new_n362), .C1(new_n230), .C2(G1698), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n330), .C1(G107), .C2(new_n289), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n357), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(G169), .B2(new_n365), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n213), .A2(new_n211), .B1(new_n264), .B2(G33), .ZN(new_n368));
  XOR2_X1   g0168(.A(new_n345), .B(KEYINPUT69), .Z(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n257), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT15), .B(G87), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n372), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n368), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n276), .A2(G77), .A3(new_n340), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G77), .B2(new_n270), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n367), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n365), .A2(G190), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n377), .B(new_n380), .C1(new_n326), .C2(new_n365), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n325), .A2(new_n355), .A3(new_n360), .A4(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n287), .A2(new_n215), .A3(new_n288), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n215), .A4(new_n288), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n231), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(G58), .B(G68), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G20), .ZN(new_n390));
  INV_X1    g0190(.A(G159), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n342), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n368), .B1(new_n393), .B2(KEYINPUT16), .ZN(new_n394));
  AND2_X1   g0194(.A1(KEYINPUT3), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT3), .A2(G33), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT7), .B1(new_n397), .B2(new_n215), .ZN(new_n398));
  INV_X1    g0198(.A(new_n387), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n257), .A2(G159), .B1(new_n389), .B2(G20), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n388), .B2(new_n392), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT75), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n394), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n345), .A2(new_n277), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT76), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n409), .B(new_n410), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(new_n276), .B1(new_n269), .B2(new_n345), .ZN(new_n412));
  OR2_X1    g0212(.A1(G223), .A2(G1698), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n413), .B1(G226), .B2(new_n331), .C1(new_n395), .C2(new_n396), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n295), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n306), .B1(new_n230), .B2(new_n308), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n323), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G200), .B2(new_n418), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n408), .A2(new_n412), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT17), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n408), .A2(new_n423), .A3(new_n412), .A4(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT77), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n408), .A2(new_n412), .ZN(new_n429));
  INV_X1    g0229(.A(G169), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n414), .A2(new_n415), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n330), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n328), .A2(G232), .B1(new_n302), .B2(new_n305), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n416), .A2(new_n417), .A3(new_n357), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n428), .B1(new_n429), .B2(new_n437), .ZN(new_n438));
  AOI211_X1 g0238(.A(KEYINPUT18), .B(new_n436), .C1(new_n408), .C2(new_n412), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n422), .A2(KEYINPUT77), .A3(new_n424), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n427), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n383), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT87), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT5), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G41), .ZN(new_n448));
  INV_X1    g0248(.A(G41), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT5), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(G264), .A3(new_n307), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n302), .A2(new_n448), .A3(new_n450), .A4(new_n446), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(G250), .B(new_n331), .C1(new_n395), .C2(new_n396), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT85), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT85), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n289), .A2(new_n458), .A3(G250), .A4(new_n331), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT86), .B(G294), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G33), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n289), .A2(G257), .A3(G1698), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n457), .A2(new_n459), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n453), .B(new_n455), .C1(new_n463), .C2(new_n330), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n444), .B1(new_n464), .B2(new_n430), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n453), .B1(new_n463), .B2(new_n330), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n454), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(KEYINPUT87), .A3(G169), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n464), .A2(G179), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n303), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n368), .A2(new_n270), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G107), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n269), .A2(new_n473), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT25), .ZN(new_n476));
  OR2_X1    g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n289), .A2(new_n215), .A3(G87), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT22), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT22), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n289), .A2(new_n480), .A3(new_n215), .A4(G87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT23), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n215), .B2(G107), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n473), .A2(KEYINPUT23), .A3(G20), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n487), .A2(G20), .B1(new_n488), .B2(KEYINPUT84), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT84), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(KEYINPUT24), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n368), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n482), .B(new_n490), .C1(new_n492), .C2(KEYINPUT24), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n477), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n470), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n463), .A2(new_n330), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n499), .A2(new_n323), .A3(new_n452), .A4(new_n454), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(KEYINPUT88), .C1(new_n464), .C2(G200), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT88), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n467), .A2(new_n502), .A3(new_n326), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n496), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n224), .A2(G1698), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n289), .B(new_n506), .C1(G238), .C2(G1698), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n295), .B1(new_n507), .B2(new_n487), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n303), .A2(G45), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G250), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT78), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT78), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n307), .A2(new_n513), .A3(G250), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n302), .A2(new_n446), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT79), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT79), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n512), .A2(new_n515), .A3(new_n518), .A4(new_n514), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n508), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(G169), .ZN(new_n521));
  INV_X1    g0321(.A(new_n357), .ZN(new_n522));
  AOI211_X1 g0322(.A(new_n522), .B(new_n508), .C1(new_n517), .C2(new_n519), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT80), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G97), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n225), .A2(new_n525), .A3(new_n473), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n292), .A2(new_n215), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT19), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n215), .B(G68), .C1(new_n395), .C2(new_n396), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n260), .B2(new_n525), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n368), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT81), .A4(new_n531), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n534), .A2(new_n535), .B1(new_n269), .B2(new_n371), .ZN(new_n536));
  INV_X1    g0336(.A(new_n472), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n372), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT82), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n536), .A2(KEYINPUT82), .A3(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n523), .A2(KEYINPUT80), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n524), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n537), .A2(G87), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n536), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n520), .A2(G190), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n548), .C1(new_n326), .C2(new_n520), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(G20), .B1(new_n253), .B2(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G283), .ZN(new_n553));
  INV_X1    g0353(.A(G116), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n552), .A2(new_n553), .B1(G20), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT20), .B1(new_n266), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n266), .A2(KEYINPUT20), .A3(new_n555), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n557), .A2(new_n558), .B1(new_n554), .B2(new_n269), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n211), .A2(new_n213), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n331), .A2(G257), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G264), .A2(G1698), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n562), .C1(new_n395), .C2(new_n396), .ZN(new_n563));
  INV_X1    g0363(.A(G303), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n287), .A2(new_n564), .A3(new_n288), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n560), .A2(new_n563), .A3(new_n294), .A4(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n451), .A2(G270), .A3(new_n307), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n454), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n368), .A2(G116), .A3(new_n270), .A4(new_n471), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n566), .A2(G190), .A3(new_n454), .A4(new_n567), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n559), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n572), .B(KEYINPUT83), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n289), .A2(G250), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n331), .B1(new_n574), .B2(KEYINPUT4), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT4), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(G1698), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n577), .B(G244), .C1(new_n396), .C2(new_n395), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n224), .B1(new_n287), .B2(new_n288), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n553), .C1(new_n579), .C2(KEYINPUT4), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n330), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n451), .A2(G257), .A3(new_n307), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n454), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n326), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT6), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n587), .A2(new_n525), .A3(G107), .ZN(new_n588));
  XNOR2_X1  g0388(.A(G97), .B(G107), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n590), .A2(new_n215), .B1(new_n202), .B2(new_n342), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n473), .B1(new_n386), .B2(new_n387), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n266), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n270), .A2(G97), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n537), .B2(G97), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n581), .A2(G190), .A3(new_n584), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n586), .A2(new_n593), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n581), .A2(new_n584), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n598), .A2(new_n430), .B1(new_n593), .B2(new_n595), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n581), .A2(new_n357), .A3(new_n584), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n568), .A2(G169), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n269), .A2(new_n554), .ZN(new_n604));
  INV_X1    g0404(.A(new_n558), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n570), .B(new_n604), .C1(new_n605), .C2(new_n556), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(G179), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n568), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n603), .A2(new_n606), .A3(KEYINPUT21), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n573), .A2(new_n602), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n551), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n443), .A2(new_n505), .A3(new_n616), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n324), .A2(new_n378), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n321), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n422), .A2(KEYINPUT77), .A3(new_n424), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT77), .B1(new_n422), .B2(new_n424), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n412), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n403), .B1(new_n402), .B2(new_n404), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n400), .A2(KEYINPUT16), .A3(new_n401), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n266), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n624), .B1(new_n628), .B2(new_n405), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT18), .B1(new_n629), .B2(new_n436), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n436), .B1(new_n408), .B2(new_n412), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n428), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(KEYINPUT91), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT91), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n438), .B2(new_n439), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n623), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n359), .B1(new_n637), .B2(new_n355), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n599), .A2(new_n600), .ZN(new_n639));
  XNOR2_X1  g0439(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n545), .A2(new_n549), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n520), .A2(new_n357), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n517), .A2(new_n519), .ZN(new_n644));
  INV_X1    g0444(.A(new_n508), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n430), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n534), .A2(new_n535), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n371), .A2(new_n269), .ZN(new_n649));
  AND4_X1   g0449(.A1(KEYINPUT82), .A2(new_n648), .A3(new_n649), .A4(new_n538), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT82), .B1(new_n536), .B2(new_n538), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n643), .B(new_n647), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n639), .A3(new_n549), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n642), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n657), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n614), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n498), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n652), .A2(new_n549), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n593), .A2(new_n595), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n585), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n665), .A2(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n662), .A2(new_n663), .A3(new_n504), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n656), .A2(new_n660), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n638), .B1(new_n443), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT92), .Z(G369));
  NAND3_X1  g0471(.A1(new_n303), .A2(new_n215), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n606), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT93), .ZN(new_n679));
  INV_X1    g0479(.A(new_n573), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n661), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n661), .A2(new_n679), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT94), .ZN(new_n684));
  INV_X1    g0484(.A(new_n505), .ZN(new_n685));
  INV_X1    g0485(.A(new_n677), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n496), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n498), .B2(new_n686), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n684), .A2(G330), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n498), .A2(new_n677), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n661), .A2(new_n677), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n685), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n206), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G1), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n526), .A2(G116), .ZN(new_n698));
  OAI22_X1  g0498(.A1(new_n697), .A2(new_n698), .B1(new_n217), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n700));
  XNOR2_X1  g0500(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n686), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n568), .A2(new_n357), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n646), .A2(new_n467), .A3(new_n598), .A4(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n397), .A2(new_n226), .ZN(new_n708));
  OAI21_X1  g0508(.A(G1698), .B1(new_n708), .B2(new_n576), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n576), .B1(new_n397), .B2(new_n224), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n578), .A2(new_n553), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n583), .B1(new_n712), .B2(new_n330), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n713), .A2(new_n520), .A3(new_n466), .A4(new_n611), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT96), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT30), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n611), .A2(new_n466), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(KEYINPUT96), .A3(new_n520), .A4(new_n713), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n707), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(KEYINPUT97), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n719), .B2(KEYINPUT97), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n704), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n551), .A2(new_n685), .A3(new_n615), .A4(new_n686), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n714), .A2(new_n715), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n718), .A3(new_n721), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n722), .A3(new_n706), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n677), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n703), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT98), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT98), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n730), .A2(new_n733), .A3(new_n703), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n702), .B1(new_n726), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n545), .A2(new_n549), .A3(new_n639), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n652), .A2(new_n549), .A3(new_n639), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n738), .A2(new_n640), .B1(new_n739), .B2(KEYINPUT26), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n666), .A2(new_n504), .A3(new_n652), .A4(new_n549), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n614), .B1(new_n497), .B2(new_n470), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n659), .B(new_n658), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n686), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n668), .A2(new_n746), .A3(new_n686), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n737), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n701), .B1(new_n749), .B2(G1), .ZN(G364));
  NAND2_X1  g0550(.A1(new_n684), .A2(G330), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n268), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n697), .B1(G45), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n684), .A2(G330), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n684), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n214), .B1(G20), .B2(new_n430), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n759), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n694), .A2(new_n289), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n445), .B2(new_n218), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(new_n248), .B2(new_n445), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n694), .A2(new_n397), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n769), .A2(G355), .B1(new_n554), .B2(new_n694), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n323), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n215), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n215), .A2(G179), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n774), .A2(new_n460), .B1(new_n777), .B2(G303), .ZN(new_n778));
  INV_X1    g0578(.A(G283), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n775), .A2(new_n323), .A3(G200), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n215), .A2(new_n323), .A3(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n522), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n215), .A2(G190), .A3(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n610), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n784), .A2(G322), .B1(new_n787), .B2(G329), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n522), .A2(new_n785), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n788), .B(new_n397), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n357), .A2(new_n326), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n215), .A2(new_n323), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n781), .B(new_n791), .C1(G326), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n215), .A2(G190), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n792), .A2(KEYINPUT100), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT100), .B1(new_n792), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n783), .A2(new_n229), .B1(new_n790), .B2(new_n202), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT99), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n777), .A2(G87), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(new_n806), .B2(new_n289), .ZN(new_n807));
  AOI211_X1 g0607(.A(KEYINPUT99), .B(new_n397), .C1(new_n777), .C2(G87), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n773), .A2(new_n525), .B1(new_n780), .B2(new_n473), .ZN(new_n809));
  NOR4_X1   g0609(.A1(new_n804), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n786), .A2(KEYINPUT32), .A3(new_n391), .ZN(new_n811));
  OAI21_X1  g0611(.A(KEYINPUT32), .B1(new_n786), .B2(new_n391), .ZN(new_n812));
  INV_X1    g0612(.A(G50), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n794), .B2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n811), .B(new_n814), .C1(new_n801), .C2(G68), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n796), .A2(new_n803), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n762), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n753), .B1(new_n764), .B2(new_n771), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n755), .A2(new_n756), .B1(new_n761), .B2(new_n818), .ZN(G396));
  OAI21_X1  g0619(.A(new_n381), .B1(new_n377), .B2(new_n686), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n379), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n378), .A2(new_n686), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n669), .B2(new_n677), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n382), .A2(new_n686), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n668), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n753), .B1(new_n737), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n737), .B2(new_n827), .ZN(new_n829));
  XOR2_X1   g0629(.A(KEYINPUT102), .B(G143), .Z(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n790), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n784), .A2(new_n831), .B1(new_n832), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n834), .B2(new_n794), .C1(new_n800), .C2(new_n343), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT34), .Z(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n289), .B1(new_n786), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT103), .Z(new_n839));
  INV_X1    g0639(.A(new_n780), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G68), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n841), .B1(new_n813), .B2(new_n776), .C1(new_n229), .C2(new_n773), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n836), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n800), .A2(new_n779), .B1(new_n554), .B2(new_n790), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n845), .A2(KEYINPUT101), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(KEYINPUT101), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n397), .B1(new_n773), .B2(new_n525), .C1(new_n794), .C2(new_n564), .ZN(new_n848));
  INV_X1    g0648(.A(G294), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n783), .A2(new_n849), .B1(new_n786), .B2(new_n789), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n780), .A2(new_n225), .B1(new_n776), .B2(new_n473), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n846), .A2(new_n847), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n817), .B1(new_n844), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n762), .A2(new_n757), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n754), .B(new_n854), .C1(new_n202), .C2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT104), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n823), .A2(new_n757), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(KEYINPUT104), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n829), .B1(new_n860), .B2(new_n861), .ZN(G384));
  INV_X1    g0662(.A(new_n590), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n863), .A2(KEYINPUT35), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(KEYINPUT35), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n864), .A2(G116), .A3(new_n216), .A4(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT36), .Z(new_n867));
  OAI211_X1 g0667(.A(new_n218), .B(G77), .C1(new_n229), .C2(new_n231), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n813), .A2(G68), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n303), .B(G13), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n394), .A2(new_n406), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n412), .ZN(new_n873));
  INV_X1    g0673(.A(new_n675), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n622), .B2(new_n440), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n873), .B1(new_n437), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n421), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  INV_X1    g0679(.A(new_n631), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n675), .B(KEYINPUT105), .Z(new_n881));
  NAND2_X1  g0681(.A1(new_n429), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n880), .A2(new_n882), .A3(new_n883), .A4(new_n421), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT38), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT106), .B1(new_n876), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n882), .B1(new_n636), .B2(new_n425), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n880), .A2(new_n882), .A3(new_n421), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(new_n883), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n888), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  INV_X1    g0693(.A(new_n875), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n442), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT106), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT38), .A4(new_n885), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n887), .A2(new_n892), .A3(new_n893), .A4(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n895), .B2(new_n885), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n886), .B1(new_n442), .B2(new_n894), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT39), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n321), .A2(new_n677), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n822), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n668), .B2(new_n825), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n283), .A2(new_n677), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n321), .A2(new_n324), .A3(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n283), .B(new_n677), .C1(new_n318), .C2(new_n320), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n899), .A2(new_n900), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n913), .A2(new_n914), .B1(new_n636), .B2(new_n881), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n904), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n638), .B1(new_n748), .B2(new_n443), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n823), .B1(new_n908), .B2(new_n909), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n686), .B1(new_n719), .B2(new_n722), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT31), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n725), .A2(new_n731), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n919), .B1(new_n914), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n919), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n887), .A2(new_n892), .A3(new_n897), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n383), .A2(new_n442), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n923), .ZN(new_n931));
  OAI21_X1  g0731(.A(G330), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n929), .B2(new_n931), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n918), .A2(new_n933), .B1(new_n303), .B2(new_n752), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n918), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n871), .B1(new_n934), .B2(new_n935), .ZN(G367));
  AOI21_X1  g0736(.A(new_n764), .B1(new_n694), .B2(new_n372), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n244), .A2(new_n765), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n754), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n780), .A2(new_n202), .B1(new_n776), .B2(new_n229), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n289), .B1(new_n783), .B2(new_n343), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n940), .B(new_n941), .C1(new_n795), .C2(new_n831), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n773), .A2(new_n231), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n786), .A2(new_n834), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(new_n832), .C2(G50), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n942), .B(new_n945), .C1(new_n391), .C2(new_n800), .ZN(new_n946));
  INV_X1    g0746(.A(G317), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n397), .B1(new_n780), .B2(new_n525), .C1(new_n947), .C2(new_n786), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT108), .Z(new_n949));
  NAND3_X1  g0749(.A1(new_n777), .A2(KEYINPUT46), .A3(G116), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n794), .B2(new_n789), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n783), .A2(new_n564), .B1(new_n773), .B2(new_n473), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n790), .A2(new_n779), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT46), .B1(new_n777), .B2(G116), .ZN(new_n954));
  NOR4_X1   g0754(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n460), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n956), .B2(new_n800), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n946), .B1(new_n949), .B2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT47), .Z(new_n959));
  OR2_X1    g0759(.A1(new_n547), .A2(new_n686), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n660), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n663), .A2(new_n960), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n939), .B1(new_n817), .B2(new_n959), .C1(new_n964), .C2(new_n760), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n752), .A2(G45), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(G1), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n664), .A2(new_n677), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n666), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n639), .A2(new_n677), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n692), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT45), .Z(new_n973));
  NOR2_X1   g0773(.A1(new_n692), .A2(new_n971), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(new_n689), .Z(new_n977));
  NAND2_X1  g0777(.A1(new_n685), .A2(new_n691), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n688), .B2(new_n691), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n751), .B(new_n979), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n749), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n749), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n695), .B(KEYINPUT41), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n967), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT43), .B1(new_n963), .B2(KEYINPUT107), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(KEYINPUT107), .B2(new_n963), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n988));
  INV_X1    g0788(.A(new_n971), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n978), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT42), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n601), .B1(new_n969), .B2(new_n498), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n686), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n987), .A2(new_n988), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n987), .B2(new_n994), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n689), .A2(new_n989), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n996), .B(new_n997), .Z(new_n998));
  OAI21_X1  g0798(.A(new_n965), .B1(new_n985), .B2(new_n998), .ZN(G387));
  NAND2_X1  g0799(.A1(new_n980), .A2(new_n967), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n769), .A2(new_n698), .B1(new_n473), .B2(new_n694), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n241), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n765), .B1(new_n1002), .B2(new_n445), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n369), .A2(new_n813), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT50), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n445), .B1(new_n231), .B2(new_n202), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1005), .A2(new_n698), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1001), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n754), .B1(new_n1008), .B2(new_n763), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n795), .A2(G159), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT109), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n774), .A2(new_n372), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n343), .B2(new_n786), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n289), .B1(new_n780), .B2(new_n525), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n784), .A2(G50), .B1(G77), .B2(new_n777), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n231), .C2(new_n790), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n800), .A2(new_n345), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1011), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G317), .A2(new_n784), .B1(new_n832), .B2(G303), .ZN(new_n1020));
  INV_X1    g0820(.A(G322), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n794), .C1(new_n800), .C2(new_n789), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n774), .A2(G283), .B1(new_n777), .B2(new_n460), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n289), .B1(new_n787), .B2(G326), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n554), .B2(new_n780), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n1028), .B2(KEYINPUT49), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1019), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1009), .B1(new_n688), .B2(new_n760), .C1(new_n1033), .C2(new_n817), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n981), .A2(new_n695), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n980), .A2(new_n749), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1000), .B(new_n1034), .C1(new_n1035), .C2(new_n1036), .ZN(G393));
  OAI21_X1  g0837(.A(new_n763), .B1(new_n525), .B2(new_n206), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n251), .A2(new_n766), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n753), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n289), .B1(new_n780), .B2(new_n225), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n774), .A2(G77), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n231), .B2(new_n776), .C1(new_n786), .C2(new_n830), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(new_n369), .C2(new_n832), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n794), .A2(new_n343), .B1(new_n783), .B2(new_n391), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1044), .B(new_n1046), .C1(new_n813), .C2(new_n800), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT110), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n774), .A2(G116), .B1(new_n777), .B2(G283), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n849), .B2(new_n790), .C1(new_n1021), .C2(new_n786), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n289), .B(new_n1051), .C1(G107), .C2(new_n840), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n794), .A2(new_n947), .B1(new_n783), .B2(new_n789), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT52), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1052), .B(new_n1054), .C1(new_n564), .C2(new_n800), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1049), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1040), .B1(new_n1057), .B2(new_n762), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n760), .B2(new_n971), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n967), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n982), .A2(new_n695), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n977), .A2(new_n981), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1059), .B1(new_n1060), .B2(new_n977), .C1(new_n1061), .C2(new_n1062), .ZN(G390));
  INV_X1    g0863(.A(KEYINPUT111), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n903), .B1(new_n906), .B2(new_n911), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n898), .A2(new_n901), .A3(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n686), .B(new_n821), .C1(new_n740), .C2(new_n743), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n822), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n910), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n927), .A2(new_n1069), .A3(new_n903), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n920), .A2(new_n923), .A3(G330), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1064), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n923), .A2(G330), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n930), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(new_n638), .C1(new_n748), .C2(new_n443), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n906), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n823), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n910), .B1(new_n736), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1078), .B1(new_n1080), .B2(new_n1072), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n923), .A2(G330), .A3(new_n1079), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1068), .B1(new_n911), .B2(new_n1082), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n921), .A2(KEYINPUT98), .A3(KEYINPUT31), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n733), .B1(new_n730), .B2(new_n703), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n725), .B(new_n724), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1086), .A2(G330), .A3(new_n1079), .A4(new_n910), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1077), .B1(new_n1081), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1073), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT111), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1066), .A2(new_n1070), .A3(new_n1087), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1074), .A2(new_n1089), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1086), .A2(G330), .A3(new_n1079), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1072), .B1(new_n1094), .B2(new_n911), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1088), .B1(new_n1095), .B2(new_n906), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1077), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1092), .B1(new_n1090), .B2(KEYINPUT111), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1064), .B(new_n1073), .C1(new_n1066), .C2(new_n1070), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1093), .A2(new_n1101), .A3(new_n695), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n902), .A2(new_n757), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n754), .B1(new_n855), .B2(new_n345), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n783), .A2(new_n837), .B1(new_n773), .B2(new_n391), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT54), .B(G143), .Z(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT113), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1107), .A2(new_n832), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1105), .B(new_n1108), .C1(G128), .C2(new_n795), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n776), .A2(new_n343), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT115), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT53), .Z(new_n1112));
  AOI21_X1  g0912(.A(new_n397), .B1(new_n787), .B2(G125), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n813), .B2(new_n780), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT114), .Z(new_n1115));
  NAND2_X1  g0915(.A1(new_n801), .A2(G137), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1109), .A2(new_n1112), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1042), .A2(new_n397), .A3(new_n806), .A4(new_n841), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G283), .B2(new_n795), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n790), .A2(new_n525), .B1(new_n786), .B2(new_n849), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G116), .B2(new_n784), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(new_n473), .C2(new_n800), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1103), .B(new_n1104), .C1(new_n817), .C2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1074), .A2(new_n967), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1125), .A2(KEYINPUT112), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(KEYINPUT112), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1102), .B(new_n1124), .C1(new_n1126), .C2(new_n1127), .ZN(G378));
  NAND3_X1  g0928(.A1(new_n925), .A2(new_n928), .A3(G330), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT118), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT118), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n925), .A2(new_n928), .A3(new_n1131), .A4(G330), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n355), .A2(new_n360), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n348), .A2(new_n874), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT55), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1133), .B(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1130), .A2(new_n1132), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT119), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT119), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1130), .A2(new_n1141), .A3(new_n1132), .A4(new_n1138), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n916), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1140), .A2(new_n916), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT120), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1099), .A2(new_n1100), .A3(new_n1098), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n1077), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1093), .A2(KEYINPUT120), .A3(new_n1097), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n696), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1156), .B2(new_n1155), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(G33), .A2(G41), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT116), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G50), .B(new_n1161), .C1(new_n449), .C2(new_n397), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n943), .A2(G41), .A3(new_n289), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n202), .B2(new_n776), .C1(new_n473), .C2(new_n783), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G116), .B2(new_n795), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n790), .A2(new_n371), .B1(new_n229), .B2(new_n780), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G283), .B2(new_n787), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(new_n525), .C2(new_n800), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT58), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n795), .A2(G125), .B1(new_n1107), .B2(new_n777), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G128), .A2(new_n784), .B1(new_n832), .B2(G137), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n343), .C2(new_n773), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G132), .B2(new_n801), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1161), .B1(new_n391), .B2(new_n780), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G124), .B2(new_n787), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT59), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1178), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1170), .B1(new_n1169), .B2(new_n1168), .C1(new_n1176), .C2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n762), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n855), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n753), .C1(G50), .C2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1138), .B2(new_n757), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1149), .B2(new_n967), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1158), .A2(new_n1186), .ZN(G375));
  NAND3_X1  g0987(.A1(new_n1081), .A2(new_n1077), .A3(new_n1088), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n1098), .A3(new_n984), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G50), .A2(new_n774), .B1(new_n787), .B2(G128), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n391), .B2(new_n776), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n397), .B1(new_n840), .B2(G58), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n790), .B2(new_n343), .C1(new_n834), .C2(new_n783), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(G132), .C2(new_n795), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n801), .A2(new_n1107), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n784), .A2(G283), .B1(new_n787), .B2(G303), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n473), .B2(new_n790), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n397), .B1(new_n780), .B2(new_n202), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT122), .Z(new_n1199));
  OAI221_X1 g0999(.A(new_n1012), .B1(new_n525), .B2(new_n776), .C1(new_n794), .C2(new_n849), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n801), .A2(G116), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1194), .A2(new_n1195), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n753), .B1(G68), .B2(new_n1183), .C1(new_n1203), .C2(new_n817), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n911), .B2(new_n757), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n967), .B(KEYINPUT121), .Z(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1205), .B1(new_n1096), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1189), .A2(new_n1208), .ZN(G381));
  INV_X1    g1009(.A(G375), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT124), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(G378), .A2(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(G378), .A2(new_n1211), .ZN(new_n1213));
  OR2_X1    g1013(.A1(G387), .A2(G390), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT123), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1214), .A2(new_n1216), .A3(G381), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .A4(new_n1217), .ZN(G407));
  NAND2_X1  g1018(.A1(new_n676), .A2(G213), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .A4(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(new_n1221), .A3(G213), .ZN(G409));
  INV_X1    g1022(.A(KEYINPUT60), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1188), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1188), .A2(new_n1223), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n695), .A3(new_n1098), .A4(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1226), .A2(new_n1208), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(G384), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(G384), .A3(new_n1208), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1229), .A2(KEYINPUT126), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT126), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1228), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1147), .A2(new_n1148), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n695), .B1(new_n1234), .B2(KEYINPUT57), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1149), .A2(KEYINPUT57), .A3(new_n1154), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G378), .B(new_n1186), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1151), .A2(new_n1150), .A3(new_n1077), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT120), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n984), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1240), .A2(new_n1206), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1213), .B(new_n1212), .C1(new_n1241), .C2(new_n1185), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT125), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1237), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1219), .B(new_n1233), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT63), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1237), .A2(new_n1242), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n1219), .A3(new_n1233), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(new_n1247), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G387), .A2(G390), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1214), .A2(new_n1252), .ZN(new_n1253));
  XOR2_X1   g1053(.A(G393), .B(G396), .Z(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1254), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1214), .A2(new_n1257), .A3(new_n1252), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1251), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT127), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1261), .B(new_n1219), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1220), .A2(G2897), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1232), .B(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1249), .A2(KEYINPUT125), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1237), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1261), .B1(new_n1268), .B2(new_n1219), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1248), .B(new_n1260), .C1(new_n1265), .C2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1255), .A2(new_n1258), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1246), .A2(KEYINPUT62), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1249), .A2(new_n1219), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT61), .B1(new_n1273), .B2(new_n1264), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1271), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1270), .A2(new_n1277), .ZN(G405));
  NAND3_X1  g1078(.A1(G375), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1237), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(new_n1255), .A3(new_n1258), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1271), .A3(new_n1237), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1232), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1281), .A2(new_n1233), .A3(new_n1282), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(G402));
endmodule


