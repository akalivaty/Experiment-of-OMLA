

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743;

  BUF_X1 U375 ( .A(n646), .Z(n352) );
  XNOR2_X1 U376 ( .A(n558), .B(n405), .ZN(n646) );
  XNOR2_X1 U377 ( .A(n500), .B(n499), .ZN(n724) );
  XNOR2_X1 U378 ( .A(n425), .B(n716), .ZN(n497) );
  XNOR2_X1 U379 ( .A(G119), .B(G128), .ZN(n507) );
  XNOR2_X2 U380 ( .A(n489), .B(KEYINPUT4), .ZN(n500) );
  XOR2_X1 U381 ( .A(G146), .B(G125), .Z(n353) );
  OR2_X2 U382 ( .A1(n384), .A2(KEYINPUT34), .ZN(n410) );
  NOR2_X2 U383 ( .A1(n568), .A2(n567), .ZN(n372) );
  XNOR2_X2 U384 ( .A(n592), .B(n593), .ZN(n383) );
  XNOR2_X2 U385 ( .A(n422), .B(KEYINPUT104), .ZN(n743) );
  XNOR2_X2 U386 ( .A(n427), .B(G101), .ZN(n382) );
  NOR2_X1 U387 ( .A1(n384), .A2(n395), .ZN(n368) );
  INV_X1 U388 ( .A(KEYINPUT25), .ZN(n515) );
  NOR2_X1 U389 ( .A1(n699), .A2(n707), .ZN(n394) );
  NOR2_X1 U390 ( .A1(n615), .A2(n707), .ZN(n403) );
  NOR2_X1 U391 ( .A1(n685), .A2(n707), .ZN(n393) );
  NOR2_X1 U392 ( .A1(n708), .A2(n666), .ZN(n671) );
  XNOR2_X1 U393 ( .A(n538), .B(n434), .ZN(n742) );
  XNOR2_X1 U394 ( .A(n368), .B(n365), .ZN(n590) );
  XNOR2_X1 U395 ( .A(n378), .B(n364), .ZN(n675) );
  OR2_X1 U396 ( .A1(n636), .A2(n377), .ZN(n378) );
  NOR2_X1 U397 ( .A1(n646), .A2(n645), .ZN(n598) );
  XNOR2_X1 U398 ( .A(n532), .B(KEYINPUT103), .ZN(n637) );
  XNOR2_X1 U399 ( .A(n444), .B(n443), .ZN(n544) );
  XNOR2_X1 U400 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U401 ( .A1(G902), .A2(n705), .ZN(n518) );
  XNOR2_X1 U402 ( .A(n513), .B(n512), .ZN(n705) );
  XNOR2_X1 U403 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U404 ( .A(n724), .B(n501), .ZN(n381) );
  XNOR2_X1 U405 ( .A(G116), .B(G113), .ZN(n376) );
  INV_X4 U406 ( .A(KEYINPUT66), .ZN(n427) );
  INV_X1 U407 ( .A(n587), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n518), .B(n517), .ZN(n649) );
  XNOR2_X1 U409 ( .A(n386), .B(n366), .ZN(n735) );
  BUF_X1 U410 ( .A(n737), .Z(n355) );
  XNOR2_X1 U411 ( .A(n414), .B(n455), .ZN(n737) );
  BUF_X1 U412 ( .A(n694), .Z(n703) );
  XNOR2_X1 U413 ( .A(n385), .B(n539), .ZN(n433) );
  NAND2_X1 U414 ( .A1(n735), .A2(n742), .ZN(n385) );
  XNOR2_X1 U415 ( .A(n375), .B(n373), .ZN(n522) );
  XNOR2_X1 U416 ( .A(n374), .B(G119), .ZN(n373) );
  XNOR2_X1 U417 ( .A(n376), .B(n490), .ZN(n375) );
  INV_X1 U418 ( .A(KEYINPUT3), .ZN(n374) );
  XNOR2_X1 U419 ( .A(n498), .B(G134), .ZN(n499) );
  XNOR2_X1 U420 ( .A(n467), .B(G475), .ZN(n443) );
  OR2_X1 U421 ( .A1(n696), .A2(G902), .ZN(n444) );
  OR2_X1 U422 ( .A1(n612), .A2(G902), .ZN(n416) );
  NOR2_X1 U423 ( .A1(n690), .A2(G902), .ZN(n406) );
  NAND2_X1 U424 ( .A1(n637), .A2(n396), .ZN(n395) );
  INV_X1 U425 ( .A(n616), .ZN(n448) );
  OR2_X2 U426 ( .A1(n737), .A2(KEYINPUT44), .ZN(n594) );
  INV_X1 U427 ( .A(KEYINPUT82), .ZN(n474) );
  XNOR2_X1 U428 ( .A(n372), .B(KEYINPUT48), .ZN(n371) );
  INV_X1 U429 ( .A(n534), .ZN(n432) );
  XNOR2_X1 U430 ( .A(n522), .B(n388), .ZN(n387) );
  XNOR2_X1 U431 ( .A(n457), .B(n389), .ZN(n388) );
  XNOR2_X1 U432 ( .A(n424), .B(n423), .ZN(n716) );
  INV_X1 U433 ( .A(G104), .ZN(n423) );
  XNOR2_X1 U434 ( .A(G107), .B(G110), .ZN(n424) );
  XNOR2_X1 U435 ( .A(n470), .B(n469), .ZN(n506) );
  XNOR2_X1 U436 ( .A(KEYINPUT8), .B(KEYINPUT68), .ZN(n468) );
  XOR2_X1 U437 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n459) );
  XNOR2_X1 U438 ( .A(G143), .B(G104), .ZN(n458) );
  XNOR2_X1 U439 ( .A(n437), .B(n435), .ZN(n461) );
  XNOR2_X1 U440 ( .A(n460), .B(n436), .ZN(n435) );
  XNOR2_X1 U441 ( .A(n439), .B(n438), .ZN(n437) );
  INV_X1 U442 ( .A(G122), .ZN(n436) );
  XOR2_X1 U443 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n464) );
  XNOR2_X1 U444 ( .A(n382), .B(n426), .ZN(n425) );
  INV_X1 U445 ( .A(KEYINPUT73), .ZN(n426) );
  INV_X1 U446 ( .A(G146), .ZN(n501) );
  NAND2_X1 U447 ( .A1(n611), .A2(n610), .ZN(n440) );
  XNOR2_X1 U448 ( .A(n400), .B(n399), .ZN(n576) );
  INV_X1 U449 ( .A(KEYINPUT39), .ZN(n399) );
  NOR2_X1 U450 ( .A1(n546), .A2(n636), .ZN(n400) );
  AND2_X1 U451 ( .A1(n413), .A2(n585), .ZN(n412) );
  NOR2_X1 U452 ( .A1(n536), .A2(n560), .ZN(n392) );
  BUF_X1 U453 ( .A(n652), .Z(n398) );
  XNOR2_X1 U454 ( .A(n652), .B(n559), .ZN(n390) );
  INV_X1 U455 ( .A(KEYINPUT1), .ZN(n405) );
  NOR2_X1 U456 ( .A1(G952), .A2(n727), .ZN(n707) );
  INV_X1 U457 ( .A(KEYINPUT72), .ZN(n490) );
  OR2_X1 U458 ( .A1(G237), .A2(G902), .ZN(n519) );
  XOR2_X1 U459 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n523) );
  INV_X1 U460 ( .A(KEYINPUT74), .ZN(n450) );
  AND2_X1 U461 ( .A1(n521), .A2(G214), .ZN(n439) );
  XNOR2_X1 U462 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n438) );
  XNOR2_X1 U463 ( .A(G113), .B(G131), .ZN(n460) );
  XNOR2_X1 U464 ( .A(G902), .B(KEYINPUT15), .ZN(n609) );
  XNOR2_X1 U465 ( .A(n370), .B(KEYINPUT86), .ZN(n451) );
  NOR2_X1 U466 ( .A1(n708), .A2(n609), .ZN(n370) );
  XOR2_X1 U467 ( .A(KEYINPUT77), .B(KEYINPUT17), .Z(n484) );
  XNOR2_X1 U468 ( .A(KEYINPUT78), .B(KEYINPUT92), .ZN(n483) );
  XNOR2_X1 U469 ( .A(n497), .B(n454), .ZN(n453) );
  INV_X1 U470 ( .A(n648), .ZN(n396) );
  AND2_X1 U471 ( .A1(n371), .A2(n575), .ZN(n421) );
  XNOR2_X1 U472 ( .A(KEYINPUT16), .B(G122), .ZN(n491) );
  XNOR2_X1 U473 ( .A(G116), .B(G134), .ZN(n471) );
  XOR2_X1 U474 ( .A(G107), .B(G122), .Z(n472) );
  INV_X1 U475 ( .A(KEYINPUT33), .ZN(n379) );
  NAND2_X1 U476 ( .A1(n598), .A2(n390), .ZN(n380) );
  BUF_X1 U477 ( .A(n574), .Z(n397) );
  NAND2_X1 U478 ( .A1(n431), .A2(n429), .ZN(n546) );
  XNOR2_X1 U479 ( .A(n430), .B(n363), .ZN(n429) );
  NOR2_X1 U480 ( .A1(n524), .A2(n432), .ZN(n431) );
  XNOR2_X1 U481 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U482 ( .A(n466), .B(n465), .ZN(n696) );
  XNOR2_X1 U483 ( .A(n381), .B(n356), .ZN(n690) );
  XNOR2_X1 U484 ( .A(n495), .B(n494), .ZN(n496) );
  INV_X1 U485 ( .A(G140), .ZN(n494) );
  XNOR2_X1 U486 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U487 ( .A1(n542), .A2(n675), .ZN(n538) );
  XNOR2_X1 U488 ( .A(n417), .B(KEYINPUT112), .ZN(n738) );
  XNOR2_X1 U489 ( .A(n419), .B(n566), .ZN(n418) );
  INV_X1 U490 ( .A(KEYINPUT36), .ZN(n566) );
  XNOR2_X1 U491 ( .A(n456), .B(KEYINPUT79), .ZN(n455) );
  INV_X1 U492 ( .A(KEYINPUT35), .ZN(n456) );
  XNOR2_X1 U493 ( .A(n599), .B(n367), .ZN(n630) );
  INV_X1 U494 ( .A(KEYINPUT31), .ZN(n367) );
  NOR2_X1 U495 ( .A1(n587), .A2(n398), .ZN(n586) );
  NAND2_X1 U496 ( .A1(n590), .A2(n361), .ZN(n616) );
  INV_X1 U497 ( .A(KEYINPUT63), .ZN(n402) );
  XNOR2_X1 U498 ( .A(n383), .B(n741), .ZN(G21) );
  NOR2_X2 U499 ( .A1(n542), .A2(n391), .ZN(n625) );
  XOR2_X1 U500 ( .A(n497), .B(n496), .Z(n356) );
  NOR2_X1 U501 ( .A1(n390), .A2(n354), .ZN(n357) );
  AND2_X1 U502 ( .A1(G210), .A2(n519), .ZN(n358) );
  NOR2_X1 U503 ( .A1(n390), .A2(n587), .ZN(n359) );
  AND2_X1 U504 ( .A1(n586), .A2(n352), .ZN(n360) );
  AND2_X1 U505 ( .A1(n357), .A2(n352), .ZN(n361) );
  AND2_X1 U506 ( .A1(n575), .A2(n608), .ZN(n362) );
  XOR2_X1 U507 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n363) );
  XOR2_X1 U508 ( .A(n533), .B(KEYINPUT110), .Z(n364) );
  XOR2_X1 U509 ( .A(KEYINPUT65), .B(KEYINPUT22), .Z(n365) );
  INV_X1 U510 ( .A(KEYINPUT34), .ZN(n415) );
  XOR2_X1 U511 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n366) );
  XNOR2_X1 U512 ( .A(n522), .B(n491), .ZN(n713) );
  NOR2_X1 U513 ( .A1(n618), .A2(n630), .ZN(n603) );
  XNOR2_X2 U514 ( .A(KEYINPUT97), .B(n602), .ZN(n618) );
  NAND2_X1 U515 ( .A1(n383), .A2(n743), .ZN(n595) );
  NAND2_X1 U516 ( .A1(n737), .A2(KEYINPUT44), .ZN(n597) );
  AND2_X2 U517 ( .A1(n369), .A2(n449), .ZN(n606) );
  NOR2_X1 U518 ( .A1(n445), .A2(n596), .ZN(n369) );
  NAND2_X1 U519 ( .A1(n371), .A2(n362), .ZN(n666) );
  NAND2_X1 U520 ( .A1(n637), .A2(n541), .ZN(n377) );
  NOR2_X1 U521 ( .A1(n636), .A2(n635), .ZN(n640) );
  XNOR2_X2 U522 ( .A(n380), .B(n379), .ZN(n674) );
  XNOR2_X1 U523 ( .A(n381), .B(n387), .ZN(n612) );
  XNOR2_X1 U524 ( .A(n382), .B(n523), .ZN(n389) );
  NOR2_X1 U525 ( .A1(n384), .A2(n657), .ZN(n599) );
  NOR2_X1 U526 ( .A1(n384), .A2(n398), .ZN(n600) );
  NAND2_X1 U527 ( .A1(n384), .A2(KEYINPUT34), .ZN(n413) );
  XNOR2_X2 U528 ( .A(n401), .B(n583), .ZN(n384) );
  NAND2_X1 U529 ( .A1(n576), .A2(n627), .ZN(n386) );
  AND2_X1 U530 ( .A1(n390), .A2(n561), .ZN(n562) );
  INV_X1 U531 ( .A(n428), .ZN(n391) );
  XNOR2_X2 U532 ( .A(n565), .B(KEYINPUT19), .ZN(n428) );
  NAND2_X1 U533 ( .A1(n590), .A2(n360), .ZN(n422) );
  XNOR2_X1 U534 ( .A(n392), .B(KEYINPUT28), .ZN(n537) );
  NAND2_X1 U535 ( .A1(n407), .A2(n412), .ZN(n414) );
  XNOR2_X1 U536 ( .A(n446), .B(KEYINPUT90), .ZN(n445) );
  NAND2_X1 U537 ( .A1(n569), .A2(n420), .ZN(n419) );
  XNOR2_X1 U538 ( .A(n393), .B(n686), .ZN(G51) );
  XNOR2_X1 U539 ( .A(n394), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X2 U540 ( .A1(n574), .A2(n541), .ZN(n565) );
  XNOR2_X2 U541 ( .A(n493), .B(n358), .ZN(n574) );
  NAND2_X1 U542 ( .A1(n694), .A2(G472), .ZN(n614) );
  NAND2_X2 U543 ( .A1(n441), .A2(n440), .ZN(n694) );
  NAND2_X1 U544 ( .A1(n428), .A2(n582), .ZN(n401) );
  XNOR2_X1 U545 ( .A(n403), .B(n402), .ZN(G57) );
  XNOR2_X1 U546 ( .A(n404), .B(n450), .ZN(n449) );
  NOR2_X2 U547 ( .A1(n595), .A2(n594), .ZN(n404) );
  XNOR2_X2 U548 ( .A(n406), .B(n502), .ZN(n558) );
  NAND2_X1 U549 ( .A1(n409), .A2(n408), .ZN(n407) );
  NAND2_X1 U550 ( .A1(n674), .A2(n415), .ZN(n408) );
  NAND2_X1 U551 ( .A1(n411), .A2(n410), .ZN(n409) );
  INV_X1 U552 ( .A(n674), .ZN(n411) );
  XNOR2_X2 U553 ( .A(n416), .B(G472), .ZN(n652) );
  NAND2_X1 U554 ( .A1(n418), .A2(n588), .ZN(n417) );
  INV_X1 U555 ( .A(n565), .ZN(n420) );
  NAND2_X1 U556 ( .A1(n421), .A2(n633), .ZN(n722) );
  NAND2_X1 U557 ( .A1(n652), .A2(n541), .ZN(n430) );
  NAND2_X1 U558 ( .A1(n597), .A2(n447), .ZN(n446) );
  NOR2_X1 U559 ( .A1(n671), .A2(n722), .ZN(n442) );
  NAND2_X1 U560 ( .A1(n442), .A2(n451), .ZN(n441) );
  NAND2_X1 U561 ( .A1(n433), .A2(n557), .ZN(n568) );
  INV_X1 U562 ( .A(KEYINPUT42), .ZN(n434) );
  NOR2_X1 U563 ( .A1(n605), .A2(n448), .ZN(n447) );
  XNOR2_X1 U564 ( .A(n452), .B(n492), .ZN(n680) );
  XNOR2_X1 U565 ( .A(n453), .B(n713), .ZN(n452) );
  INV_X1 U566 ( .A(n500), .ZN(n454) );
  XNOR2_X1 U567 ( .A(n684), .B(n683), .ZN(n685) );
  AND2_X1 U568 ( .A1(n521), .A2(G210), .ZN(n457) );
  XNOR2_X1 U569 ( .A(n612), .B(KEYINPUT62), .ZN(n613) );
  XNOR2_X1 U570 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U571 ( .A(n698), .B(n697), .ZN(n699) );
  XOR2_X2 U572 ( .A(G953), .B(KEYINPUT64), .Z(n727) );
  XNOR2_X1 U573 ( .A(n459), .B(n458), .ZN(n462) );
  NOR2_X1 U574 ( .A1(G953), .A2(G237), .ZN(n521) );
  XNOR2_X1 U575 ( .A(n462), .B(n461), .ZN(n466) );
  XNOR2_X1 U576 ( .A(n353), .B(G140), .ZN(n463) );
  XNOR2_X1 U577 ( .A(n464), .B(n463), .ZN(n723) );
  INV_X1 U578 ( .A(n723), .ZN(n465) );
  XNOR2_X1 U579 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n467) );
  XNOR2_X1 U580 ( .A(KEYINPUT101), .B(n544), .ZN(n540) );
  XNOR2_X1 U581 ( .A(KEYINPUT102), .B(G478), .ZN(n482) );
  NAND2_X1 U582 ( .A1(G234), .A2(n727), .ZN(n470) );
  XNOR2_X1 U583 ( .A(n468), .B(KEYINPUT69), .ZN(n469) );
  NAND2_X1 U584 ( .A1(G217), .A2(n506), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U586 ( .A(n473), .B(KEYINPUT7), .Z(n478) );
  XNOR2_X2 U587 ( .A(G143), .B(G128), .ZN(n475) );
  XNOR2_X2 U588 ( .A(n475), .B(n474), .ZN(n489) );
  INV_X1 U589 ( .A(n489), .ZN(n476) );
  XNOR2_X1 U590 ( .A(n476), .B(KEYINPUT9), .ZN(n477) );
  XNOR2_X1 U591 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U592 ( .A(n480), .B(n479), .ZN(n701) );
  NOR2_X1 U593 ( .A1(G902), .A2(n701), .ZN(n481) );
  XNOR2_X1 U594 ( .A(n482), .B(n481), .ZN(n545) );
  NAND2_X1 U595 ( .A1(n540), .A2(n545), .ZN(n564) );
  INV_X1 U596 ( .A(n564), .ZN(n627) );
  XNOR2_X1 U597 ( .A(n484), .B(n483), .ZN(n488) );
  XOR2_X1 U598 ( .A(n353), .B(KEYINPUT18), .Z(n486) );
  NAND2_X1 U599 ( .A1(G224), .A2(n727), .ZN(n485) );
  XNOR2_X1 U600 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U601 ( .A(n488), .B(n487), .Z(n492) );
  NAND2_X1 U602 ( .A1(n680), .A2(n609), .ZN(n493) );
  XNOR2_X1 U603 ( .A(n397), .B(KEYINPUT38), .ZN(n636) );
  NAND2_X1 U604 ( .A1(G227), .A2(n727), .ZN(n495) );
  XOR2_X1 U605 ( .A(G137), .B(G131), .Z(n498) );
  XNOR2_X1 U606 ( .A(KEYINPUT71), .B(G469), .ZN(n502) );
  XOR2_X1 U607 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n505) );
  NAND2_X1 U608 ( .A1(n609), .A2(G234), .ZN(n503) );
  XNOR2_X1 U609 ( .A(n503), .B(KEYINPUT20), .ZN(n514) );
  NAND2_X1 U610 ( .A1(G221), .A2(n514), .ZN(n504) );
  XNOR2_X1 U611 ( .A(n505), .B(n504), .ZN(n648) );
  XNOR2_X1 U612 ( .A(n723), .B(KEYINPUT24), .ZN(n513) );
  NAND2_X1 U613 ( .A1(G221), .A2(n506), .ZN(n511) );
  XOR2_X1 U614 ( .A(G110), .B(G137), .Z(n508) );
  XNOR2_X1 U615 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U616 ( .A(n509), .B(KEYINPUT23), .Z(n510) );
  NAND2_X1 U617 ( .A1(G217), .A2(n514), .ZN(n516) );
  NOR2_X1 U618 ( .A1(n648), .A2(n649), .ZN(n584) );
  AND2_X1 U619 ( .A1(n558), .A2(n584), .ZN(n601) );
  XNOR2_X1 U620 ( .A(n601), .B(KEYINPUT107), .ZN(n524) );
  NAND2_X1 U621 ( .A1(G214), .A2(n519), .ZN(n520) );
  XOR2_X1 U622 ( .A(KEYINPUT93), .B(n520), .Z(n541) );
  NAND2_X1 U623 ( .A1(G234), .A2(G237), .ZN(n525) );
  XNOR2_X1 U624 ( .A(n525), .B(KEYINPUT14), .ZN(n526) );
  XNOR2_X1 U625 ( .A(KEYINPUT76), .B(n526), .ZN(n528) );
  NAND2_X1 U626 ( .A1(G952), .A2(n528), .ZN(n664) );
  NOR2_X1 U627 ( .A1(G953), .A2(n664), .ZN(n527) );
  XOR2_X1 U628 ( .A(KEYINPUT94), .B(n527), .Z(n581) );
  NAND2_X1 U629 ( .A1(n528), .A2(G902), .ZN(n577) );
  NOR2_X1 U630 ( .A1(G900), .A2(n577), .ZN(n530) );
  INV_X1 U631 ( .A(n727), .ZN(n529) );
  NAND2_X1 U632 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U633 ( .A1(n581), .A2(n531), .ZN(n534) );
  XOR2_X1 U634 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n533) );
  INV_X1 U635 ( .A(n541), .ZN(n635) );
  NAND2_X1 U636 ( .A1(n545), .A2(n544), .ZN(n532) );
  INV_X1 U637 ( .A(n652), .ZN(n536) );
  INV_X1 U638 ( .A(n649), .ZN(n587) );
  NOR2_X1 U639 ( .A1(n648), .A2(n587), .ZN(n535) );
  NAND2_X1 U640 ( .A1(n535), .A2(n534), .ZN(n560) );
  NAND2_X1 U641 ( .A1(n537), .A2(n558), .ZN(n542) );
  XOR2_X1 U642 ( .A(KEYINPUT46), .B(KEYINPUT88), .Z(n539) );
  NOR2_X1 U643 ( .A1(n545), .A2(n540), .ZN(n629) );
  OR2_X1 U644 ( .A1(n627), .A2(n629), .ZN(n639) );
  NAND2_X1 U645 ( .A1(n639), .A2(n625), .ZN(n543) );
  NAND2_X1 U646 ( .A1(n543), .A2(KEYINPUT47), .ZN(n549) );
  NOR2_X1 U647 ( .A1(n545), .A2(n544), .ZN(n585) );
  INV_X1 U648 ( .A(n397), .ZN(n547) );
  NOR2_X1 U649 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U650 ( .A1(n585), .A2(n548), .ZN(n624) );
  NAND2_X1 U651 ( .A1(n549), .A2(n624), .ZN(n550) );
  XNOR2_X1 U652 ( .A(n550), .B(KEYINPUT84), .ZN(n556) );
  INV_X1 U653 ( .A(n625), .ZN(n554) );
  XNOR2_X1 U654 ( .A(KEYINPUT85), .B(n639), .ZN(n604) );
  XOR2_X1 U655 ( .A(KEYINPUT67), .B(KEYINPUT47), .Z(n551) );
  NOR2_X1 U656 ( .A1(n604), .A2(n551), .ZN(n552) );
  XNOR2_X1 U657 ( .A(KEYINPUT75), .B(n552), .ZN(n553) );
  NOR2_X1 U658 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U659 ( .A1(n556), .A2(n555), .ZN(n557) );
  INV_X1 U660 ( .A(KEYINPUT6), .ZN(n559) );
  INV_X1 U661 ( .A(n560), .ZN(n561) );
  XNOR2_X1 U662 ( .A(n562), .B(KEYINPUT105), .ZN(n563) );
  NOR2_X1 U663 ( .A1(n564), .A2(n563), .ZN(n569) );
  XNOR2_X1 U664 ( .A(n738), .B(KEYINPUT89), .ZN(n567) );
  XNOR2_X1 U665 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n572) );
  NAND2_X1 U666 ( .A1(n352), .A2(n569), .ZN(n570) );
  NOR2_X1 U667 ( .A1(n635), .A2(n570), .ZN(n571) );
  XNOR2_X1 U668 ( .A(n572), .B(n571), .ZN(n573) );
  NOR2_X1 U669 ( .A1(n397), .A2(n573), .ZN(n634) );
  INV_X1 U670 ( .A(n634), .ZN(n575) );
  NAND2_X1 U671 ( .A1(n629), .A2(n576), .ZN(n633) );
  INV_X1 U672 ( .A(n577), .ZN(n579) );
  INV_X1 U673 ( .A(G953), .ZN(n578) );
  NOR2_X1 U674 ( .A1(G898), .A2(n578), .ZN(n718) );
  NAND2_X1 U675 ( .A1(n579), .A2(n718), .ZN(n580) );
  NAND2_X1 U676 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U677 ( .A(KEYINPUT91), .B(KEYINPUT0), .Z(n583) );
  INV_X1 U678 ( .A(n584), .ZN(n645) );
  XNOR2_X1 U679 ( .A(KEYINPUT80), .B(KEYINPUT32), .ZN(n593) );
  INV_X1 U680 ( .A(n352), .ZN(n588) );
  NAND2_X1 U681 ( .A1(n359), .A2(n588), .ZN(n589) );
  XNOR2_X1 U682 ( .A(n589), .B(KEYINPUT81), .ZN(n591) );
  NAND2_X1 U683 ( .A1(n591), .A2(n590), .ZN(n592) );
  AND2_X1 U684 ( .A1(n595), .A2(KEYINPUT44), .ZN(n596) );
  NAND2_X1 U685 ( .A1(n398), .A2(n598), .ZN(n657) );
  NAND2_X1 U686 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X2 U688 ( .A(n606), .B(KEYINPUT45), .ZN(n708) );
  NAND2_X1 U689 ( .A1(KEYINPUT2), .A2(n633), .ZN(n607) );
  XNOR2_X1 U690 ( .A(KEYINPUT83), .B(n607), .ZN(n608) );
  INV_X1 U691 ( .A(n671), .ZN(n611) );
  INV_X1 U692 ( .A(KEYINPUT2), .ZN(n670) );
  NOR2_X1 U693 ( .A1(n609), .A2(n670), .ZN(n610) );
  XNOR2_X1 U694 ( .A(G101), .B(n616), .ZN(G3) );
  NAND2_X1 U695 ( .A1(n618), .A2(n627), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n617), .B(G104), .ZN(G6) );
  XOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n620) );
  NAND2_X1 U698 ( .A1(n618), .A2(n629), .ZN(n619) );
  XNOR2_X1 U699 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U700 ( .A(G107), .B(n621), .ZN(G9) );
  XOR2_X1 U701 ( .A(G128), .B(KEYINPUT29), .Z(n623) );
  NAND2_X1 U702 ( .A1(n625), .A2(n629), .ZN(n622) );
  XNOR2_X1 U703 ( .A(n623), .B(n622), .ZN(G30) );
  XNOR2_X1 U704 ( .A(G143), .B(n624), .ZN(G45) );
  NAND2_X1 U705 ( .A1(n625), .A2(n627), .ZN(n626) );
  XNOR2_X1 U706 ( .A(n626), .B(G146), .ZN(G48) );
  NAND2_X1 U707 ( .A1(n630), .A2(n627), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n628), .B(G113), .ZN(G15) );
  XOR2_X1 U709 ( .A(G116), .B(KEYINPUT113), .Z(n632) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U711 ( .A(n632), .B(n631), .ZN(G18) );
  XNOR2_X1 U712 ( .A(G134), .B(n633), .ZN(G36) );
  XOR2_X1 U713 ( .A(G140), .B(n634), .Z(G42) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U718 ( .A(KEYINPUT116), .B(n643), .Z(n644) );
  NOR2_X1 U719 ( .A1(n674), .A2(n644), .ZN(n661) );
  NAND2_X1 U720 ( .A1(n352), .A2(n645), .ZN(n647) );
  XNOR2_X1 U721 ( .A(KEYINPUT50), .B(n647), .ZN(n655) );
  XOR2_X1 U722 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n651) );
  NAND2_X1 U723 ( .A1(n354), .A2(n648), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(n653) );
  NOR2_X1 U725 ( .A1(n653), .A2(n398), .ZN(n654) );
  NAND2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U728 ( .A(KEYINPUT51), .B(n658), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n675), .A2(n659), .ZN(n660) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT52), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(KEYINPUT117), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n722), .A2(n708), .ZN(n667) );
  NAND2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n673) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n678) );
  NOR2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U740 ( .A1(G953), .A2(n676), .ZN(n677) );
  NAND2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U742 ( .A(KEYINPUT53), .B(n679), .Z(G75) );
  NAND2_X1 U743 ( .A1(n694), .A2(G210), .ZN(n684) );
  INV_X1 U744 ( .A(n680), .ZN(n682) );
  XOR2_X1 U745 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n681) );
  XOR2_X1 U746 ( .A(KEYINPUT87), .B(KEYINPUT56), .Z(n686) );
  XOR2_X1 U747 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n688) );
  XNOR2_X1 U748 ( .A(KEYINPUT119), .B(KEYINPUT118), .ZN(n687) );
  XNOR2_X1 U749 ( .A(n688), .B(n687), .ZN(n689) );
  XOR2_X1 U750 ( .A(n690), .B(n689), .Z(n692) );
  NAND2_X1 U751 ( .A1(n703), .A2(G469), .ZN(n691) );
  XNOR2_X1 U752 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U753 ( .A1(n707), .A2(n693), .ZN(G54) );
  NAND2_X1 U754 ( .A1(n694), .A2(G475), .ZN(n698) );
  XOR2_X1 U755 ( .A(KEYINPUT59), .B(KEYINPUT120), .Z(n695) );
  NAND2_X1 U756 ( .A1(G478), .A2(n703), .ZN(n700) );
  XNOR2_X1 U757 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U758 ( .A1(n707), .A2(n702), .ZN(G63) );
  NAND2_X1 U759 ( .A1(G217), .A2(n703), .ZN(n704) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U761 ( .A1(n707), .A2(n706), .ZN(G66) );
  OR2_X1 U762 ( .A1(G953), .A2(n708), .ZN(n712) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n709) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n709), .ZN(n710) );
  NAND2_X1 U765 ( .A1(n710), .A2(G898), .ZN(n711) );
  NAND2_X1 U766 ( .A1(n712), .A2(n711), .ZN(n721) );
  XNOR2_X1 U767 ( .A(G101), .B(n713), .ZN(n714) );
  XNOR2_X1 U768 ( .A(n714), .B(KEYINPUT122), .ZN(n715) );
  XOR2_X1 U769 ( .A(n716), .B(n715), .Z(n717) );
  NOR2_X1 U770 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U771 ( .A(KEYINPUT121), .B(n719), .Z(n720) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(G69) );
  XNOR2_X1 U773 ( .A(KEYINPUT123), .B(n722), .ZN(n726) );
  XOR2_X1 U774 ( .A(n724), .B(n723), .Z(n729) );
  INV_X1 U775 ( .A(n729), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n726), .B(n725), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n728), .A2(n727), .ZN(n734) );
  XNOR2_X1 U778 ( .A(G227), .B(n729), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n730), .A2(G900), .ZN(n731) );
  XNOR2_X1 U780 ( .A(KEYINPUT124), .B(n731), .ZN(n732) );
  NAND2_X1 U781 ( .A1(n732), .A2(G953), .ZN(n733) );
  NAND2_X1 U782 ( .A1(n734), .A2(n733), .ZN(G72) );
  XNOR2_X1 U783 ( .A(n735), .B(G131), .ZN(n736) );
  XNOR2_X1 U784 ( .A(n736), .B(KEYINPUT126), .ZN(G33) );
  XOR2_X1 U785 ( .A(n355), .B(G122), .Z(G24) );
  XOR2_X1 U786 ( .A(KEYINPUT114), .B(KEYINPUT37), .Z(n740) );
  XNOR2_X1 U787 ( .A(n738), .B(G125), .ZN(n739) );
  XNOR2_X1 U788 ( .A(n740), .B(n739), .ZN(G27) );
  XOR2_X1 U789 ( .A(G119), .B(KEYINPUT125), .Z(n741) );
  XNOR2_X1 U790 ( .A(G137), .B(n742), .ZN(G39) );
  XNOR2_X1 U791 ( .A(n743), .B(G110), .ZN(G12) );
endmodule

