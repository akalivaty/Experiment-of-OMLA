//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(G110), .B(G122), .Z(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT78), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n194), .A3(KEYINPUT78), .A4(new_n195), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(G101), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT4), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT79), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n191), .A2(new_n194), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(KEYINPUT80), .A3(new_n206), .A4(new_n195), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n191), .A2(new_n194), .A3(new_n206), .A4(new_n195), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n198), .A2(G101), .A3(new_n202), .A4(new_n199), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G116), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT2), .B(G113), .ZN(new_n219));
  XOR2_X1   g033(.A(new_n218), .B(new_n219), .Z(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n213), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n218), .A2(new_n219), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G113), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n226));
  INV_X1    g040(.A(new_n215), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n218), .A2(new_n226), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n224), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n193), .A2(G104), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n206), .B1(new_n195), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n208), .A2(new_n209), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n208), .A2(new_n209), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT82), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n207), .A2(new_n210), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n234), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n231), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n189), .B1(new_n222), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n231), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n240), .B1(new_n239), .B2(new_n234), .ZN(new_n245));
  AOI211_X1 g059(.A(KEYINPUT82), .B(new_n233), .C1(new_n207), .C2(new_n210), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n213), .A2(new_n221), .ZN(new_n248));
  INV_X1    g062(.A(new_n189), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n243), .A2(KEYINPUT6), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G143), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G143), .B(G146), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT0), .B(G128), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G125), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n255), .ZN(new_n262));
  INV_X1    g076(.A(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G125), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n252), .A2(KEYINPUT1), .A3(G146), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n263), .A2(KEYINPUT1), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n253), .A3(new_n255), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n264), .A2(new_n265), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G953), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G224), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n270), .B(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n275), .B(new_n189), .C1(new_n222), .C2(new_n242), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n251), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT86), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT5), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n223), .B1(new_n228), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n237), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n233), .B1(new_n207), .B2(new_n210), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(new_n231), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n189), .B(KEYINPUT8), .Z(new_n285));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n270), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n261), .A2(new_n269), .A3(KEYINPUT85), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n272), .A4(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n261), .A2(new_n269), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n290), .B(KEYINPUT85), .C1(new_n291), .C2(new_n273), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n284), .A2(new_n285), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n250), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n278), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI211_X1 g110(.A(KEYINPUT86), .B(G902), .C1(new_n293), .C2(new_n250), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n277), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G210), .B1(G237), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n299), .B(new_n277), .C1(new_n296), .C2(new_n297), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n188), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G952), .ZN(new_n304));
  AOI211_X1 g118(.A(G953), .B(new_n304), .C1(G234), .C2(G237), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT69), .B(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI211_X1 g122(.A(new_n271), .B(new_n308), .C1(G234), .C2(G237), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(KEYINPUT21), .B(G898), .Z(new_n311));
  OAI21_X1  g125(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n252), .A2(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n263), .A2(G143), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT93), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT93), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G134), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n316), .A2(G134), .A3(new_n318), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G122), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n324), .A2(KEYINPUT91), .A3(G116), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT91), .B1(new_n324), .B2(G116), .ZN(new_n326));
  OAI22_X1  g140(.A1(new_n325), .A2(new_n326), .B1(G116), .B2(new_n324), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n327), .A2(G107), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n324), .A2(KEYINPUT14), .A3(G116), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT94), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT14), .B1(new_n324), .B2(G116), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n325), .B2(new_n326), .ZN(new_n332));
  OAI21_X1  g146(.A(G107), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n323), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n327), .B(G107), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT13), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n313), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT92), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT92), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n313), .A2(new_n339), .A3(new_n336), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n314), .A3(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n313), .A2(new_n336), .ZN(new_n342));
  OAI21_X1  g156(.A(G134), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n335), .A2(new_n321), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n334), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT9), .B(G234), .Z(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G217), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n347), .A2(new_n348), .A3(G953), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n334), .A2(new_n344), .A3(new_n349), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G478), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n354), .A2(KEYINPUT15), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n308), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n353), .B2(new_n308), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT89), .ZN(new_n360));
  NOR2_X1   g174(.A1(G237), .A2(G953), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G143), .A3(G214), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(G143), .B1(new_n361), .B2(G214), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT18), .B(G131), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G140), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G125), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n265), .A2(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G146), .ZN(new_n370));
  XNOR2_X1  g184(.A(G125), .B(G140), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n254), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n364), .ZN(new_n374));
  NAND2_X1  g188(.A1(KEYINPUT18), .A2(G131), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n362), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n365), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT88), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT88), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n365), .A2(new_n376), .A3(new_n373), .A4(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT16), .ZN(new_n381));
  OR3_X1    g195(.A1(new_n265), .A2(KEYINPUT16), .A3(G140), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G146), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT73), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n265), .A2(KEYINPUT16), .A3(G140), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n371), .B2(KEYINPUT16), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT73), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G146), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n371), .B(KEYINPUT19), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n384), .A2(new_n388), .B1(new_n389), .B2(new_n254), .ZN(new_n390));
  OAI21_X1  g204(.A(G131), .B1(new_n363), .B2(new_n364), .ZN(new_n391));
  INV_X1    g205(.A(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n374), .A2(new_n392), .A3(new_n362), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n378), .A2(new_n380), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n190), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n360), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n378), .A2(new_n380), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n390), .A2(new_n394), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n397), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(KEYINPUT89), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(G146), .B1(new_n381), .B2(new_n382), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT17), .B(G131), .C1(new_n363), .C2(new_n364), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n383), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT90), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT90), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n405), .A2(new_n406), .A3(new_n409), .A4(new_n383), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n408), .B(new_n410), .C1(KEYINPUT17), .C2(new_n394), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n399), .A3(new_n397), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n398), .A2(new_n403), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G475), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n295), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n413), .A2(new_n418), .A3(new_n414), .A4(new_n295), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n411), .A2(new_n399), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n402), .ZN(new_n422));
  AOI21_X1  g236(.A(G902), .B1(new_n422), .B2(new_n412), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n423), .A2(new_n414), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n303), .A2(new_n312), .A3(new_n359), .A4(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n268), .B(new_n266), .C1(G128), .C2(new_n258), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT66), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT66), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n264), .A2(new_n429), .A3(new_n266), .A4(new_n268), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n320), .A2(G137), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n320), .A2(G137), .ZN(new_n434));
  OAI21_X1  g248(.A(G131), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT11), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n320), .B2(G137), .ZN(new_n437));
  INV_X1    g251(.A(G137), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT11), .A3(G134), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n437), .A2(new_n439), .A3(new_n392), .A4(new_n432), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n432), .A3(new_n439), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G131), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n260), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n443), .A2(KEYINPUT30), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT65), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n260), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n440), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n257), .B(KEYINPUT65), .C1(new_n258), .C2(new_n259), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n442), .A2(new_n427), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(new_n221), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n361), .A2(G210), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT26), .B(G101), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n443), .A2(new_n220), .A3(new_n447), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT31), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT28), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n455), .A2(new_n221), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n446), .B1(new_n431), .B2(new_n442), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT28), .A3(new_n220), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n463), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT31), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n458), .A2(new_n475), .A3(new_n464), .A4(new_n465), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n467), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(G472), .A2(G902), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT32), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(KEYINPUT32), .A3(new_n478), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n469), .A2(new_n483), .A3(new_n470), .A4(new_n472), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT28), .B1(new_n471), .B2(new_n220), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT68), .B1(new_n471), .B2(new_n220), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT68), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n441), .B1(new_n428), .B2(new_n430), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n487), .B(new_n221), .C1(new_n488), .C2(new_n446), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n465), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n485), .B1(new_n490), .B2(KEYINPUT28), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n464), .B(new_n484), .C1(new_n491), .C2(new_n483), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n458), .A2(new_n465), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(new_n464), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n307), .B1(new_n494), .B2(new_n483), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G472), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n481), .B(new_n482), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n271), .A2(G221), .A3(G234), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT75), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n438), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(G137), .A3(new_n502), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(KEYINPUT72), .A2(G110), .ZN(new_n507));
  NOR2_X1   g321(.A1(KEYINPUT72), .A2(G110), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n263), .B(G119), .C1(KEYINPUT71), .C2(KEYINPUT23), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT23), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n214), .B2(G128), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n214), .B2(G128), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n509), .B(new_n510), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n263), .A2(KEYINPUT70), .A3(G119), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n263), .A2(G119), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT70), .B1(new_n263), .B2(G119), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT24), .B(G110), .Z(new_n520));
  OAI21_X1  g334(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n387), .B1(new_n386), .B2(G146), .ZN(new_n522));
  AND4_X1   g336(.A1(new_n387), .A2(new_n381), .A3(G146), .A4(new_n382), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n521), .B(new_n372), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n519), .A2(new_n520), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G110), .ZN(new_n527));
  INV_X1    g341(.A(new_n383), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n525), .B(new_n527), .C1(new_n528), .C2(new_n404), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n524), .A2(KEYINPUT74), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT74), .B1(new_n524), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n506), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT76), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n504), .A2(new_n505), .A3(new_n529), .A4(new_n524), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT76), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n535), .B(new_n506), .C1(new_n530), .C2(new_n531), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n348), .B1(new_n308), .B2(G234), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n537), .A2(G902), .A3(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n533), .A2(new_n536), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n540), .A2(KEYINPUT25), .A3(new_n308), .A4(new_n534), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n533), .A2(new_n308), .A3(new_n534), .A4(new_n536), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n539), .B1(new_n545), .B2(new_n538), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n498), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G221), .B1(new_n347), .B2(G902), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n271), .A2(G227), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n549), .B(KEYINPUT77), .Z(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(G110), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(new_n366), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT10), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n428), .B2(new_n430), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n245), .B2(new_n246), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n427), .B(new_n234), .C1(new_n235), .C2(new_n236), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT81), .ZN(new_n559));
  INV_X1    g373(.A(new_n260), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n213), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT81), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(new_n562), .A3(new_n554), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n556), .A2(new_n559), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(new_n451), .ZN(new_n565));
  INV_X1    g379(.A(new_n451), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n238), .A2(new_n241), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n567), .A2(new_n555), .B1(new_n560), .B2(new_n213), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n557), .A2(new_n562), .A3(new_n554), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n562), .B1(new_n557), .B2(new_n554), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n566), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n553), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n427), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n237), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n557), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT12), .B1(new_n576), .B2(new_n451), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n578), .B(new_n566), .C1(new_n575), .C2(new_n557), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT83), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n568), .A2(new_n566), .A3(new_n571), .ZN(new_n581));
  INV_X1    g395(.A(new_n557), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n427), .B1(new_n239), .B2(new_n234), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n451), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n578), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT83), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n576), .A2(KEYINPUT12), .A3(new_n451), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n580), .A2(new_n581), .A3(new_n588), .A4(new_n552), .ZN(new_n589));
  AOI211_X1 g403(.A(G469), .B(new_n307), .C1(new_n573), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G469), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n577), .A2(new_n579), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n553), .B1(new_n565), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n564), .A2(new_n451), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n581), .A3(new_n552), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n591), .B1(new_n596), .B2(new_n295), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n548), .B1(new_n590), .B2(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n426), .A2(new_n547), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n206), .ZN(G3));
  AND2_X1   g414(.A1(new_n542), .A2(new_n543), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n542), .A2(new_n543), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n538), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n539), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n477), .A2(new_n308), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G472), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n479), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n598), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n353), .A2(new_n354), .A3(new_n308), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n352), .B2(KEYINPUT95), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n353), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n351), .B(new_n352), .C1(KEYINPUT95), .C2(new_n611), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n307), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n610), .B1(new_n615), .B2(new_n354), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n420), .B2(new_n424), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n303), .A2(new_n312), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT96), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT34), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(new_n190), .ZN(G6));
  NOR2_X1   g436(.A1(new_n423), .A2(new_n414), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n415), .A2(new_n416), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n359), .B(new_n623), .C1(new_n624), .C2(new_n417), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n303), .A2(new_n625), .A3(new_n312), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n609), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NOR2_X1   g444(.A1(new_n530), .A2(new_n531), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n506), .A2(KEYINPUT36), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n631), .B(new_n632), .Z(new_n633));
  NOR2_X1   g447(.A1(new_n538), .A2(G902), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n603), .A2(new_n635), .ZN(new_n636));
  OR4_X1    g450(.A1(new_n598), .A2(new_n426), .A3(new_n608), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT97), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  NAND2_X1  g454(.A1(new_n301), .A2(new_n302), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n187), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n497), .B1(new_n492), .B2(new_n495), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n477), .A2(KEYINPUT32), .A3(new_n478), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT32), .B1(new_n477), .B2(new_n478), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n636), .A2(new_n598), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n306), .B1(new_n310), .B2(G900), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n625), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n641), .B(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT38), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n493), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n463), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n490), .A2(new_n464), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n660), .A2(new_n295), .A3(new_n661), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n481), .B(new_n482), .C1(new_n662), .C2(new_n497), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT99), .Z(new_n664));
  INV_X1    g478(.A(new_n548), .ZN(new_n665));
  INV_X1    g479(.A(new_n597), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n573), .A2(new_n589), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n591), .A3(new_n308), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n665), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n649), .B(KEYINPUT100), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT39), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n359), .B1(new_n420), .B2(new_n424), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n636), .A2(new_n187), .A3(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n657), .A2(new_n664), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  NAND2_X1  g493(.A1(new_n617), .A2(new_n649), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n647), .A2(new_n648), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  NAND2_X1  g497(.A1(new_n667), .A2(new_n308), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n591), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n686), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n667), .A2(new_n308), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n687), .A2(new_n548), .A3(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n690), .A2(new_n646), .A3(new_n605), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n618), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT102), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT41), .B(G113), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  NAND2_X1  g509(.A1(new_n691), .A2(new_n627), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  AOI21_X1  g511(.A(new_n688), .B1(new_n667), .B2(new_n308), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n307), .B(new_n686), .C1(new_n573), .C2(new_n589), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n603), .A2(new_n635), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n498), .A2(new_n700), .A3(new_n548), .A4(new_n701), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(new_n426), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  OAI211_X1 g518(.A(new_n476), .B(new_n467), .C1(new_n491), .C2(new_n464), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n606), .A2(G472), .B1(new_n705), .B2(new_n478), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n700), .A2(new_n546), .A3(new_n548), .A4(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n641), .A2(new_n675), .A3(new_n187), .A4(new_n312), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n324), .ZN(G24));
  NOR2_X1   g524(.A1(new_n642), .A2(new_n690), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n617), .A2(new_n649), .A3(new_n706), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n701), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G125), .ZN(G27));
  NOR4_X1   g528(.A1(new_n646), .A2(new_n605), .A3(new_n641), .A4(new_n188), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(KEYINPUT42), .A3(new_n669), .A4(new_n681), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n641), .A2(new_n188), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n669), .A3(new_n546), .A4(new_n498), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n717), .B1(new_n719), .B2(new_n680), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G131), .ZN(G33));
  INV_X1    g536(.A(new_n547), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n669), .A3(new_n650), .A4(new_n718), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  NAND2_X1  g539(.A1(new_n420), .A2(new_n424), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n616), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n727), .A2(KEYINPUT43), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(KEYINPUT43), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n608), .B(new_n701), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(KEYINPUT44), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT103), .ZN(new_n733));
  INV_X1    g547(.A(new_n718), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n731), .B2(KEYINPUT44), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n596), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n593), .A2(KEYINPUT45), .A3(new_n595), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(G469), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n591), .A2(new_n295), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT46), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n590), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n741), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n745), .A2(new_n548), .A3(new_n671), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n733), .A2(new_n735), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT104), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G137), .ZN(G39));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n745), .B2(new_n548), .ZN(new_n751));
  AOI211_X1 g565(.A(KEYINPUT105), .B(new_n665), .C1(new_n743), .C2(new_n744), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n751), .B2(new_n752), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n734), .A2(new_n546), .A3(new_n498), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n754), .A2(new_n756), .A3(new_n681), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT106), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G140), .ZN(G42));
  NAND2_X1  g574(.A1(new_n754), .A2(new_n756), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n700), .A2(new_n665), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n305), .B1(new_n728), .B2(new_n729), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n706), .A2(new_n603), .A3(new_n604), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n718), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT114), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n654), .A2(KEYINPUT38), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n654), .A2(KEYINPUT38), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n769), .A2(new_n770), .A3(new_n187), .ZN(new_n771));
  INV_X1    g585(.A(new_n690), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(new_n766), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n718), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n764), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n764), .A2(new_n776), .A3(KEYINPUT116), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n701), .B(new_n706), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n771), .A2(new_n772), .A3(new_n766), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n664), .A2(new_n605), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n776), .A2(new_n306), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n425), .A3(new_n616), .A4(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n775), .A2(new_n781), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n734), .B1(new_n761), .B2(new_n762), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n790), .A3(new_n766), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n768), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n777), .B(new_n778), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n795), .B1(new_n796), .B2(new_n723), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT48), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n784), .A2(new_n617), .A3(new_n785), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(G952), .A3(new_n271), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n796), .A2(new_n795), .A3(new_n723), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT48), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n799), .B(new_n801), .C1(new_n803), .C2(new_n797), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n788), .A2(KEYINPUT117), .B1(new_n789), .B2(new_n766), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n793), .B1(new_n787), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n624), .A2(new_n417), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n359), .A3(new_n649), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n646), .A2(new_n810), .A3(new_n623), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n648), .B(new_n718), .C1(new_n811), .C2(new_n712), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT108), .B1(new_n812), .B2(new_n724), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(KEYINPUT108), .A3(new_n724), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n814), .A2(new_n815), .B1(new_n720), .B2(new_n716), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n303), .A2(new_n312), .A3(new_n617), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT107), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n303), .A2(KEYINPUT107), .A3(new_n312), .A4(new_n617), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n303), .A2(new_n312), .ZN(new_n821));
  INV_X1    g635(.A(new_n359), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n425), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n819), .B(new_n820), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n599), .B1(new_n824), .B2(new_n609), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n498), .A2(new_n700), .A3(new_n546), .A4(new_n548), .ZN(new_n826));
  OAI22_X1  g640(.A1(new_n426), .A2(new_n702), .B1(new_n826), .B2(new_n626), .ZN(new_n827));
  OAI22_X1  g641(.A1(new_n826), .A2(new_n817), .B1(new_n707), .B2(new_n708), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n825), .A2(new_n637), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n816), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n647), .B(new_n648), .C1(new_n650), .C2(new_n681), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n636), .A2(new_n663), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n303), .A2(new_n675), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n649), .B(KEYINPUT109), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n835), .A3(new_n669), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n833), .A2(new_n837), .A3(new_n713), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(KEYINPUT110), .B(KEYINPUT111), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n833), .A2(new_n837), .A3(KEYINPUT52), .A4(new_n713), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n840), .B(new_n841), .C1(KEYINPUT110), .C2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(KEYINPUT110), .B2(new_n842), .ZN(new_n844));
  INV_X1    g658(.A(new_n841), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n831), .A2(new_n832), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n840), .A2(new_n842), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n816), .A2(new_n830), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(KEYINPUT54), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n708), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n690), .A2(new_n765), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n691), .A2(new_n618), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n854), .A2(new_n855), .A3(new_n696), .A4(new_n703), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT112), .B1(new_n827), .B2(new_n828), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n721), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n856), .A2(new_n857), .A3(new_n721), .A4(KEYINPUT113), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n812), .A2(KEYINPUT108), .A3(new_n724), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT53), .B1(new_n863), .B2(new_n813), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n825), .A2(new_n637), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n862), .A2(new_n843), .A3(new_n846), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n849), .A2(new_n832), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n794), .A2(new_n808), .A3(new_n851), .A4(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n766), .A2(new_n711), .ZN(new_n872));
  OAI22_X1  g686(.A1(new_n871), .A2(new_n872), .B1(G952), .B2(G953), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n656), .A2(new_n548), .A3(new_n187), .A4(new_n727), .ZN(new_n874));
  INV_X1    g688(.A(new_n700), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(KEYINPUT49), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT49), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n546), .B1(new_n700), .B2(new_n877), .ZN(new_n878));
  OR4_X1    g692(.A1(new_n664), .A2(new_n874), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n879), .ZN(G75));
  NAND2_X1  g694(.A1(new_n251), .A2(new_n276), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n274), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT55), .Z(new_n883));
  AOI211_X1 g697(.A(new_n308), .B(new_n299), .C1(new_n867), .C2(new_n868), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(KEYINPUT56), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n867), .A2(new_n868), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n307), .A3(new_n300), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  INV_X1    g702(.A(new_n883), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n271), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n885), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n885), .A2(new_n890), .A3(KEYINPUT119), .A4(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(G51));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n308), .B(new_n739), .C1(new_n867), .C2(new_n868), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n740), .B(KEYINPUT57), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n867), .A2(new_n869), .A3(new_n868), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n869), .B1(new_n867), .B2(new_n868), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n903), .B2(new_n667), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n898), .B1(new_n904), .B2(new_n891), .ZN(new_n905));
  INV_X1    g719(.A(new_n667), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n870), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n908), .B2(new_n900), .ZN(new_n909));
  OAI211_X1 g723(.A(KEYINPUT120), .B(new_n892), .C1(new_n909), .C2(new_n899), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n910), .ZN(G54));
  NAND4_X1  g725(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .A4(new_n307), .ZN(new_n912));
  INV_X1    g726(.A(new_n413), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n912), .A2(new_n915), .A3(new_n913), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n912), .B2(new_n913), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n891), .B(new_n914), .C1(new_n916), .C2(new_n917), .ZN(G60));
  NAND2_X1  g732(.A1(new_n613), .A2(new_n614), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT122), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n851), .A2(new_n870), .ZN(new_n921));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT59), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n920), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n908), .A2(new_n920), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n891), .B(new_n924), .C1(new_n925), .C2(new_n923), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT60), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n886), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n633), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n892), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n933));
  OR2_X1    g747(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n929), .A2(new_n537), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n935), .ZN(new_n937));
  OAI211_X1 g751(.A(KEYINPUT123), .B(KEYINPUT61), .C1(new_n937), .C2(new_n931), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n936), .A2(new_n938), .ZN(G66));
  NOR2_X1   g753(.A1(new_n830), .A2(G953), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n271), .B1(new_n311), .B2(G224), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n881), .B1(G898), .B2(new_n271), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n942), .B(new_n943), .Z(G69));
  AND2_X1   g758(.A1(new_n448), .A2(new_n457), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(new_n389), .Z(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(G900), .B1(new_n947), .B2(G227), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n271), .B(new_n948), .C1(G227), .C2(new_n947), .ZN(new_n949));
  INV_X1    g763(.A(new_n833), .ZN(new_n950));
  INV_X1    g764(.A(new_n713), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT124), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n833), .A2(new_n953), .A3(new_n713), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n678), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(new_n747), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n823), .B1(new_n425), .B2(new_n616), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n715), .A2(new_n669), .A3(new_n671), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n759), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(G953), .B1(new_n961), .B2(new_n946), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n746), .A2(new_n723), .A3(new_n835), .ZN(new_n963));
  AND4_X1   g777(.A1(new_n747), .A2(new_n952), .A3(new_n954), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n721), .A2(new_n724), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT125), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n964), .A2(new_n759), .A3(new_n947), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n949), .B1(new_n962), .B2(new_n967), .ZN(G72));
  NAND4_X1  g782(.A1(new_n958), .A2(new_n759), .A3(new_n830), .A4(new_n960), .ZN(new_n969));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT63), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT126), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n660), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n494), .B(KEYINPUT127), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n964), .A2(new_n759), .A3(new_n830), .A4(new_n966), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n847), .A2(new_n850), .ZN(new_n977));
  NOR4_X1   g791(.A1(new_n977), .A2(new_n494), .A3(new_n659), .A4(new_n971), .ZN(new_n978));
  NOR4_X1   g792(.A1(new_n973), .A2(new_n976), .A3(new_n891), .A4(new_n978), .ZN(G57));
endmodule


