//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  OR3_X1    g0003(.A1(new_n203), .A2(KEYINPUT64), .A3(G13), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(new_n203), .B2(G13), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AOI22_X1  g0008(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(G58), .A2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n208), .B(new_n226), .C1(new_n229), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G264), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  AND2_X1   g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  OAI21_X1  g0050(.A(KEYINPUT66), .B1(new_n250), .B2(new_n227), .ZN(new_n251));
  AND2_X1   g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(G274), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n256), .A2(G244), .A3(new_n258), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n250), .A2(new_n227), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT67), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(KEYINPUT67), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G107), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n267), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n265), .A2(new_n266), .A3(new_n264), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT67), .B1(new_n270), .B2(new_n271), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G238), .A2(G1698), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(new_n217), .B2(G1698), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n263), .B(new_n274), .C1(new_n277), .C2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(G169), .B1(new_n262), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n282), .A2(new_n227), .ZN(new_n283));
  XOR2_X1   g0083(.A(KEYINPUT15), .B(G87), .Z(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT69), .B1(new_n269), .B2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(new_n228), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT8), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G58), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n216), .A2(KEYINPUT8), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n284), .A2(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G20), .A2(G77), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n283), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G1), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G20), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G77), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n283), .A2(new_n299), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT70), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n228), .B2(G1), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n257), .A2(KEYINPUT70), .A3(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n301), .A2(new_n305), .A3(new_n212), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n296), .A2(new_n300), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT71), .B1(new_n281), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  INV_X1    g0109(.A(new_n274), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n279), .B1(new_n267), .B2(new_n272), .ZN(new_n311));
  INV_X1    g0111(.A(new_n263), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n260), .A2(new_n261), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n300), .ZN(new_n316));
  INV_X1    g0116(.A(new_n306), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n294), .A2(new_n295), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n316), .B(new_n317), .C1(new_n318), .C2(new_n283), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n315), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n262), .A2(new_n322), .A3(new_n280), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n308), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n262), .A2(new_n280), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G200), .ZN(new_n326));
  INV_X1    g0126(.A(G190), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n326), .B(new_n307), .C1(new_n327), .C2(new_n325), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT72), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n259), .B1(new_n251), .B2(new_n255), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G226), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n267), .A2(new_n272), .ZN(new_n333));
  INV_X1    g0133(.A(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G222), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G223), .A2(G1698), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n263), .B1(new_n333), .B2(G77), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n260), .B(new_n332), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n309), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n337), .B(new_n263), .C1(G77), .C2(new_n333), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n342), .A2(new_n322), .A3(new_n260), .A4(new_n332), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n297), .A2(new_n228), .A3(G1), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n282), .A2(new_n227), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n346), .A2(G50), .A3(new_n304), .A4(new_n303), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n210), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n293), .A2(G150), .ZN(new_n349));
  NOR3_X1   g0149(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n228), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n216), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT8), .B(G58), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(KEYINPUT68), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n354), .B2(new_n288), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n347), .B(new_n348), .C1(new_n355), .C2(new_n283), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n341), .A2(new_n343), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n340), .A2(G200), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n355), .A2(new_n283), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n359), .A2(KEYINPUT9), .A3(new_n347), .A4(new_n348), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n342), .A2(G190), .A3(new_n260), .A4(new_n332), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT9), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n358), .A2(new_n360), .A3(new_n361), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT10), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n340), .A2(G200), .B1(new_n356), .B2(new_n362), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT10), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n360), .A4(new_n361), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n357), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n324), .A2(new_n370), .A3(new_n328), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n330), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT73), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n330), .A2(new_n369), .A3(KEYINPUT73), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT77), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT18), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n211), .A2(G1698), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n379), .B1(G223), .B2(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n380), .A2(KEYINPUT76), .A3(new_n381), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n263), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G274), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n251), .B2(new_n255), .ZN(new_n388));
  AOI22_X1  g0188(.A1(G232), .A2(new_n331), .B1(new_n388), .B2(new_n259), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G169), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(new_n389), .A3(G179), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n219), .A2(G58), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n231), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(G20), .B1(G159), .B2(new_n293), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  NOR4_X1   g0196(.A1(new_n265), .A2(new_n266), .A3(new_n396), .A4(G20), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n267), .A2(new_n272), .A3(new_n228), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(new_n396), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n395), .B1(new_n399), .B2(new_n220), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n265), .A2(new_n266), .A3(G20), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT75), .B1(new_n403), .B2(KEYINPUT7), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n270), .A2(new_n228), .A3(new_n271), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT75), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n396), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n397), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G68), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT16), .B(new_n395), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n402), .A2(new_n345), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n301), .A2(new_n305), .ZN(new_n412));
  MUX2_X1   g0212(.A(new_n344), .B(new_n412), .S(new_n354), .Z(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI221_X4 g0214(.A(new_n378), .B1(new_n391), .B2(new_n392), .C1(new_n411), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n414), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n391), .A2(new_n392), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT18), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n410), .A2(new_n345), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n413), .B1(new_n420), .B2(new_n402), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n390), .A2(G200), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n386), .A2(new_n389), .A3(G190), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n421), .A2(KEYINPUT17), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n411), .A2(new_n422), .A3(new_n423), .A4(new_n414), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n377), .B1(new_n419), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n391), .A2(new_n392), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n378), .B1(new_n421), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT18), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n433), .A2(KEYINPUT77), .A3(new_n427), .A4(new_n424), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT13), .ZN(new_n436));
  NOR2_X1   g0236(.A1(G226), .A2(G1698), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n334), .A2(G232), .ZN(new_n438));
  AOI211_X1 g0238(.A(new_n437), .B(new_n438), .C1(new_n267), .C2(new_n272), .ZN(new_n439));
  AND2_X1   g0239(.A1(G33), .A2(G97), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n263), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n256), .A2(G238), .A3(new_n258), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n260), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n436), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n437), .ZN(new_n445));
  INV_X1    g0245(.A(new_n438), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n446), .C1(new_n275), .C2(new_n276), .ZN(new_n447));
  INV_X1    g0247(.A(new_n440), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n312), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n260), .A2(new_n442), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT13), .ZN(new_n451));
  OAI21_X1  g0251(.A(G169), .B1(new_n444), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT14), .ZN(new_n453));
  OR3_X1    g0253(.A1(new_n444), .A2(new_n451), .A3(new_n322), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT14), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(G169), .C1(new_n444), .C2(new_n451), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT74), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n288), .A2(G77), .B1(G50), .B2(new_n293), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n220), .A2(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n283), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT12), .B1(new_n301), .B2(new_n305), .ZN(new_n463));
  AOI22_X1  g0263(.A1(KEYINPUT11), .A2(new_n462), .B1(new_n463), .B2(G68), .ZN(new_n464));
  OAI221_X1 g0264(.A(new_n464), .B1(KEYINPUT11), .B2(new_n462), .C1(KEYINPUT12), .C2(new_n344), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT12), .ZN(new_n466));
  INV_X1    g0266(.A(new_n298), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n461), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT74), .A4(new_n456), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n459), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n444), .A2(new_n451), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G200), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n469), .B(new_n474), .C1(new_n473), .C2(new_n327), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n376), .A2(new_n435), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT78), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n376), .A2(new_n435), .A3(new_n476), .A4(KEYINPUT78), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n267), .A2(new_n272), .A3(G303), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n270), .A2(new_n271), .ZN(new_n483));
  OR2_X1    g0283(.A1(G257), .A2(G1698), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n484), .C1(G264), .C2(new_n334), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n263), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n257), .A2(G45), .ZN(new_n488));
  OR2_X1    g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n251), .B2(new_n255), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G270), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n388), .A2(new_n491), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n487), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n346), .B(G116), .C1(G1), .C2(new_n269), .ZN(new_n496));
  INV_X1    g0296(.A(G116), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n344), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n282), .A2(new_n227), .B1(G20), .B2(new_n497), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  INV_X1    g0300(.A(G97), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n500), .B(new_n228), .C1(G33), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT20), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n499), .A2(KEYINPUT20), .A3(new_n502), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n496), .B(new_n498), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n495), .A2(G169), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT85), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n506), .B2(new_n507), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT86), .ZN(new_n512));
  INV_X1    g0312(.A(new_n495), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G179), .A3(new_n505), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n495), .A2(G200), .ZN(new_n515));
  INV_X1    g0315(.A(new_n505), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(new_n327), .C2(new_n495), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n511), .A2(new_n512), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n506), .A2(new_n507), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT21), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(new_n514), .A4(new_n517), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT86), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(KEYINPUT22), .B(G87), .C1(new_n265), .C2(new_n266), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n228), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n228), .A2(G107), .B1(KEYINPUT88), .B2(KEYINPUT23), .ZN(new_n529));
  AND2_X1   g0329(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n228), .A2(G87), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n267), .B2(new_n272), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n528), .B(new_n531), .C1(KEYINPUT22), .C2(new_n533), .ZN(new_n534));
  XNOR2_X1  g0334(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n277), .B2(new_n532), .ZN(new_n538));
  INV_X1    g0338(.A(new_n535), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n538), .A2(new_n539), .A3(new_n528), .A4(new_n531), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n345), .A3(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n283), .B(new_n299), .C1(G1), .C2(new_n269), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G107), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n298), .A2(G20), .A3(new_n273), .ZN(new_n546));
  XOR2_X1   g0346(.A(new_n546), .B(KEYINPUT25), .Z(new_n547));
  NAND2_X1  g0347(.A1(new_n223), .A2(new_n334), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n483), .B(new_n548), .C1(G257), .C2(new_n334), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G294), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(new_n263), .B1(new_n492), .B2(G264), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n494), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n327), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n545), .A2(new_n547), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n288), .A2(G97), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT82), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT81), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT81), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT19), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n558), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n501), .B1(new_n285), .B2(new_n287), .ZN(new_n566));
  INV_X1    g0366(.A(new_n564), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT82), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n561), .A2(new_n563), .A3(new_n440), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n228), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n222), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n483), .A2(new_n228), .A3(G68), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n565), .A2(new_n568), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n284), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n575), .A2(new_n345), .B1(new_n344), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n218), .A2(new_n334), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n483), .B(new_n578), .C1(G244), .C2(new_n334), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n526), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n263), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n488), .A2(KEYINPUT80), .A3(G250), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT80), .ZN(new_n583));
  AOI21_X1  g0383(.A(G274), .B1(new_n583), .B2(G250), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n582), .B1(new_n584), .B2(new_n488), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n256), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n543), .A2(G87), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n577), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n586), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n312), .B1(new_n579), .B2(new_n526), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT84), .B1(new_n593), .B2(G190), .ZN(new_n594));
  AND4_X1   g0394(.A1(KEYINPUT84), .A2(new_n581), .A3(G190), .A4(new_n586), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(G169), .B1(new_n581), .B2(new_n586), .ZN(new_n597));
  OR3_X1    g0397(.A1(new_n542), .A2(KEYINPUT83), .A3(new_n576), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT83), .B1(new_n542), .B2(new_n576), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n597), .B1(new_n577), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n593), .A2(new_n322), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n590), .A2(new_n596), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n541), .A2(new_n544), .A3(new_n547), .ZN(new_n604));
  AOI21_X1  g0404(.A(G169), .B1(new_n552), .B2(new_n494), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n551), .A2(new_n263), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n492), .A2(G264), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n494), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n605), .B1(new_n322), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n557), .A2(new_n603), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n293), .A2(G77), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n273), .A2(KEYINPUT6), .A3(G97), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n501), .A2(new_n273), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n571), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n617), .B2(KEYINPUT6), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G20), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n614), .B(new_n619), .C1(new_n399), .C2(new_n273), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n345), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n344), .A2(new_n501), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n542), .B2(new_n501), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT79), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n623), .B1(new_n620), .B2(new_n345), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT79), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n223), .B1(new_n267), .B2(new_n272), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT4), .ZN(new_n631));
  OAI21_X1  g0431(.A(G1698), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n213), .B1(new_n270), .B2(new_n271), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n500), .B1(new_n633), .B2(KEYINPUT4), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n213), .B1(new_n267), .B2(new_n272), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n631), .A2(G1698), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n632), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n609), .B1(new_n639), .B2(new_n263), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n492), .A2(G257), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n309), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n634), .B1(new_n637), .B2(new_n636), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n312), .B1(new_n643), .B2(new_n632), .ZN(new_n644));
  INV_X1    g0444(.A(new_n641), .ZN(new_n645));
  NOR4_X1   g0445(.A1(new_n644), .A2(new_n322), .A3(new_n609), .A4(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n627), .B(new_n629), .C1(new_n642), .C2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n640), .A2(G190), .A3(new_n641), .ZN(new_n648));
  INV_X1    g0448(.A(G200), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n644), .A2(new_n609), .A3(new_n645), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n648), .B(new_n628), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n613), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n481), .A2(new_n524), .A3(new_n653), .ZN(G372));
  INV_X1    g0454(.A(new_n324), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n475), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n472), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n433), .B1(new_n657), .B2(new_n428), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n365), .A2(new_n368), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n357), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n481), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n649), .B1(new_n640), .B2(new_n641), .ZN(new_n662));
  NOR4_X1   g0462(.A1(new_n644), .A2(new_n327), .A3(new_n609), .A4(new_n645), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT79), .B1(new_n621), .B2(new_n624), .ZN(new_n665));
  AOI211_X1 g0465(.A(new_n626), .B(new_n623), .C1(new_n620), .C2(new_n345), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n639), .A2(new_n263), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(G179), .A3(new_n494), .A4(new_n641), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n650), .B2(new_n309), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n628), .A2(new_n664), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT89), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n575), .A2(new_n345), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n576), .A2(new_n344), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n600), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n597), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n602), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n593), .A2(G190), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n577), .A2(new_n588), .A3(new_n678), .A4(new_n589), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n604), .A2(new_n555), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n554), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n671), .A2(new_n672), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n672), .B1(new_n671), .B2(new_n682), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT90), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n520), .A2(new_n521), .A3(new_n514), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n604), .A2(new_n611), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n511), .A2(KEYINPUT90), .A3(new_n514), .A4(new_n612), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n683), .A2(new_n684), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n625), .B1(new_n642), .B2(new_n646), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n680), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT91), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n603), .A2(KEYINPUT26), .A3(new_n670), .A4(new_n667), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT91), .B(new_n692), .C1(new_n693), .C2(new_n680), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n677), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n691), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n660), .B1(new_n661), .B2(new_n701), .ZN(G369));
  OR3_X1    g0502(.A1(new_n467), .A2(KEYINPUT27), .A3(G20), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT27), .B1(new_n467), .B2(G20), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT92), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G343), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n516), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n511), .B2(new_n514), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n524), .B2(new_n709), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT93), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n710), .A2(KEYINPUT93), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n707), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n612), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n604), .A2(new_n716), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n557), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n717), .B1(new_n719), .B2(new_n612), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n715), .A2(G330), .A3(new_n720), .ZN(new_n721));
  AND4_X1   g0521(.A1(new_n686), .A2(new_n557), .A3(new_n612), .A4(new_n707), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n717), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n206), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n726), .A2(G116), .A3(new_n572), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n727), .A2(G1), .B1(new_n233), .B2(new_n726), .ZN(new_n728));
  XNOR2_X1  g0528(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n731), .B(new_n707), .C1(new_n691), .C2(new_n700), .ZN(new_n732));
  INV_X1    g0532(.A(G330), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n640), .A2(G179), .A3(new_n513), .A4(new_n641), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n587), .A2(new_n608), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n646), .A2(KEYINPUT30), .A3(new_n513), .A4(new_n737), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n640), .A2(new_n641), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n513), .A2(new_n593), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n322), .A4(new_n553), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n740), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n734), .B1(new_n744), .B2(new_n716), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(new_n734), .A3(new_n716), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n653), .A2(new_n524), .A3(new_n707), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n733), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n671), .A2(new_n682), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n686), .A2(new_n687), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n603), .A2(new_n692), .A3(new_n670), .A4(new_n667), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT26), .B1(new_n693), .B2(new_n680), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(new_n756), .A3(new_n677), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n707), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT29), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n732), .A2(new_n751), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n730), .B1(new_n761), .B2(G1), .ZN(G364));
  NOR2_X1   g0562(.A1(new_n297), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n257), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n726), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n206), .A2(new_n333), .A3(G355), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n725), .A2(new_n483), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G45), .B2(new_n232), .ZN(new_n770));
  INV_X1    g0570(.A(G45), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n245), .A2(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n768), .B1(G116), .B2(new_n206), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT95), .Z(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n227), .B1(G20), .B2(new_n309), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n767), .B1(new_n773), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT96), .Z(new_n781));
  NOR2_X1   g0581(.A1(new_n228), .A2(new_n322), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n783), .A2(new_n649), .A3(G190), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n228), .A2(G179), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G190), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n784), .A2(new_n785), .B1(G329), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G303), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n327), .A2(new_n649), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n786), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n790), .B(new_n277), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n327), .A2(G179), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n228), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n794), .B1(G294), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n782), .A2(new_n792), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G326), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n783), .A2(new_n327), .A3(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n782), .A2(new_n787), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n802), .A2(G322), .B1(G311), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n798), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n786), .A2(new_n327), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT97), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n806), .B1(G283), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(G107), .ZN(new_n814));
  INV_X1    g0614(.A(G159), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n788), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT32), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n277), .B1(G50), .B2(new_n800), .ZN(new_n818));
  INV_X1    g0618(.A(new_n793), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G87), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n814), .A2(new_n817), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n796), .A2(new_n501), .ZN(new_n822));
  INV_X1    g0622(.A(new_n784), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n409), .ZN(new_n824));
  INV_X1    g0624(.A(new_n802), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n825), .A2(new_n216), .B1(new_n803), .B2(new_n212), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n821), .A2(new_n822), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n778), .B1(new_n813), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n777), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n781), .B(new_n828), .C1(new_n715), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n715), .A2(G330), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n713), .A2(new_n714), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n733), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n830), .B1(new_n834), .B2(new_n766), .ZN(G396));
  NOR2_X1   g0635(.A1(new_n707), .A2(new_n307), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n329), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n655), .A2(new_n836), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(new_n701), .C2(new_n716), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n707), .B(new_n840), .C1(new_n691), .C2(new_n700), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n751), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n839), .A2(new_n750), .A3(new_n841), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n767), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n811), .A2(new_n409), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n802), .A2(G143), .B1(G159), .B2(new_n804), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  INV_X1    g0648(.A(G150), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n847), .B1(new_n848), .B2(new_n799), .C1(new_n849), .C2(new_n823), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT34), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n483), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n846), .B(new_n852), .C1(new_n851), .C2(new_n850), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n216), .B2(new_n796), .C1(new_n854), .C2(new_n788), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G50), .B2(new_n819), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n799), .A2(new_n791), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n811), .A2(new_n222), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G311), .B2(new_n789), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT99), .Z(new_n860));
  AOI211_X1 g0660(.A(new_n333), .B(new_n822), .C1(G116), .C2(new_n804), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n784), .A2(G283), .B1(G107), .B2(new_n819), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n857), .B(new_n863), .C1(G294), .C2(new_n802), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n778), .B1(new_n856), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n778), .A2(new_n774), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n766), .B1(G77), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT98), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT100), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n776), .B2(new_n840), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n845), .A2(new_n872), .ZN(G384));
  NAND2_X1  g0673(.A1(new_n472), .A2(new_n475), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n469), .A2(new_n707), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n875), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n472), .A2(new_n475), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n748), .A2(new_n749), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n879), .A2(new_n880), .A3(new_n840), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n395), .B1(new_n408), .B2(new_n409), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n401), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(KEYINPUT102), .A3(new_n345), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n410), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT102), .B1(new_n883), .B2(new_n345), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n414), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n706), .B(new_n887), .C1(new_n419), .C2(new_n428), .ZN(new_n888));
  INV_X1    g0688(.A(new_n706), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n430), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n416), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n892), .A3(new_n425), .ZN(new_n893));
  INV_X1    g0693(.A(new_n425), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n887), .B2(new_n890), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n893), .B1(new_n895), .B2(new_n892), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n888), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n888), .A2(new_n896), .A3(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n881), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n891), .A2(new_n425), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n893), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n416), .B(new_n706), .C1(new_n419), .C2(new_n428), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n903), .B1(new_n909), .B2(new_n900), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n902), .A2(new_n903), .B1(new_n910), .B2(new_n881), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n481), .A2(new_n880), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(G330), .ZN(new_n914));
  INV_X1    g0714(.A(new_n878), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n877), .B1(new_n472), .B2(new_n475), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n324), .A2(new_n716), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT101), .Z(new_n919));
  AOI21_X1  g0719(.A(new_n917), .B1(new_n841), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n901), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n888), .A2(new_n896), .A3(KEYINPUT38), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n922), .B1(new_n923), .B2(new_n908), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n472), .A2(new_n716), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n924), .B(new_n925), .C1(new_n901), .C2(new_n922), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n419), .A2(new_n889), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n921), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n660), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n732), .A2(new_n759), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n481), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n928), .B(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n914), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n257), .B2(new_n763), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n497), .B1(new_n618), .B2(KEYINPUT35), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(new_n229), .C1(KEYINPUT35), .C2(new_n618), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT36), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n233), .A2(new_n393), .A3(G77), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(G50), .B2(new_n409), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(G1), .A3(new_n297), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n934), .A2(new_n937), .A3(new_n940), .ZN(G367));
  OR2_X1    g0741(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n686), .A2(new_n707), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n942), .B(new_n943), .C1(new_n720), .C2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n833), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n761), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n671), .B1(new_n628), .B2(new_n707), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n670), .A2(new_n625), .A3(new_n716), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n723), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT45), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT45), .B1(new_n951), .B2(new_n723), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT44), .B1(new_n951), .B2(new_n723), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n951), .A2(new_n723), .A3(KEYINPUT44), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n721), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n958), .B(new_n957), .C1(new_n954), .C2(new_n955), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(new_n833), .A3(new_n720), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT105), .B1(new_n948), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n959), .A2(new_n961), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT105), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n833), .A2(new_n946), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n833), .A2(new_n946), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n760), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n964), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n760), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n726), .B(KEYINPUT41), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n764), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n951), .A2(new_n722), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT42), .Z(new_n975));
  AOI21_X1  g0775(.A(new_n612), .B1(new_n949), .B2(new_n950), .ZN(new_n976));
  INV_X1    g0776(.A(new_n647), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n707), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n707), .B1(new_n577), .B2(new_n589), .ZN(new_n979));
  MUX2_X1   g0779(.A(new_n680), .B(new_n677), .S(new_n979), .Z(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT103), .Z(new_n981));
  AOI22_X1  g0781(.A1(new_n975), .A2(new_n978), .B1(KEYINPUT43), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n833), .A2(new_n720), .A3(new_n951), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n973), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n981), .A2(new_n829), .ZN(new_n988));
  INV_X1    g0788(.A(new_n769), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n779), .B1(new_n206), .B2(new_n576), .C1(new_n237), .C2(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n784), .A2(G294), .B1(G283), .B2(new_n804), .ZN(new_n991));
  INV_X1    g0791(.A(new_n483), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n791), .C2(new_n825), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n797), .A2(G107), .B1(new_n800), .B2(G311), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n995), .B2(new_n788), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n811), .A2(new_n501), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n793), .A2(new_n497), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT46), .ZN(new_n999));
  NOR4_X1   g0799(.A1(new_n993), .A2(new_n996), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n793), .A2(new_n216), .B1(new_n788), .B2(new_n848), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT106), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n812), .A2(G77), .B1(G143), .B2(new_n800), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n796), .A2(new_n409), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n277), .B(new_n1004), .C1(G150), .C2(new_n802), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1002), .B(new_n1006), .C1(G159), .C2(new_n784), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n804), .A2(G50), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1000), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n778), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n766), .B(new_n990), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n988), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n987), .A2(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(new_n726), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n966), .A2(new_n760), .A3(new_n967), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT109), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1019), .B(new_n948), .C1(new_n1018), .C2(new_n1017), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n947), .A2(new_n765), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n784), .A2(G311), .B1(new_n800), .B2(G322), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n791), .B2(new_n803), .C1(new_n995), .C2(new_n825), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT48), .ZN(new_n1024));
  INV_X1    g0824(.A(G283), .ZN(new_n1025));
  INV_X1    g0825(.A(G294), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1024), .B1(new_n1025), .B2(new_n796), .C1(new_n1026), .C2(new_n793), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT49), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n483), .B1(new_n789), .B2(G326), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n811), .B2(new_n497), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n576), .A2(new_n796), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n825), .A2(new_n210), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1032), .B(new_n997), .C1(new_n354), .C2(new_n784), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n483), .B1(new_n803), .B2(new_n409), .C1(new_n815), .C2(new_n799), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G77), .B2(new_n819), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1033), .B(new_n1035), .C1(new_n849), .C2(new_n788), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1028), .A2(new_n1030), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n778), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n572), .A2(G116), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n771), .C1(new_n409), .C2(new_n212), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT107), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n292), .A2(new_n210), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT50), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n769), .B1(new_n1041), .B2(new_n1043), .C1(new_n241), .C2(new_n771), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n206), .A2(new_n333), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1044), .B1(G107), .B2(new_n206), .C1(new_n1039), .C2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n767), .B1(new_n1046), .B2(new_n779), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT108), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1038), .B(new_n1048), .C1(new_n720), .C2(new_n829), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1020), .A2(new_n1021), .A3(new_n1049), .ZN(G393));
  NAND2_X1  g0850(.A1(new_n964), .A2(new_n765), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n951), .A2(KEYINPUT110), .A3(new_n829), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n779), .B1(new_n501), .B2(new_n206), .C1(new_n248), .C2(new_n989), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT111), .Z(new_n1054));
  AOI211_X1 g0854(.A(new_n992), .B(new_n858), .C1(new_n292), .C2(new_n804), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n819), .A2(new_n219), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n802), .A2(G159), .B1(new_n800), .B2(G150), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT51), .Z(new_n1058));
  AOI22_X1  g0858(.A1(new_n784), .A2(G50), .B1(G143), .B2(new_n789), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n796), .A2(new_n212), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n802), .A2(G311), .B1(new_n800), .B2(G317), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT112), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n277), .B1(new_n1026), .B2(new_n803), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G303), .B2(new_n784), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n819), .A2(G283), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n797), .A2(G116), .B1(G322), .B2(new_n789), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1066), .A2(new_n814), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1060), .A2(new_n1061), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n767), .B(new_n1054), .C1(new_n1070), .C2(new_n778), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT110), .B1(new_n951), .B2(new_n829), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1052), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1016), .B1(new_n963), .B2(new_n969), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT113), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n948), .A2(new_n962), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1051), .B(new_n1073), .C1(new_n1078), .C2(new_n1079), .ZN(G390));
  INV_X1    g0880(.A(KEYINPUT115), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT114), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n653), .A2(new_n524), .A3(new_n707), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n744), .A2(new_n734), .A3(new_n716), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1084), .A2(new_n745), .ZN(new_n1085));
  OAI211_X1 g0885(.A(G330), .B(new_n840), .C1(new_n1083), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n917), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n752), .A2(new_n753), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n757), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n716), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n918), .B1(new_n1090), .B2(new_n840), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n750), .A2(new_n879), .A3(new_n840), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1087), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1087), .A2(new_n1092), .B1(new_n841), .B2(new_n919), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n481), .A2(new_n930), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n874), .B1(new_n429), .B2(new_n434), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT78), .B1(new_n1097), .B2(new_n376), .ZN(new_n1098));
  AND4_X1   g0898(.A1(KEYINPUT78), .A2(new_n376), .A3(new_n435), .A4(new_n476), .ZN(new_n1099));
  OAI211_X1 g0899(.A(G330), .B(new_n880), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1096), .A2(new_n1100), .A3(new_n660), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1082), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n841), .A2(new_n919), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1086), .A2(new_n917), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n879), .B1(new_n750), .B2(new_n840), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1087), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1108), .A2(new_n931), .A3(KEYINPUT114), .A4(new_n1100), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1102), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n924), .B1(new_n901), .B2(new_n922), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n920), .B2(new_n925), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n925), .B1(new_n909), .B2(new_n900), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1091), .B2(new_n917), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1112), .A2(new_n1114), .A3(new_n1092), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1092), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1081), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n1104), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1112), .A2(new_n1114), .A3(new_n1092), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1122), .A2(KEYINPUT115), .A3(new_n1102), .A4(new_n1109), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1110), .A2(new_n1117), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1118), .A2(new_n726), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n846), .B1(G97), .B2(new_n804), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n277), .C1(new_n273), .C2(new_n823), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n825), .A2(new_n497), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n799), .A2(new_n1025), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n820), .B1(new_n212), .B2(new_n796), .C1(new_n1026), .C2(new_n788), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n277), .B1(G137), .B2(new_n784), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n793), .A2(new_n849), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .C1(new_n210), .C2(new_n811), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT54), .B(G143), .Z(new_n1137));
  AND2_X1   g0937(.A1(new_n804), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n797), .A2(G159), .B1(G125), .B2(new_n789), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(new_n854), .C2(new_n825), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n800), .A2(G128), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n1136), .A2(new_n1138), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n778), .B1(new_n1131), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1144), .B(new_n766), .C1(new_n354), .C2(new_n867), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1111), .B2(new_n775), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n1117), .B2(new_n765), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1125), .A2(new_n1147), .ZN(G378));
  INV_X1    g0948(.A(new_n1101), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1124), .A2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1151));
  XNOR2_X1  g0951(.A(new_n369), .B(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n706), .A2(new_n356), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n911), .A2(G330), .A3(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n899), .A2(new_n900), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n879), .A2(new_n880), .A3(new_n840), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n903), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n910), .A2(new_n881), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1154), .B1(new_n1161), .B2(new_n733), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n928), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1156), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1156), .B2(new_n1162), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1150), .A2(KEYINPUT57), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1101), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1155), .B1(new_n911), .B2(G330), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1161), .A2(new_n733), .A3(new_n1154), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n928), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1156), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1168), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1167), .A2(new_n726), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1155), .A2(new_n775), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n804), .A2(new_n284), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n823), .B2(new_n501), .C1(new_n811), .C2(new_n216), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1004), .B(new_n1179), .C1(G283), .C2(new_n789), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n992), .B1(new_n825), .B2(new_n273), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G41), .B(new_n1181), .C1(G116), .C2(new_n800), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(new_n212), .C2(new_n793), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT58), .Z(new_n1184));
  OAI21_X1  g0984(.A(new_n210), .B1(new_n265), .B2(G41), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n797), .A2(G150), .B1(new_n819), .B2(new_n1137), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G125), .A2(new_n800), .B1(new_n804), .B2(G137), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n802), .A2(G128), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n784), .A2(G132), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G41), .B1(new_n1190), .B2(KEYINPUT59), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G33), .B1(new_n789), .B2(G124), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(new_n815), .C2(new_n811), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1185), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n778), .B1(new_n1184), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n767), .B1(new_n210), .B2(new_n866), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1177), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1166), .B2(new_n765), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1176), .A2(new_n1200), .ZN(G375));
  NAND2_X1  g1001(.A1(new_n1095), .A2(new_n1101), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1102), .A2(new_n1109), .A3(new_n971), .A4(new_n1202), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT117), .Z(new_n1204));
  XNOR2_X1  g1004(.A(new_n764), .B(KEYINPUT118), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1095), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT119), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n812), .A2(G58), .B1(G150), .B2(new_n804), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n210), .B2(new_n796), .C1(new_n854), .C2(new_n799), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n784), .B2(new_n1137), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n789), .A2(G128), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n819), .A2(G159), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n992), .B1(new_n802), .B2(G137), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n277), .B1(new_n273), .B2(new_n803), .C1(new_n823), .C2(new_n497), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n811), .A2(new_n212), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n825), .A2(new_n1025), .B1(new_n788), .B2(new_n791), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1031), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n501), .B2(new_n793), .C1(new_n1026), .C2(new_n799), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1011), .B1(new_n1215), .B2(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n767), .B(new_n1221), .C1(new_n409), .C2(new_n866), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n774), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n879), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1208), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1204), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(G381));
  INV_X1    g1027(.A(KEYINPUT120), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G378), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1125), .A2(KEYINPUT120), .A3(new_n1147), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G375), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1073), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT113), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1232), .B1(new_n1234), .B2(new_n1077), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1013), .B1(new_n973), .B2(new_n986), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n1051), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1231), .A2(new_n1226), .A3(new_n1238), .ZN(new_n1239));
  OR4_X1    g1039(.A1(G396), .A2(new_n1239), .A3(G384), .A4(G393), .ZN(G407));
  INV_X1    g1040(.A(G343), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(G213), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT121), .Z(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1231), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(G407), .A2(G213), .A3(new_n1245), .ZN(G409));
  AND2_X1   g1046(.A1(new_n1208), .A2(new_n1224), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n1101), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1109), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(new_n1202), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n726), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1247), .A2(new_n1251), .A3(G384), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G384), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1206), .B1(new_n1169), .B2(new_n972), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1199), .B1(new_n1255), .B2(new_n1166), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1176), .A2(G378), .A3(new_n1200), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1242), .B(new_n1254), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(G384), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1250), .A2(new_n726), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n1225), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1247), .A2(new_n1251), .A3(G384), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1264), .A2(KEYINPUT62), .A3(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1243), .B(new_n1266), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT125), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1125), .A2(KEYINPUT120), .A3(new_n1147), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT120), .B1(new_n1125), .B2(new_n1147), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1255), .A2(new_n1166), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1270), .A2(new_n1271), .B1(new_n1272), .B2(new_n1199), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1176), .A2(G378), .A3(new_n1200), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1275), .A2(KEYINPUT125), .A3(new_n1243), .A4(new_n1266), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1261), .A2(new_n1269), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1243), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1243), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1241), .A2(G213), .A3(G2897), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1279), .A2(G2897), .B1(new_n1254), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1277), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  XOR2_X1   g1085(.A(G393), .B(G396), .Z(new_n1286));
  INV_X1    g1086(.A(KEYINPUT122), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(G390), .B2(G387), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1236), .B1(new_n1235), .B2(new_n1051), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1286), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1286), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G390), .A2(G387), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1237), .A4(new_n1287), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1277), .A2(KEYINPUT126), .A3(new_n1282), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1285), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1297), .B(new_n1244), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1254), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n1290), .A3(new_n1293), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1242), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1297), .B1(new_n1302), .B2(new_n1281), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1259), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1301), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT123), .B1(new_n1300), .B2(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1302), .A2(new_n1281), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1259), .B1(new_n1307), .B2(new_n1297), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1294), .B1(new_n1254), .B2(new_n1298), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT123), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .A4(new_n1301), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1306), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1296), .A2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(new_n1254), .A2(KEYINPUT127), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1294), .B(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1258), .B1(G375), .B2(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1315), .B(new_n1317), .ZN(G402));
endmodule


