//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT76), .B(G107), .ZN(new_n189));
  OR3_X1    g003(.A1(new_n189), .A2(KEYINPUT80), .A3(G104), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G104), .ZN(new_n192));
  OAI211_X1 g006(.A(KEYINPUT80), .B(new_n192), .C1(new_n189), .C2(G104), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(G101), .A3(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  OAI21_X1  g013(.A(G128), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT81), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n195), .A2(new_n199), .A3(G128), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT81), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n196), .A2(new_n200), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT3), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n191), .A2(KEYINPUT76), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT76), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT77), .B1(new_n192), .B2(KEYINPUT3), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n189), .A2(KEYINPUT77), .A3(new_n209), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT78), .A2(G101), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT78), .A2(G101), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n218), .B(new_n219), .C1(G104), .C2(new_n191), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n207), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  AOI211_X1 g036(.A(KEYINPUT79), .B(new_n220), .C1(new_n215), .C2(new_n216), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n194), .B(new_n206), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT10), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT64), .B1(new_n197), .B2(G146), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n197), .A2(G146), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n232), .A2(new_n235), .B1(new_n195), .B2(new_n233), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G101), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n191), .A2(G104), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n238), .B1(new_n217), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n237), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n222), .A2(new_n223), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n239), .B1(new_n215), .B2(new_n216), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT4), .B1(new_n245), .B2(new_n238), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n243), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G137), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(G137), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT11), .A3(G134), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G131), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n250), .A2(new_n253), .A3(new_n256), .A4(new_n251), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n232), .A2(new_n200), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n225), .B1(new_n260), .B2(new_n203), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n261), .B(new_n194), .C1(new_n222), .C2(new_n223), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n226), .A2(new_n247), .A3(new_n259), .A4(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G110), .B(G140), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n265), .A2(G227), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n264), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n194), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n217), .A2(new_n221), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT79), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n217), .A2(new_n207), .A3(new_n221), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n260), .A2(new_n203), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n224), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT12), .A3(new_n258), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n258), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n269), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n226), .A2(new_n247), .A3(new_n262), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n258), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n268), .B1(new_n283), .B2(new_n263), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n187), .B(new_n188), .C1(new_n281), .C2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n268), .A3(new_n263), .ZN(new_n286));
  INV_X1    g100(.A(new_n263), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n280), .B2(new_n277), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n286), .B(G469), .C1(new_n288), .C2(new_n268), .ZN(new_n289));
  NAND2_X1  g103(.A1(G469), .A2(G902), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT9), .B(G234), .ZN(new_n292));
  OAI21_X1  g106(.A(G221), .B1(new_n292), .B2(G902), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n293), .B(KEYINPUT75), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT82), .ZN(new_n297));
  OAI21_X1  g111(.A(G214), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n300), .B(KEYINPUT86), .Z(new_n301));
  XNOR2_X1  g115(.A(G110), .B(G122), .ZN(new_n302));
  XNOR2_X1  g116(.A(G116), .B(G119), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT2), .B(G113), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n305), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n303), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(new_n241), .B2(new_n242), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(new_n244), .B2(new_n246), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n303), .A2(KEYINPUT5), .ZN(new_n313));
  INV_X1    g127(.A(G116), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n314), .A2(KEYINPUT5), .A3(G119), .ZN(new_n315));
  INV_X1    g129(.A(G113), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n313), .A2(new_n317), .B1(new_n307), .B2(new_n303), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n194), .B(new_n318), .C1(new_n222), .C2(new_n223), .ZN(new_n319));
  AOI211_X1 g133(.A(KEYINPUT6), .B(new_n302), .C1(new_n312), .C2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n275), .A2(G125), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT84), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n236), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n321), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT84), .B1(new_n236), .B2(new_n323), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n265), .A2(G224), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n312), .A2(new_n319), .A3(new_n302), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT83), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n312), .A2(KEYINPUT83), .A3(new_n319), .A4(new_n302), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n302), .B1(new_n312), .B2(new_n319), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT6), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI211_X1 g151(.A(new_n320), .B(new_n329), .C1(new_n334), .C2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT7), .ZN(new_n339));
  INV_X1    g153(.A(new_n328), .ZN(new_n340));
  OAI22_X1  g154(.A1(new_n321), .A2(new_n324), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n340), .B2(KEYINPUT85), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(KEYINPUT85), .B2(new_n340), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n341), .B1(new_n327), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n274), .B(new_n318), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n302), .B(KEYINPUT8), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n334), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n188), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n301), .B1(new_n338), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n334), .A2(new_n337), .ZN(new_n351));
  INV_X1    g165(.A(new_n320), .ZN(new_n352));
  INV_X1    g166(.A(new_n329), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(G902), .B1(new_n334), .B2(new_n347), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n300), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n299), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G140), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n323), .B2(KEYINPUT72), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT72), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(G125), .A3(G140), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(KEYINPUT16), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT16), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n323), .B2(G140), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G146), .ZN(new_n366));
  XNOR2_X1  g180(.A(G125), .B(G140), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT19), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n359), .A2(KEYINPUT19), .A3(new_n361), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n229), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G237), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n265), .A3(G214), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT87), .A3(new_n197), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n197), .A2(KEYINPUT87), .ZN(new_n375));
  NOR2_X1   g189(.A1(G237), .A2(G953), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(G214), .A3(new_n376), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n374), .A2(new_n256), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n256), .B1(new_n374), .B2(new_n377), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n366), .B(new_n371), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n374), .A2(new_n377), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT18), .A3(G131), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n367), .A2(new_n229), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n359), .A2(G146), .A3(new_n361), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT18), .A2(G131), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n374), .A2(new_n386), .A3(new_n377), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n380), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(G113), .B(G122), .Z(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n208), .ZN(new_n391));
  XNOR2_X1  g205(.A(G113), .B(G122), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n391), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n396), .B1(new_n391), .B2(new_n393), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n362), .A2(new_n229), .A3(new_n364), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n401), .A3(new_n366), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT17), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n399), .B(new_n388), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT89), .ZN(new_n406));
  NOR2_X1   g220(.A1(G475), .A2(G902), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n395), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT20), .ZN(new_n411));
  NOR3_X1   g225(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n388), .B1(new_n402), .B2(new_n403), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n394), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n404), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n188), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n419), .A2(G475), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n414), .A2(new_n415), .A3(new_n421), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n410), .A2(KEYINPUT20), .B1(new_n405), .B2(new_n412), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT90), .B1(new_n423), .B2(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT92), .ZN(new_n426));
  INV_X1    g240(.A(G122), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G116), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT91), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n314), .A2(G122), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT14), .ZN(new_n432));
  OAI21_X1  g246(.A(G107), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n189), .A3(new_n431), .ZN(new_n434));
  XNOR2_X1  g248(.A(G128), .B(G143), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(new_n249), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G128), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT13), .B1(new_n438), .B2(G143), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(new_n249), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(new_n435), .ZN(new_n441));
  INV_X1    g255(.A(new_n434), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n189), .B1(new_n429), .B2(new_n431), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n437), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G217), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n292), .A2(new_n446), .A3(G953), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n437), .A2(new_n444), .A3(new_n447), .ZN(new_n450));
  AOI21_X1  g264(.A(G902), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G478), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT15), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n451), .A2(new_n454), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n426), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n451), .A2(new_n454), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT92), .A3(new_n455), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT93), .B(G952), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(G953), .ZN(new_n463));
  NAND2_X1  g277(.A1(G234), .A2(G237), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT21), .B(G898), .Z(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT94), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(G902), .A3(G953), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n425), .A2(new_n461), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n291), .A2(new_n472), .A3(new_n295), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n297), .A2(new_n357), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n252), .A2(G134), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n249), .A2(G137), .ZN(new_n476));
  OAI21_X1  g290(.A(G131), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n257), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n275), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n258), .A2(new_n236), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n309), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n480), .A3(new_n310), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT28), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n376), .A2(G210), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT27), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT26), .B(G101), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n479), .A2(new_n480), .A3(new_n310), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n490), .A2(KEYINPUT28), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n485), .A2(KEYINPUT29), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n188), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT67), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(KEYINPUT67), .A3(new_n188), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT66), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n310), .B1(new_n479), .B2(new_n480), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n498), .B(KEYINPUT28), .C1(new_n490), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n491), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n498), .B1(new_n484), .B2(KEYINPUT28), .ZN(new_n502));
  INV_X1    g316(.A(new_n489), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n479), .A2(new_n480), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n479), .B2(new_n480), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n309), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n483), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n503), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT29), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G472), .B1(new_n497), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n489), .A3(new_n483), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT31), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT65), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n503), .B1(new_n501), .B2(new_n502), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n508), .A2(new_n520), .A3(new_n489), .A4(new_n483), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n515), .A2(KEYINPUT65), .A3(KEYINPUT31), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n518), .A2(new_n519), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT32), .ZN(new_n524));
  NOR2_X1   g338(.A1(G472), .A2(G902), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n514), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT68), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT68), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n514), .B(new_n530), .C1(new_n526), .C2(new_n527), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n446), .B1(G234), .B2(new_n188), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT22), .B(G137), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n265), .A2(G221), .A3(G234), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT23), .ZN(new_n537));
  INV_X1    g351(.A(G119), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n537), .B1(new_n538), .B2(G128), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(G128), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n438), .A2(KEYINPUT23), .A3(G119), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G110), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n362), .A2(new_n229), .A3(new_n364), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n229), .B1(new_n362), .B2(new_n364), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n438), .A2(G119), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n540), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT69), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT24), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(G110), .ZN(new_n551));
  INV_X1    g365(.A(G110), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT24), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT70), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT69), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n547), .A2(new_n540), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(KEYINPUT24), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n550), .A2(G110), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT70), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n549), .A2(new_n554), .A3(new_n556), .A4(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n549), .A2(new_n556), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n554), .A2(new_n560), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT71), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n546), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n366), .A2(new_n383), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n549), .A2(new_n556), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n554), .A2(new_n560), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n542), .A2(G110), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n569), .A2(new_n570), .B1(new_n571), .B2(KEYINPUT73), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n542), .B2(G110), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n568), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n567), .A2(new_n575), .A3(KEYINPUT74), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT74), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n366), .A2(new_n401), .B1(G110), .B2(new_n542), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT71), .B1(new_n564), .B2(new_n565), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n561), .A2(new_n562), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n569), .A2(new_n570), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n571), .A2(KEYINPUT73), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n574), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n545), .B1(new_n229), .B2(new_n367), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n577), .B1(new_n581), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n536), .B1(new_n576), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n536), .B1(new_n581), .B2(new_n586), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT25), .B1(new_n591), .B2(new_n188), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT25), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n593), .B(G902), .C1(new_n588), .C2(new_n590), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n532), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT74), .B1(new_n567), .B2(new_n575), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n581), .A2(new_n577), .A3(new_n586), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n589), .B1(new_n598), .B2(new_n536), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n532), .A2(G902), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n595), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n529), .A2(new_n531), .A3(new_n603), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n474), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n218), .A2(new_n219), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G3));
  NAND2_X1  g421(.A1(new_n523), .A2(new_n188), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G472), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n523), .A2(new_n525), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND4_X1   g425(.A1(new_n603), .A2(new_n297), .A3(new_n473), .A4(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT95), .Z(new_n613));
  INV_X1    g427(.A(new_n300), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n338), .B2(new_n349), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n299), .B1(new_n615), .B2(new_n356), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n469), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT97), .B(G478), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n451), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n449), .A2(new_n450), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n450), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n620), .B(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n452), .A2(G902), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n619), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n422), .B2(new_n424), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n617), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n613), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT98), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  AND3_X1   g447(.A1(new_n410), .A2(KEYINPUT99), .A3(KEYINPUT20), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT99), .B1(new_n410), .B2(KEYINPUT20), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT20), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n406), .A2(new_n637), .A3(new_n407), .A4(new_n409), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT100), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n640));
  OR3_X1    g454(.A1(new_n636), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n640), .B1(new_n636), .B2(new_n639), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n641), .A2(new_n642), .A3(new_n421), .A4(new_n461), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n617), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n613), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  NAND3_X1  g461(.A1(new_n297), .A2(new_n473), .A3(new_n611), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n649));
  INV_X1    g463(.A(new_n532), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n593), .B1(new_n599), .B2(G902), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n591), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n536), .A2(KEYINPUT36), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n576), .A2(new_n587), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n654), .B1(new_n596), .B2(new_n597), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n600), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n655), .B1(new_n576), .B2(new_n587), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n596), .A2(new_n597), .A3(new_n654), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(KEYINPUT102), .A3(new_n600), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n649), .B1(new_n653), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT102), .B1(new_n663), .B2(new_n600), .ZN(new_n667));
  AOI211_X1 g481(.A(new_n659), .B(new_n601), .C1(new_n661), .C2(new_n662), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n595), .A2(KEYINPUT103), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n357), .A3(new_n471), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n648), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT37), .B(G110), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  AND3_X1   g489(.A1(new_n529), .A2(new_n531), .A3(new_n671), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n465), .B1(G900), .B2(new_n468), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n643), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n473), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n472), .B1(new_n291), .B2(new_n295), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n676), .A2(new_n679), .A3(new_n682), .A4(new_n616), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  NAND2_X1  g498(.A1(new_n297), .A2(new_n473), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n677), .B(KEYINPUT39), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  OR3_X1    g501(.A1(new_n685), .A2(KEYINPUT40), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n350), .A2(new_n356), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n689), .B(KEYINPUT38), .Z(new_n690));
  AOI21_X1  g504(.A(new_n299), .B1(new_n458), .B2(new_n460), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n425), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT40), .B1(new_n685), .B2(new_n687), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n610), .A2(KEYINPUT32), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n509), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n503), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n188), .B1(new_n484), .B2(new_n489), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n653), .A2(new_n665), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n688), .A2(new_n693), .A3(new_n694), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  NAND2_X1  g520(.A1(new_n627), .A2(new_n677), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n676), .A2(new_n682), .A3(new_n616), .A4(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n529), .A2(new_n671), .A3(new_n531), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n685), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(KEYINPUT104), .A3(new_n616), .A4(new_n708), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  AND3_X1   g530(.A1(new_n529), .A2(new_n531), .A3(new_n603), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n188), .B1(new_n281), .B2(new_n284), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G469), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n295), .A3(new_n285), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n717), .A2(new_n629), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND3_X1  g538(.A1(new_n717), .A2(new_n644), .A3(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND3_X1  g540(.A1(new_n721), .A2(new_n616), .A3(new_n471), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n676), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT105), .B1(new_n712), .B2(new_n727), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  AOI21_X1  g547(.A(new_n692), .B1(new_n356), .B2(new_n615), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n485), .A2(new_n491), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n521), .B1(new_n735), .B2(new_n489), .ZN(new_n736));
  INV_X1    g550(.A(new_n516), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n525), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n609), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n602), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n720), .A2(new_n470), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n734), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NOR2_X1   g557(.A1(new_n739), .A2(new_n703), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n708), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n721), .A2(new_n616), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  NAND3_X1  g562(.A1(new_n350), .A2(new_n298), .A3(new_n356), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n296), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n529), .A3(new_n531), .A4(new_n603), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n528), .A2(new_n603), .A3(new_n627), .A4(new_n677), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n750), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n752), .A2(new_n753), .B1(KEYINPUT42), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n642), .A2(new_n421), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n461), .A3(new_n641), .A4(new_n677), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n758), .B1(new_n751), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n717), .A2(new_n679), .A3(KEYINPUT106), .A4(new_n750), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  INV_X1    g578(.A(new_n425), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT109), .ZN(new_n766));
  INV_X1    g580(.A(new_n626), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n425), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(KEYINPUT43), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n425), .B2(new_n626), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n611), .A2(new_n703), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(KEYINPUT112), .A3(KEYINPUT44), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n773), .A2(new_n774), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT110), .B1(new_n770), .B2(new_n772), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n778), .B(KEYINPUT44), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n775), .A2(new_n778), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n749), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n286), .B1(new_n288), .B2(new_n268), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n187), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n789), .A2(new_n790), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n290), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT108), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n795), .A2(new_n798), .A3(KEYINPUT46), .A4(new_n290), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT46), .B1(new_n795), .B2(new_n290), .ZN(new_n801));
  INV_X1    g615(.A(new_n285), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n294), .B(new_n687), .C1(new_n800), .C2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n785), .A2(new_n788), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  INV_X1    g620(.A(new_n749), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n708), .A2(new_n807), .A3(new_n602), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n529), .B2(new_n531), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n294), .B1(new_n800), .B2(new_n803), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(KEYINPUT47), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n812), .B(new_n294), .C1(new_n800), .C2(new_n803), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n809), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G140), .ZN(G42));
  INV_X1    g629(.A(new_n702), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n749), .A2(new_n720), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n602), .A2(new_n465), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n425), .A3(new_n767), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n465), .B1(new_n770), .B2(new_n772), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n817), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n820), .B1(new_n822), .B2(new_n744), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n740), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n690), .A2(new_n299), .A3(new_n721), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  OAI211_X1 g643(.A(KEYINPUT51), .B(new_n823), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n811), .A2(new_n813), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n719), .A2(new_n285), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n831), .B1(new_n295), .B2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT116), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n824), .A2(new_n749), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n833), .B2(KEYINPUT116), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n830), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n822), .A2(new_n528), .A3(new_n603), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT48), .Z(new_n840));
  OAI221_X1 g654(.A(new_n463), .B1(new_n628), .B2(new_n819), .C1(new_n824), .C2(new_n746), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n823), .B1(new_n828), .B2(new_n829), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n833), .B2(new_n835), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n842), .B1(new_n844), .B2(KEYINPUT51), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n459), .A2(new_n455), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n678), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n759), .A2(new_n641), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n712), .A2(new_n685), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n745), .A2(new_n296), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n807), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n854), .A2(new_n756), .A3(new_n763), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n717), .B(new_n721), .C1(new_n644), .C2(new_n629), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n648), .A2(new_n672), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n605), .A3(new_n857), .A4(new_n742), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n338), .A2(new_n349), .A3(new_n614), .ZN(new_n859));
  INV_X1    g673(.A(new_n301), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n354), .B2(new_n355), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n298), .B(new_n469), .C1(new_n859), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n765), .A2(new_n849), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT113), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n425), .B1(new_n459), .B2(new_n455), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n357), .A3(new_n866), .A4(new_n469), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n357), .A2(new_n469), .A3(new_n627), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n612), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n729), .B1(new_n676), .B2(new_n728), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n712), .A2(new_n727), .A3(KEYINPUT105), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n858), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n855), .A2(new_n874), .A3(KEYINPUT114), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n854), .A2(new_n763), .A3(new_n756), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n742), .B1(new_n474), .B2(new_n604), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n673), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n732), .A3(new_n856), .A4(new_n870), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n876), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n296), .A2(new_n678), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n704), .A2(new_n734), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT115), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n683), .A2(new_n747), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n715), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT52), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n711), .B2(new_n714), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n891), .A3(new_n885), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n848), .B1(new_n882), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n891), .B1(new_n890), .B2(new_n885), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n891), .A2(new_n715), .A3(new_n887), .A4(new_n885), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n875), .A2(new_n881), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n848), .B1(new_n887), .B2(new_n891), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n847), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT53), .B1(new_n897), .B2(new_n898), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n877), .A2(new_n880), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n848), .B1(new_n886), .B2(KEYINPUT52), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n892), .A2(new_n889), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n902), .A2(KEYINPUT54), .A3(new_n905), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  OAI22_X1  g721(.A1(new_n846), .A2(new_n907), .B1(G952), .B2(G953), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n603), .A2(new_n298), .A3(new_n295), .A4(new_n767), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n832), .A2(KEYINPUT49), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n832), .A2(KEYINPUT49), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n766), .A2(new_n769), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n690), .A3(new_n816), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n908), .A2(new_n914), .ZN(G75));
  NOR2_X1   g729(.A1(new_n265), .A2(G952), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT119), .Z(new_n917));
  INV_X1    g731(.A(new_n905), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n188), .B1(new_n894), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n320), .B1(new_n334), .B2(new_n337), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n353), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n338), .ZN(new_n923));
  XOR2_X1   g737(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n917), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(G902), .B1(new_n902), .B2(new_n905), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT118), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT118), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n930), .B(G902), .C1(new_n902), .C2(new_n905), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n301), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n925), .A2(KEYINPUT56), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(G51));
  XOR2_X1   g748(.A(new_n795), .B(KEYINPUT120), .Z(new_n935));
  NAND3_X1  g749(.A1(new_n929), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n290), .B(KEYINPUT57), .Z(new_n937));
  AOI21_X1  g751(.A(new_n847), .B1(new_n894), .B2(new_n918), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n906), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n281), .A2(new_n284), .ZN(new_n940));
  AOI22_X1  g754(.A1(new_n936), .A2(KEYINPUT121), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n929), .A2(new_n942), .A3(new_n931), .A4(new_n935), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n916), .B1(new_n941), .B2(new_n943), .ZN(G54));
  AND2_X1   g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n929), .A2(new_n931), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n406), .A2(new_n409), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n916), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n947), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n929), .A2(new_n949), .A3(new_n931), .A4(new_n945), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(G60));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT59), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n624), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n894), .A2(new_n847), .A3(new_n918), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT54), .B1(new_n902), .B2(new_n905), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n917), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n952), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n954), .B1(new_n901), .B2(new_n906), .ZN(new_n961));
  INV_X1    g775(.A(new_n624), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n958), .A2(new_n952), .A3(new_n959), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(G63));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT60), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n894), .B2(new_n918), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(new_n591), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n663), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n917), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n970), .A2(KEYINPUT61), .A3(new_n917), .A4(new_n971), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(G66));
  AOI21_X1  g790(.A(new_n265), .B1(new_n467), .B2(G224), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n880), .B2(new_n265), .ZN(new_n978));
  INV_X1    g792(.A(G898), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n921), .B1(new_n979), .B2(G953), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n978), .B(new_n980), .ZN(new_n981));
  XOR2_X1   g795(.A(KEYINPUT123), .B(KEYINPUT124), .Z(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G69));
  OR2_X1    g797(.A1(new_n506), .A2(new_n507), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n369), .A2(new_n370), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n984), .B(new_n985), .Z(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT125), .Z(new_n987));
  AOI21_X1  g801(.A(new_n749), .B1(new_n863), .B2(new_n628), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n717), .A2(new_n682), .A3(new_n686), .A4(new_n988), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n805), .A2(new_n814), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n890), .A2(new_n705), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n987), .B1(new_n994), .B2(G953), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n763), .A2(new_n756), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n890), .A2(new_n996), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n734), .A2(new_n528), .A3(new_n603), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n804), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n805), .A3(new_n814), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(KEYINPUT126), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n999), .A2(new_n1002), .A3(new_n814), .A4(new_n805), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n1001), .A2(new_n265), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(G900), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n986), .B1(new_n1005), .B2(new_n265), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n995), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n265), .B1(G227), .B2(G900), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(G72));
  NAND3_X1  g823(.A1(new_n1001), .A2(new_n874), .A3(new_n1003), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  AOI211_X1 g826(.A(new_n489), .B(new_n509), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n990), .A2(new_n874), .A3(new_n993), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n1012), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n699), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n894), .A2(new_n900), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1012), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(new_n510), .B2(new_n515), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n916), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(KEYINPUT127), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1023), .A2(new_n503), .A3(new_n698), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT127), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1024), .A2(new_n1025), .A3(new_n1016), .A4(new_n1020), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1022), .A2(new_n1026), .ZN(G57));
endmodule


