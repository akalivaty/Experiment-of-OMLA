//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203));
  XOR2_X1   g002(.A(G1gat), .B(G29gat), .Z(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n206), .B(new_n207), .Z(new_n208));
  INV_X1    g007(.A(KEYINPUT5), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  INV_X1    g009(.A(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT2), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n214), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(KEYINPUT71), .A2(KEYINPUT2), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n212), .A2(new_n222), .A3(new_n213), .A4(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT72), .ZN(new_n225));
  XOR2_X1   g024(.A(G155gat), .B(G162gat), .Z(new_n226));
  AND3_X1   g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n225), .B1(new_n224), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n219), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT73), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT73), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n231), .B(new_n219), .C1(new_n227), .C2(new_n228), .ZN(new_n232));
  OR2_X1    g031(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(KEYINPUT65), .A2(G134gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(G127gat), .A3(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(KEYINPUT66), .A2(G127gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT66), .A2(G127gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(G134gat), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240));
  INV_X1    g039(.A(G120gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G113gat), .ZN(new_n242));
  INV_X1    g041(.A(G113gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G120gat), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT1), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  MUX2_X1   g044(.A(new_n239), .B(new_n240), .S(new_n245), .Z(new_n246));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n232), .A3(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n214), .A2(new_n215), .A3(new_n218), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n224), .A2(new_n226), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT72), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n245), .B1(new_n235), .B2(new_n238), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n245), .A2(new_n240), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n247), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n209), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n230), .A2(KEYINPUT3), .A3(new_n232), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n255), .B1(new_n252), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(new_n229), .B2(new_n246), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n255), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n268), .A3(new_n258), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n260), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n264), .A2(new_n268), .A3(new_n209), .A4(new_n258), .ZN(new_n271));
  AOI211_X1 g070(.A(new_n203), .B(new_n208), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  INV_X1    g072(.A(new_n208), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT6), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n270), .A2(new_n208), .A3(new_n271), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G8gat), .B(G36gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT70), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(G190gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT28), .A3(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT27), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(G190gat), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n284), .B1(new_n290), .B2(KEYINPUT28), .ZN(new_n291));
  INV_X1    g090(.A(G169gat), .ZN(new_n292));
  INV_X1    g091(.A(G176gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT26), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n291), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT23), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  AND4_X1   g104(.A1(KEYINPUT25), .A2(new_n303), .A3(new_n305), .A4(new_n296), .ZN(new_n306));
  OR2_X1    g105(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n283), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n298), .A2(KEYINPUT24), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  NOR2_X1   g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n310), .B2(new_n312), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n305), .A3(new_n296), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n322), .A2(new_n323), .B1(G226gat), .B2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G197gat), .B(G204gat), .ZN(new_n326));
  INV_X1    g125(.A(G211gat), .ZN(new_n327));
  INV_X1    g126(.A(G218gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n326), .B1(KEYINPUT22), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n330), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G226gat), .ZN(new_n334));
  INV_X1    g133(.A(G233gat), .ZN(new_n335));
  AOI211_X1 g134(.A(new_n334), .B(new_n335), .C1(new_n302), .C2(new_n321), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n325), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n330), .B(new_n331), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n324), .B2(new_n336), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n281), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n340), .A3(new_n281), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT30), .A4(new_n281), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n202), .B1(new_n277), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT69), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT32), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n282), .A2(KEYINPUT28), .A3(new_n283), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT27), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n307), .B2(new_n308), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n283), .B1(new_n352), .B2(new_n288), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT28), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n321), .B(new_n255), .C1(new_n355), .C2(new_n300), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n302), .A2(KEYINPUT67), .A3(new_n255), .A4(new_n321), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n354), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n300), .B1(new_n360), .B2(new_n284), .ZN(new_n361));
  INV_X1    g160(.A(new_n321), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n246), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n349), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT33), .B1(new_n364), .B2(new_n366), .ZN(new_n368));
  XOR2_X1   g167(.A(G15gat), .B(G43gat), .Z(new_n369));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n367), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  AOI221_X4 g172(.A(new_n349), .B1(KEYINPUT33), .B2(new_n371), .C1(new_n364), .C2(new_n366), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n348), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n358), .A2(new_n363), .A3(new_n365), .A4(new_n359), .ZN(new_n376));
  XOR2_X1   g175(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n381), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n383), .B(new_n348), .C1(new_n373), .C2(new_n374), .ZN(new_n384));
  INV_X1    g183(.A(G22gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n262), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n323), .B1(new_n229), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT78), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(new_n323), .C1(new_n229), .C2(new_n386), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n339), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n339), .A2(KEYINPUT29), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n230), .B(new_n232), .C1(new_n392), .C2(KEYINPUT3), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n391), .A2(G228gat), .A3(G233gat), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n252), .A2(new_n262), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n333), .B1(new_n396), .B2(new_n323), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n333), .A2(new_n323), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n252), .B1(new_n398), .B2(new_n262), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n395), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n385), .B1(new_n394), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n388), .A2(new_n339), .A3(new_n390), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n393), .A2(G228gat), .A3(G233gat), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n400), .B(new_n385), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(G50gat), .ZN(new_n407));
  XOR2_X1   g206(.A(G78gat), .B(G106gat), .Z(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  NAND4_X1  g208(.A1(new_n402), .A2(KEYINPUT79), .A3(new_n405), .A4(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT79), .B1(new_n411), .B2(G22gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n409), .ZN(new_n413));
  INV_X1    g212(.A(new_n405), .ZN(new_n414));
  OAI22_X1  g213(.A1(new_n412), .A2(new_n413), .B1(new_n414), .B2(new_n401), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n382), .A2(new_n384), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n343), .A2(new_n342), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n338), .A2(new_n340), .ZN(new_n418));
  INV_X1    g217(.A(new_n281), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n417), .A2(new_n345), .A3(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n270), .A2(new_n208), .A3(new_n271), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n208), .B1(new_n270), .B2(new_n271), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT6), .ZN(new_n424));
  OAI211_X1 g223(.A(KEYINPUT76), .B(new_n421), .C1(new_n424), .C2(new_n272), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n347), .A2(new_n416), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT86), .B1(new_n426), .B2(KEYINPUT35), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n272), .B(KEYINPUT85), .ZN(new_n428));
  NOR4_X1   g227(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT82), .A4(KEYINPUT6), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n275), .B2(new_n276), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n428), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n410), .A2(new_n415), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n383), .B1(new_n373), .B2(new_n374), .ZN(new_n434));
  OR3_X1    g233(.A1(new_n367), .A2(new_n368), .A3(new_n372), .ZN(new_n435));
  INV_X1    g234(.A(new_n374), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n381), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT80), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n346), .A2(new_n440), .ZN(new_n441));
  AND4_X1   g240(.A1(KEYINPUT80), .A2(new_n417), .A3(new_n345), .A4(new_n420), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT35), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n432), .A2(new_n439), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n427), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n426), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n347), .A2(new_n425), .ZN(new_n448));
  INV_X1    g247(.A(new_n433), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OR2_X1    g249(.A1(new_n438), .A2(KEYINPUT36), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n382), .A2(new_n384), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT36), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT80), .B1(new_n344), .B2(new_n345), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(new_n442), .ZN(new_n457));
  INV_X1    g256(.A(new_n423), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n264), .A2(new_n268), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n259), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT81), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(KEYINPUT81), .A3(new_n259), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT39), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n247), .A2(new_n258), .A3(new_n256), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n462), .A2(KEYINPUT39), .A3(new_n463), .A4(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n208), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n466), .A2(KEYINPUT40), .A3(new_n208), .A4(new_n468), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n457), .A2(new_n458), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT83), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n474), .A2(KEYINPUT37), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n281), .B1(new_n474), .B2(KEYINPUT37), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT84), .B1(new_n477), .B2(KEYINPUT38), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(new_n476), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n477), .A2(KEYINPUT38), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n478), .A2(new_n481), .A3(new_n343), .A4(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n473), .B(new_n433), .C1(new_n432), .C2(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n446), .A2(new_n447), .B1(new_n455), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT15), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT14), .B(G29gat), .ZN(new_n487));
  INV_X1    g286(.A(G36gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G29gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(G43gat), .B(G50gat), .Z(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT88), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n489), .A2(new_n493), .A3(new_n491), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n486), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n486), .B2(new_n495), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n501), .A2(G1gat), .ZN(new_n502));
  AOI21_X1  g301(.A(G8gat), .B1(new_n502), .B2(KEYINPUT89), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT16), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n501), .B1(new_n504), .B2(G1gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n503), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n509), .A2(KEYINPUT90), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n509), .A2(KEYINPUT90), .B1(new_n508), .B2(new_n498), .ZN(new_n511));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n508), .B(new_n498), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n512), .B(KEYINPUT13), .Z(new_n516));
  AOI22_X1  g315(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G197gat), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT11), .B(G169gat), .Z(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n521), .B(new_n522), .Z(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT18), .A4(new_n512), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n517), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n517), .B2(new_n525), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n485), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(KEYINPUT97), .B(G92gat), .Z(new_n530));
  INV_X1    g329(.A(G85gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n530), .A2(new_n531), .B1(KEYINPUT8), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT98), .ZN(new_n534));
  NAND2_X1  g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G99gat), .B(G106gat), .Z(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n537), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n498), .ZN(new_n541));
  NAND3_X1  g340(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n541), .B(new_n542), .C1(new_n500), .C2(new_n540), .ZN(new_n543));
  XOR2_X1   g342(.A(G190gat), .B(G218gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT99), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT100), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n543), .A2(new_n545), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT96), .ZN(new_n551));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  OR4_X1    g352(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n553), .ZN(new_n554));
  OAI22_X1  g353(.A1(new_n548), .A2(new_n553), .B1(new_n547), .B2(new_n549), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G71gat), .B(G78gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT91), .Z(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT92), .Z(new_n560));
  AOI21_X1  g359(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT93), .Z(new_n562));
  OAI21_X1  g361(.A(new_n558), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n557), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G127gat), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n507), .B1(new_n567), .B2(new_n568), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT95), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT94), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G155gat), .ZN(new_n578));
  XOR2_X1   g377(.A(G183gat), .B(G211gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n575), .A2(new_n580), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n556), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G230gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(new_n335), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n537), .B(new_n538), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT101), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n567), .B1(new_n588), .B2(new_n538), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n540), .A2(new_n589), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n540), .A2(KEYINPUT10), .A3(new_n563), .A4(new_n566), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n586), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n592), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n586), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  OR2_X1    g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n596), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n586), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n584), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n529), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n277), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(G1gat), .Z(G1324gat));
  INV_X1    g410(.A(new_n457), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT16), .B(G8gat), .Z(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(KEYINPUT42), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT103), .ZN(new_n616));
  INV_X1    g415(.A(G8gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n613), .B(KEYINPUT102), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n618), .A2(new_n614), .ZN(new_n619));
  OAI221_X1 g418(.A(new_n616), .B1(new_n617), .B2(new_n618), .C1(new_n619), .C2(KEYINPUT42), .ZN(G1325gat));
  AND2_X1   g419(.A1(new_n451), .A2(new_n453), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT104), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(G15gat), .B1(new_n608), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G15gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n438), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n624), .B1(new_n608), .B2(new_n626), .ZN(G1326gat));
  NOR2_X1   g426(.A1(new_n608), .A2(new_n433), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT43), .B(G22gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1327gat));
  AND3_X1   g429(.A1(new_n426), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n631), .A2(new_n427), .A3(new_n445), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n484), .A2(new_n454), .A3(new_n450), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT106), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n427), .ZN(new_n635));
  INV_X1    g434(.A(new_n445), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n447), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n455), .A2(new_n484), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT106), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n556), .A2(KEYINPUT44), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n634), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT44), .B1(new_n485), .B2(new_n556), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT105), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(new_n526), .B2(new_n527), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n517), .A2(new_n525), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n523), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n517), .A2(new_n524), .A3(new_n525), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(KEYINPUT105), .A3(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n583), .A2(new_n606), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n644), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT107), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n644), .A2(KEYINPUT107), .A3(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(G29gat), .B1(new_n659), .B2(new_n609), .ZN(new_n660));
  INV_X1    g459(.A(new_n556), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n529), .A2(new_n661), .A3(new_n652), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(new_n490), .A3(new_n277), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT45), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(G1328gat));
  OAI21_X1  g464(.A(G36gat), .B1(new_n659), .B2(new_n612), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n662), .A2(new_n488), .A3(new_n457), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(KEYINPUT108), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n668), .A2(KEYINPUT108), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n666), .B(new_n671), .C1(new_n669), .C2(new_n667), .ZN(G1329gat));
  INV_X1    g471(.A(G43gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n662), .A2(new_n673), .A3(new_n438), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT47), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n657), .A2(new_n622), .A3(new_n658), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(G43gat), .ZN(new_n678));
  OAI21_X1  g477(.A(G43gat), .B1(new_n655), .B2(new_n454), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n679), .B2(new_n674), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n678), .A2(KEYINPUT109), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n682));
  INV_X1    g481(.A(new_n676), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT107), .B1(new_n644), .B2(new_n654), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n656), .B(new_n653), .C1(new_n642), .C2(new_n643), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n684), .A2(new_n685), .A3(new_n623), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n683), .B1(new_n686), .B2(new_n673), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n679), .A2(new_n674), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT47), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n682), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n681), .A2(new_n690), .ZN(G1330gat));
  OAI21_X1  g490(.A(G50gat), .B1(new_n655), .B2(new_n433), .ZN(new_n692));
  INV_X1    g491(.A(G50gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n662), .A2(new_n693), .A3(new_n449), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(KEYINPUT48), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n694), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n657), .A2(new_n449), .A3(new_n658), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(G50gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n695), .B1(new_n698), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g498(.A1(new_n651), .A2(new_n584), .ZN(new_n700));
  AND4_X1   g499(.A1(new_n606), .A2(new_n634), .A3(new_n640), .A4(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(KEYINPUT110), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(KEYINPUT110), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n277), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g506(.A1(new_n704), .A2(new_n612), .ZN(new_n708));
  NOR2_X1   g507(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n709));
  AND2_X1   g508(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n708), .B2(new_n709), .ZN(G1333gat));
  OAI21_X1  g511(.A(G71gat), .B1(new_n704), .B2(new_n623), .ZN(new_n713));
  INV_X1    g512(.A(G71gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n438), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n704), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT50), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n713), .B(KEYINPUT50), .C1(new_n704), .C2(new_n715), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(G1334gat));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n449), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g521(.A1(new_n651), .A2(new_n583), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n644), .A2(new_n606), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(G85gat), .B1(new_n724), .B2(new_n609), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n723), .B(new_n661), .C1(new_n633), .C2(new_n632), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n730), .B2(new_n729), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n606), .A2(new_n531), .A3(new_n277), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n725), .B1(new_n732), .B2(new_n733), .ZN(G1336gat));
  INV_X1    g533(.A(new_n530), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n724), .B2(new_n612), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737));
  INV_X1    g536(.A(new_n606), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n738), .A2(G92gat), .A3(new_n612), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n736), .B(new_n737), .C1(new_n732), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n726), .A2(KEYINPUT112), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(new_n727), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n736), .B1(new_n742), .B2(new_n739), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT52), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n744), .ZN(G1337gat));
  OAI21_X1  g544(.A(G99gat), .B1(new_n724), .B2(new_n623), .ZN(new_n746));
  INV_X1    g545(.A(G99gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n606), .A2(new_n747), .A3(new_n438), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n732), .B2(new_n748), .ZN(G1338gat));
  OAI21_X1  g548(.A(G106gat), .B1(new_n724), .B2(new_n433), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n738), .A2(G106gat), .A3(new_n433), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n750), .B(new_n751), .C1(new_n732), .C2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n750), .B1(new_n742), .B2(new_n752), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT53), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1339gat));
  INV_X1    g555(.A(new_n583), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n594), .A2(new_n586), .A3(new_n595), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n603), .A2(KEYINPUT54), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n601), .B1(new_n596), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(KEYINPUT55), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n605), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT55), .B1(new_n760), .B2(new_n762), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n758), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n760), .A2(new_n762), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n769), .A2(KEYINPUT113), .A3(new_n605), .A4(new_n763), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n646), .A2(new_n650), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n512), .B1(new_n510), .B2(new_n511), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n515), .A2(new_n516), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n521), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n606), .A2(new_n649), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n661), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n649), .A2(new_n774), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n556), .A2(new_n777), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n778), .A2(new_n766), .A3(new_n770), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n757), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n651), .A2(new_n584), .A3(new_n606), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n457), .A2(new_n609), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n439), .A3(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n785), .A2(new_n243), .A3(new_n528), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n609), .B1(new_n780), .B2(new_n782), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n787), .A2(new_n612), .A3(new_n416), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n651), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n786), .B1(new_n789), .B2(new_n243), .ZN(G1340gat));
  NOR3_X1   g589(.A1(new_n785), .A2(new_n241), .A3(new_n738), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n606), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n241), .ZN(G1341gat));
  NAND4_X1  g592(.A1(new_n788), .A2(new_n236), .A3(new_n237), .A4(new_n583), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n236), .A2(new_n237), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n785), .B2(new_n757), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1342gat));
  NAND4_X1  g596(.A1(new_n788), .A2(new_n233), .A3(new_n234), .A4(new_n661), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n798), .A2(KEYINPUT56), .ZN(new_n799));
  OAI21_X1  g598(.A(G134gat), .B1(new_n785), .B2(new_n556), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n798), .A2(KEYINPUT114), .A3(KEYINPUT56), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT114), .B1(new_n798), .B2(KEYINPUT56), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n799), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(G1343gat));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n769), .A2(new_n605), .A3(new_n763), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n775), .B1(new_n528), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n556), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n778), .A2(new_n766), .A3(new_n770), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(KEYINPUT115), .A3(new_n556), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n781), .B1(new_n812), .B2(new_n757), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT57), .B1(new_n813), .B2(new_n433), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n783), .A2(new_n815), .A3(new_n449), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n454), .A2(new_n784), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n804), .B(G141gat), .C1(new_n819), .C2(new_n528), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n622), .A2(new_n433), .A3(new_n457), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n787), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n528), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n210), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT116), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(KEYINPUT117), .B2(KEYINPUT58), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n651), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n830), .A2(G141gat), .B1(KEYINPUT117), .B2(new_n826), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n828), .B1(new_n831), .B2(new_n804), .ZN(G1344gat));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833));
  OR3_X1    g632(.A1(new_n556), .A2(new_n777), .A3(new_n805), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n583), .B1(new_n807), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n584), .A2(new_n823), .A3(new_n606), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n815), .B(new_n449), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n433), .B1(new_n780), .B2(new_n782), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n606), .B(new_n837), .C1(new_n838), .C2(new_n815), .ZN(new_n839));
  OAI21_X1  g638(.A(G148gat), .B1(new_n839), .B2(new_n817), .ZN(new_n840));
  XOR2_X1   g639(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n814), .A2(new_n606), .A3(new_n816), .A4(new_n818), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n211), .A2(KEYINPUT59), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n840), .A2(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n822), .A2(G148gat), .A3(new_n738), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n833), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n846), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n783), .A2(new_n449), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT57), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n850), .A2(new_n606), .A3(new_n818), .A4(new_n837), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n841), .B1(new_n851), .B2(G148gat), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n843), .A2(new_n844), .ZN(new_n853));
  OAI211_X1 g652(.A(KEYINPUT119), .B(new_n848), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n847), .A2(new_n854), .ZN(G1345gat));
  OAI21_X1  g654(.A(G155gat), .B1(new_n819), .B2(new_n757), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n583), .A2(new_n216), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n822), .B2(new_n857), .ZN(G1346gat));
  NAND3_X1  g657(.A1(new_n829), .A2(G162gat), .A3(new_n661), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n217), .B1(new_n822), .B2(new_n556), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(KEYINPUT120), .A3(new_n860), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1347gat));
  NOR2_X1   g664(.A1(new_n612), .A2(new_n277), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n783), .A2(new_n416), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n292), .A3(new_n651), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT121), .Z(new_n869));
  NAND3_X1  g668(.A1(new_n783), .A2(new_n439), .A3(new_n866), .ZN(new_n870));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870), .B2(new_n528), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT122), .Z(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(G1348gat));
  NAND3_X1  g672(.A1(new_n867), .A2(new_n293), .A3(new_n606), .ZN(new_n874));
  OAI21_X1  g673(.A(G176gat), .B1(new_n870), .B2(new_n738), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1349gat));
  NAND3_X1  g675(.A1(new_n867), .A2(new_n282), .A3(new_n583), .ZN(new_n877));
  OAI22_X1  g676(.A1(new_n870), .A2(new_n757), .B1(new_n286), .B2(new_n285), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n879), .B(new_n880), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n867), .A2(new_n283), .A3(new_n661), .ZN(new_n882));
  OAI21_X1  g681(.A(G190gat), .B1(new_n870), .B2(new_n556), .ZN(new_n883));
  XNOR2_X1  g682(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n883), .A2(new_n885), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(G1351gat));
  NAND2_X1  g687(.A1(new_n623), .A2(new_n866), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n849), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(new_n651), .ZN(new_n891));
  INV_X1    g690(.A(new_n889), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n837), .B(new_n892), .C1(new_n838), .C2(new_n815), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n823), .A2(G197gat), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n891), .A2(G197gat), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(G1352gat));
  XOR2_X1   g695(.A(KEYINPUT125), .B(G204gat), .Z(new_n897));
  NOR2_X1   g696(.A1(new_n738), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n890), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT62), .Z(new_n900));
  OR3_X1    g699(.A1(new_n839), .A2(KEYINPUT126), .A3(new_n889), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT126), .B1(new_n839), .B2(new_n889), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n902), .A3(new_n897), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(G1353gat));
  OAI21_X1  g703(.A(G211gat), .B1(new_n893), .B2(new_n757), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT63), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT63), .B(G211gat), .C1(new_n893), .C2(new_n757), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(KEYINPUT127), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n890), .A2(new_n327), .A3(new_n583), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n909), .B(new_n910), .C1(KEYINPUT127), .C2(new_n907), .ZN(G1354gat));
  OAI21_X1  g710(.A(G218gat), .B1(new_n893), .B2(new_n556), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n890), .A2(new_n328), .A3(new_n661), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1355gat));
endmodule


