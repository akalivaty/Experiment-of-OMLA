

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n663, n665, n666, n667, n668, n670, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774;

  BUF_X1 U373 ( .A(n655), .Z(n359) );
  INV_X1 U374 ( .A(n670), .ZN(n353) );
  INV_X1 U375 ( .A(n663), .ZN(n351) );
  XNOR2_X1 U376 ( .A(n649), .B(n355), .ZN(n653) );
  INV_X1 U377 ( .A(n747), .ZN(n356) );
  INV_X1 U378 ( .A(n747), .ZN(n360) );
  INV_X1 U379 ( .A(n648), .ZN(n355) );
  AND2_X1 U380 ( .A1(n384), .A2(n387), .ZN(n383) );
  NAND2_X1 U381 ( .A1(n382), .A2(n381), .ZN(n380) );
  AND2_X1 U382 ( .A1(n726), .A2(n386), .ZN(n382) );
  NAND2_X1 U383 ( .A1(n400), .A2(n423), .ZN(n379) );
  AND2_X1 U384 ( .A1(n556), .A2(n557), .ZN(n575) );
  NOR2_X1 U385 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U386 ( .A(n363), .B(n374), .ZN(n543) );
  NOR2_X1 U387 ( .A1(n563), .A2(n504), .ZN(n363) );
  NAND2_X1 U388 ( .A1(n600), .A2(n706), .ZN(n590) );
  NAND2_X1 U389 ( .A1(n428), .A2(n425), .ZN(n393) );
  OR2_X1 U390 ( .A1(n666), .A2(n642), .ZN(n459) );
  OR2_X1 U391 ( .A1(n733), .A2(n426), .ZN(n425) );
  XNOR2_X1 U392 ( .A(n521), .B(n520), .ZN(n647) );
  XNOR2_X1 U393 ( .A(n521), .B(n512), .ZN(n733) );
  XOR2_X1 U394 ( .A(KEYINPUT10), .B(n481), .Z(n526) );
  XNOR2_X1 U395 ( .A(n403), .B(n506), .ZN(n402) );
  XNOR2_X1 U396 ( .A(n505), .B(KEYINPUT4), .ZN(n403) );
  XNOR2_X1 U397 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n438) );
  XNOR2_X1 U398 ( .A(G110), .B(G107), .ZN(n445) );
  BUF_X1 U399 ( .A(n492), .Z(n762) );
  INV_X1 U400 ( .A(KEYINPUT71), .ZN(n476) );
  INV_X1 U401 ( .A(G131), .ZN(n475) );
  XNOR2_X1 U402 ( .A(n352), .B(n351), .ZN(G60) );
  XNOR2_X1 U403 ( .A(n354), .B(n353), .ZN(G51) );
  NAND2_X1 U404 ( .A1(n357), .A2(n356), .ZN(n352) );
  NAND2_X1 U405 ( .A1(n361), .A2(n360), .ZN(n354) );
  AND2_X2 U406 ( .A1(n419), .A2(n371), .ZN(n635) );
  AND2_X2 U407 ( .A1(n433), .A2(n641), .ZN(n761) );
  XNOR2_X1 U408 ( .A(n661), .B(n358), .ZN(n357) );
  INV_X1 U409 ( .A(n660), .ZN(n358) );
  XNOR2_X1 U410 ( .A(n668), .B(n362), .ZN(n361) );
  INV_X1 U411 ( .A(n667), .ZN(n362) );
  NOR2_X1 U412 ( .A1(n371), .A2(n683), .ZN(n711) );
  XNOR2_X1 U413 ( .A(n445), .B(G104), .ZN(n754) );
  NOR2_X1 U414 ( .A1(n714), .A2(n563), .ZN(n550) );
  NAND2_X1 U415 ( .A1(n694), .A2(n695), .ZN(n691) );
  XNOR2_X1 U416 ( .A(n616), .B(n401), .ZN(n618) );
  INV_X1 U417 ( .A(G953), .ZN(n492) );
  XOR2_X1 U418 ( .A(KEYINPUT73), .B(G137), .Z(n506) );
  XNOR2_X1 U419 ( .A(KEYINPUT30), .B(KEYINPUT110), .ZN(n594) );
  XNOR2_X1 U420 ( .A(n539), .B(n538), .ZN(n364) );
  NAND2_X1 U421 ( .A1(n592), .A2(n632), .ZN(n687) );
  XNOR2_X1 U422 ( .A(KEYINPUT3), .B(G119), .ZN(n450) );
  XNOR2_X1 U423 ( .A(G101), .B(KEYINPUT75), .ZN(n448) );
  AND2_X1 U424 ( .A1(n618), .A2(n368), .ZN(n405) );
  NAND2_X1 U425 ( .A1(n619), .A2(n411), .ZN(n410) );
  NAND2_X1 U426 ( .A1(n619), .A2(KEYINPUT86), .ZN(n407) );
  NOR2_X1 U427 ( .A1(n620), .A2(KEYINPUT47), .ZN(n621) );
  NAND2_X1 U428 ( .A1(n431), .A2(G902), .ZN(n429) );
  XNOR2_X1 U429 ( .A(n539), .B(n538), .ZN(n587) );
  XNOR2_X1 U430 ( .A(n537), .B(KEYINPUT25), .ZN(n538) );
  XNOR2_X1 U431 ( .A(G128), .B(G137), .ZN(n529) );
  XOR2_X1 U432 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n494) );
  XNOR2_X1 U433 ( .A(n453), .B(n753), .ZN(n666) );
  INV_X1 U434 ( .A(n638), .ZN(n417) );
  BUF_X1 U435 ( .A(n547), .Z(n692) );
  NAND2_X1 U436 ( .A1(n412), .A2(KEYINPUT86), .ZN(n411) );
  INV_X1 U437 ( .A(n617), .ZN(n412) );
  OR2_X1 U438 ( .A1(n619), .A2(n414), .ZN(n409) );
  XNOR2_X1 U439 ( .A(G116), .B(G113), .ZN(n449) );
  XNOR2_X1 U440 ( .A(n687), .B(KEYINPUT92), .ZN(n615) );
  AND2_X1 U441 ( .A1(n367), .A2(n413), .ZN(n628) );
  XNOR2_X1 U442 ( .A(n439), .B(G128), .ZN(n488) );
  INV_X1 U443 ( .A(G143), .ZN(n439) );
  XNOR2_X1 U444 ( .A(n643), .B(KEYINPUT68), .ZN(n644) );
  AND2_X1 U445 ( .A1(n761), .A2(n424), .ZN(n423) );
  NAND2_X1 U446 ( .A1(n500), .A2(KEYINPUT88), .ZN(n424) );
  XNOR2_X1 U447 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n442) );
  AND2_X1 U448 ( .A1(n430), .A2(n429), .ZN(n428) );
  NAND2_X1 U449 ( .A1(n513), .A2(n427), .ZN(n426) );
  XNOR2_X1 U450 ( .A(G116), .B(G107), .ZN(n489) );
  XNOR2_X1 U451 ( .A(n488), .B(n404), .ZN(n507) );
  INV_X1 U452 ( .A(G134), .ZN(n404) );
  INV_X1 U453 ( .A(KEYINPUT65), .ZN(n386) );
  AND2_X1 U454 ( .A1(n599), .A2(n416), .ZN(n603) );
  XNOR2_X1 U455 ( .A(n487), .B(n486), .ZN(n568) );
  XNOR2_X1 U456 ( .A(n485), .B(G475), .ZN(n486) );
  XNOR2_X1 U457 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U458 ( .A(n531), .B(n436), .ZN(n532) );
  XNOR2_X1 U459 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U460 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X1 U461 ( .A1(n568), .A2(n566), .ZN(n617) );
  INV_X1 U462 ( .A(KEYINPUT111), .ZN(n401) );
  AND2_X1 U463 ( .A1(n415), .A2(n599), .ZN(n616) );
  AND2_X1 U464 ( .A1(n598), .A2(n417), .ZN(n415) );
  INV_X1 U465 ( .A(KEYINPUT106), .ZN(n390) );
  NAND2_X1 U466 ( .A1(n543), .A2(n692), .ZN(n571) );
  XOR2_X1 U467 ( .A(n600), .B(n601), .Z(n365) );
  XOR2_X1 U468 ( .A(n466), .B(KEYINPUT97), .Z(n366) );
  AND2_X1 U469 ( .A1(n627), .A2(n626), .ZN(n367) );
  AND2_X1 U470 ( .A1(n617), .A2(n414), .ZN(n368) );
  AND2_X1 U471 ( .A1(n410), .A2(n409), .ZN(n369) );
  AND2_X1 U472 ( .A1(n562), .A2(n364), .ZN(n370) );
  NOR2_X2 U473 ( .A1(n568), .A2(n567), .ZN(n371) );
  AND2_X1 U474 ( .A1(n641), .A2(KEYINPUT2), .ZN(n372) );
  AND2_X1 U475 ( .A1(n692), .A2(n370), .ZN(n373) );
  XOR2_X1 U476 ( .A(KEYINPUT67), .B(KEYINPUT22), .Z(n374) );
  INV_X1 U477 ( .A(KEYINPUT86), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n391), .B(n390), .ZN(n656) );
  INV_X1 U479 ( .A(G902), .ZN(n427) );
  XOR2_X1 U480 ( .A(KEYINPUT35), .B(KEYINPUT90), .Z(n375) );
  INV_X1 U481 ( .A(KEYINPUT88), .ZN(n580) );
  AND2_X1 U482 ( .A1(n644), .A2(KEYINPUT65), .ZN(n376) );
  AND2_X1 U483 ( .A1(n389), .A2(n553), .ZN(n377) );
  NAND2_X1 U484 ( .A1(n642), .A2(n580), .ZN(n378) );
  NAND2_X1 U485 ( .A1(n379), .A2(n376), .ZN(n384) );
  NAND2_X1 U486 ( .A1(n379), .A2(n644), .ZN(n381) );
  NAND2_X2 U487 ( .A1(n383), .A2(n380), .ZN(n739) );
  NAND2_X1 U488 ( .A1(n388), .A2(n748), .ZN(n726) );
  NAND2_X1 U489 ( .A1(n385), .A2(n388), .ZN(n387) );
  AND2_X1 U490 ( .A1(n748), .A2(KEYINPUT65), .ZN(n385) );
  XNOR2_X2 U491 ( .A(n434), .B(KEYINPUT89), .ZN(n388) );
  NAND2_X1 U492 ( .A1(n394), .A2(n377), .ZN(n555) );
  OR2_X2 U493 ( .A1(n394), .A2(n389), .ZN(n554) );
  INV_X1 U494 ( .A(KEYINPUT69), .ZN(n389) );
  XNOR2_X1 U495 ( .A(n394), .B(G122), .ZN(n771) );
  XNOR2_X2 U496 ( .A(n552), .B(n375), .ZN(n394) );
  NAND2_X1 U497 ( .A1(n543), .A2(n373), .ZN(n391) );
  XNOR2_X2 U498 ( .A(n392), .B(G146), .ZN(n521) );
  XNOR2_X1 U499 ( .A(n392), .B(KEYINPUT123), .ZN(n760) );
  XNOR2_X2 U500 ( .A(n402), .B(n507), .ZN(n392) );
  NOR2_X1 U501 ( .A1(n691), .A2(n393), .ZN(n561) );
  XNOR2_X1 U502 ( .A(n393), .B(KEYINPUT1), .ZN(n547) );
  NOR2_X1 U503 ( .A1(n607), .A2(n393), .ZN(n609) );
  NAND2_X1 U504 ( .A1(n395), .A2(n394), .ZN(n576) );
  NOR2_X1 U505 ( .A1(n656), .A2(n396), .ZN(n395) );
  NAND2_X1 U506 ( .A1(n655), .A2(n389), .ZN(n396) );
  XNOR2_X1 U507 ( .A(n398), .B(n549), .ZN(n714) );
  NAND2_X1 U508 ( .A1(n548), .A2(n558), .ZN(n398) );
  NOR2_X2 U509 ( .A1(n547), .A2(n691), .ZN(n558) );
  XNOR2_X2 U510 ( .A(n545), .B(n544), .ZN(n655) );
  NAND2_X1 U511 ( .A1(n615), .A2(n399), .ZN(n630) );
  XNOR2_X1 U512 ( .A(n613), .B(n614), .ZN(n399) );
  NAND2_X1 U513 ( .A1(n421), .A2(n420), .ZN(n400) );
  XNOR2_X1 U514 ( .A(n635), .B(KEYINPUT113), .ZN(n418) );
  XNOR2_X1 U515 ( .A(n589), .B(KEYINPUT108), .ZN(n419) );
  XNOR2_X1 U516 ( .A(n561), .B(KEYINPUT98), .ZN(n598) );
  XNOR2_X2 U517 ( .A(n605), .B(n540), .ZN(n588) );
  XNOR2_X2 U518 ( .A(n590), .B(KEYINPUT19), .ZN(n467) );
  NOR2_X1 U519 ( .A1(n740), .A2(G902), .ZN(n499) );
  XNOR2_X1 U520 ( .A(n497), .B(n498), .ZN(n740) );
  NAND2_X1 U521 ( .A1(n422), .A2(n580), .ZN(n421) );
  NOR2_X1 U522 ( .A1(n405), .A2(n369), .ZN(n408) );
  NAND2_X1 U523 ( .A1(n618), .A2(n617), .ZN(n679) );
  NAND2_X1 U524 ( .A1(n408), .A2(n406), .ZN(n413) );
  OR2_X1 U525 ( .A1(n618), .A2(n407), .ZN(n406) );
  AND2_X1 U526 ( .A1(n598), .A2(n365), .ZN(n416) );
  NOR2_X1 U527 ( .A1(n418), .A2(n590), .ZN(n591) );
  INV_X2 U528 ( .A(n587), .ZN(n694) );
  XNOR2_X2 U529 ( .A(n441), .B(G125), .ZN(n481) );
  NAND2_X1 U530 ( .A1(n645), .A2(n378), .ZN(n420) );
  INV_X1 U531 ( .A(n645), .ZN(n422) );
  NAND2_X1 U532 ( .A1(n733), .A2(n431), .ZN(n430) );
  INV_X1 U533 ( .A(n513), .ZN(n431) );
  NAND2_X1 U534 ( .A1(n773), .A2(n774), .ZN(n613) );
  XNOR2_X2 U535 ( .A(n432), .B(KEYINPUT40), .ZN(n773) );
  NAND2_X1 U536 ( .A1(n640), .A2(n371), .ZN(n432) );
  XNOR2_X1 U537 ( .A(n603), .B(n602), .ZN(n640) );
  XNOR2_X1 U538 ( .A(n631), .B(KEYINPUT48), .ZN(n433) );
  NAND2_X1 U539 ( .A1(n433), .A2(n372), .ZN(n434) );
  BUF_X1 U540 ( .A(n739), .Z(n743) );
  INV_X1 U541 ( .A(n605), .ZN(n593) );
  BUF_X1 U542 ( .A(n605), .Z(n562) );
  AND2_X1 U543 ( .A1(n565), .A2(n564), .ZN(n435) );
  XNOR2_X1 U544 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n436) );
  XNOR2_X1 U545 ( .A(KEYINPUT93), .B(KEYINPUT33), .ZN(n549) );
  INV_X1 U546 ( .A(G104), .ZN(n482) );
  BUF_X1 U547 ( .A(n593), .Z(n698) );
  INV_X1 U548 ( .A(KEYINPUT112), .ZN(n608) );
  INV_X1 U549 ( .A(n747), .ZN(n652) );
  INV_X1 U550 ( .A(KEYINPUT42), .ZN(n611) );
  XNOR2_X1 U551 ( .A(n612), .B(n611), .ZN(n774) );
  NAND2_X1 U552 ( .A1(n492), .A2(G224), .ZN(n437) );
  XNOR2_X1 U553 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U554 ( .A(n440), .B(n488), .ZN(n444) );
  INV_X1 U555 ( .A(G146), .ZN(n441) );
  XNOR2_X1 U556 ( .A(n481), .B(n442), .ZN(n443) );
  XNOR2_X1 U557 ( .A(n444), .B(n443), .ZN(n447) );
  XNOR2_X1 U558 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n446) );
  XNOR2_X1 U559 ( .A(n754), .B(n446), .ZN(n510) );
  XNOR2_X1 U560 ( .A(n447), .B(n510), .ZN(n453) );
  XNOR2_X1 U561 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U562 ( .A(n451), .B(n450), .ZN(n518) );
  XNOR2_X1 U563 ( .A(KEYINPUT16), .B(G122), .ZN(n452) );
  XNOR2_X1 U564 ( .A(n518), .B(n452), .ZN(n753) );
  XNOR2_X1 U565 ( .A(KEYINPUT15), .B(G902), .ZN(n500) );
  INV_X1 U566 ( .A(n500), .ZN(n642) );
  NOR2_X1 U567 ( .A1(G237), .A2(G902), .ZN(n454) );
  XOR2_X1 U568 ( .A(KEYINPUT82), .B(n454), .Z(n460) );
  NAND2_X1 U569 ( .A1(n460), .A2(G210), .ZN(n457) );
  INV_X1 U570 ( .A(KEYINPUT85), .ZN(n455) );
  XNOR2_X1 U571 ( .A(n455), .B(KEYINPUT95), .ZN(n456) );
  XNOR2_X1 U572 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X2 U573 ( .A(n459), .B(n458), .ZN(n600) );
  NAND2_X1 U574 ( .A1(n460), .A2(G214), .ZN(n461) );
  XNOR2_X1 U575 ( .A(n461), .B(KEYINPUT96), .ZN(n706) );
  NAND2_X1 U576 ( .A1(G234), .A2(G237), .ZN(n462) );
  XNOR2_X1 U577 ( .A(n462), .B(KEYINPUT14), .ZN(n464) );
  NAND2_X1 U578 ( .A1(G952), .A2(n464), .ZN(n720) );
  NOR2_X1 U579 ( .A1(G953), .A2(n720), .ZN(n584) );
  AND2_X1 U580 ( .A1(G953), .A2(G902), .ZN(n463) );
  NAND2_X1 U581 ( .A1(n464), .A2(n463), .ZN(n581) );
  NOR2_X1 U582 ( .A1(G898), .A2(n581), .ZN(n465) );
  OR2_X1 U583 ( .A1(n584), .A2(n465), .ZN(n466) );
  NAND2_X1 U584 ( .A1(n467), .A2(n366), .ZN(n468) );
  XNOR2_X2 U585 ( .A(n468), .B(KEYINPUT0), .ZN(n563) );
  XOR2_X1 U586 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n470) );
  NOR2_X1 U587 ( .A1(G953), .A2(G237), .ZN(n514) );
  NAND2_X1 U588 ( .A1(G214), .A2(n514), .ZN(n469) );
  XNOR2_X1 U589 ( .A(n470), .B(n469), .ZN(n474) );
  XOR2_X1 U590 ( .A(KEYINPUT12), .B(G122), .Z(n472) );
  XNOR2_X1 U591 ( .A(G113), .B(G140), .ZN(n471) );
  XNOR2_X1 U592 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U593 ( .A(n474), .B(n473), .ZN(n480) );
  NAND2_X1 U594 ( .A1(n475), .A2(KEYINPUT71), .ZN(n478) );
  NAND2_X1 U595 ( .A1(n476), .A2(G131), .ZN(n477) );
  NAND2_X2 U596 ( .A1(n478), .A2(n477), .ZN(n505) );
  XNOR2_X1 U597 ( .A(n505), .B(G143), .ZN(n479) );
  XNOR2_X1 U598 ( .A(n480), .B(n479), .ZN(n484) );
  XNOR2_X1 U599 ( .A(n526), .B(n482), .ZN(n483) );
  XNOR2_X1 U600 ( .A(n484), .B(n483), .ZN(n659) );
  NOR2_X1 U601 ( .A1(G902), .A2(n659), .ZN(n487) );
  XNOR2_X1 U602 ( .A(KEYINPUT13), .B(KEYINPUT103), .ZN(n485) );
  XOR2_X1 U603 ( .A(KEYINPUT9), .B(G122), .Z(n490) );
  XNOR2_X1 U604 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U605 ( .A(n507), .B(n491), .ZN(n498) );
  XOR2_X1 U606 ( .A(KEYINPUT7), .B(KEYINPUT104), .Z(n496) );
  NAND2_X1 U607 ( .A1(G234), .A2(n762), .ZN(n493) );
  XNOR2_X1 U608 ( .A(n493), .B(n494), .ZN(n528) );
  NAND2_X1 U609 ( .A1(G217), .A2(n528), .ZN(n495) );
  XNOR2_X1 U610 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U611 ( .A(G478), .B(n499), .ZN(n566) );
  NAND2_X1 U612 ( .A1(n568), .A2(n566), .ZN(n709) );
  NAND2_X1 U613 ( .A1(n500), .A2(G234), .ZN(n501) );
  XNOR2_X1 U614 ( .A(n501), .B(KEYINPUT20), .ZN(n536) );
  AND2_X1 U615 ( .A1(n536), .A2(G221), .ZN(n503) );
  INV_X1 U616 ( .A(KEYINPUT21), .ZN(n502) );
  XNOR2_X1 U617 ( .A(n503), .B(n502), .ZN(n585) );
  OR2_X1 U618 ( .A1(n709), .A2(n585), .ZN(n504) );
  NAND2_X1 U619 ( .A1(G227), .A2(n762), .ZN(n508) );
  XOR2_X1 U620 ( .A(n508), .B(G101), .Z(n509) );
  XNOR2_X1 U621 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U622 ( .A(KEYINPUT72), .B(G140), .Z(n527) );
  XNOR2_X1 U623 ( .A(n511), .B(n527), .ZN(n512) );
  XNOR2_X1 U624 ( .A(KEYINPUT74), .B(G469), .ZN(n513) );
  AND2_X1 U625 ( .A1(n514), .A2(G210), .ZN(n517) );
  XOR2_X1 U626 ( .A(KEYINPUT83), .B(KEYINPUT99), .Z(n515) );
  XNOR2_X1 U627 ( .A(n515), .B(KEYINPUT5), .ZN(n516) );
  XNOR2_X1 U628 ( .A(n517), .B(n516), .ZN(n519) );
  XNOR2_X1 U629 ( .A(n519), .B(n518), .ZN(n520) );
  NAND2_X1 U630 ( .A1(n647), .A2(n427), .ZN(n525) );
  XNOR2_X1 U631 ( .A(KEYINPUT78), .B(KEYINPUT100), .ZN(n523) );
  INV_X1 U632 ( .A(G472), .ZN(n522) );
  XNOR2_X1 U633 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X2 U634 ( .A(n525), .B(n524), .ZN(n605) );
  XNOR2_X1 U635 ( .A(n527), .B(n526), .ZN(n759) );
  NAND2_X1 U636 ( .A1(G221), .A2(n528), .ZN(n533) );
  XOR2_X1 U637 ( .A(G110), .B(G119), .Z(n530) );
  XNOR2_X1 U638 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U639 ( .A(n534), .B(n759), .ZN(n744) );
  NOR2_X1 U640 ( .A1(n744), .A2(G902), .ZN(n535) );
  INV_X1 U641 ( .A(n535), .ZN(n539) );
  NAND2_X1 U642 ( .A1(n536), .A2(G217), .ZN(n537) );
  INV_X1 U643 ( .A(KEYINPUT6), .ZN(n540) );
  NOR2_X1 U644 ( .A1(n692), .A2(n694), .ZN(n541) );
  AND2_X1 U645 ( .A1(n588), .A2(n541), .ZN(n542) );
  NAND2_X1 U646 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U647 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n544) );
  INV_X1 U648 ( .A(n655), .ZN(n546) );
  NOR2_X1 U649 ( .A1(n656), .A2(n546), .ZN(n557) );
  INV_X1 U650 ( .A(n585), .ZN(n695) );
  INV_X1 U651 ( .A(n588), .ZN(n548) );
  XNOR2_X1 U652 ( .A(n550), .B(KEYINPUT34), .ZN(n551) );
  NAND2_X1 U653 ( .A1(n551), .A2(n617), .ZN(n552) );
  INV_X1 U654 ( .A(KEYINPUT44), .ZN(n553) );
  NAND2_X1 U655 ( .A1(n554), .A2(n555), .ZN(n556) );
  NAND2_X1 U656 ( .A1(n558), .A2(n698), .ZN(n701) );
  NOR2_X1 U657 ( .A1(n701), .A2(n563), .ZN(n560) );
  XNOR2_X1 U658 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n559) );
  XNOR2_X1 U659 ( .A(n560), .B(n559), .ZN(n684) );
  AND2_X1 U660 ( .A1(n562), .A2(n598), .ZN(n565) );
  INV_X1 U661 ( .A(n563), .ZN(n564) );
  NOR2_X1 U662 ( .A1(n684), .A2(n435), .ZN(n569) );
  INV_X1 U663 ( .A(n566), .ZN(n567) );
  AND2_X1 U664 ( .A1(n568), .A2(n567), .ZN(n683) );
  XOR2_X1 U665 ( .A(n711), .B(KEYINPUT87), .Z(n620) );
  OR2_X1 U666 ( .A1(n569), .A2(n620), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n588), .A2(n694), .ZN(n570) );
  NOR2_X1 U668 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U669 ( .A(n572), .B(KEYINPUT105), .ZN(n772) );
  NAND2_X1 U670 ( .A1(n573), .A2(n772), .ZN(n574) );
  NOR2_X1 U671 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U672 ( .A1(n576), .A2(KEYINPUT44), .ZN(n577) );
  NAND2_X1 U673 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X2 U674 ( .A(n579), .B(KEYINPUT45), .ZN(n645) );
  XOR2_X1 U675 ( .A(KEYINPUT107), .B(n581), .Z(n582) );
  NOR2_X1 U676 ( .A1(G900), .A2(n582), .ZN(n583) );
  NOR2_X1 U677 ( .A1(n584), .A2(n583), .ZN(n597) );
  NOR2_X1 U678 ( .A1(n585), .A2(n597), .ZN(n586) );
  NAND2_X1 U679 ( .A1(n364), .A2(n586), .ZN(n604) );
  NOR2_X1 U680 ( .A1(n588), .A2(n604), .ZN(n589) );
  XNOR2_X1 U681 ( .A(n591), .B(KEYINPUT36), .ZN(n592) );
  INV_X1 U682 ( .A(n692), .ZN(n632) );
  XOR2_X1 U683 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n614) );
  NAND2_X1 U684 ( .A1(n593), .A2(n706), .ZN(n595) );
  XNOR2_X1 U685 ( .A(n595), .B(n594), .ZN(n596) );
  XOR2_X1 U686 ( .A(KEYINPUT38), .B(KEYINPUT81), .Z(n601) );
  INV_X1 U687 ( .A(KEYINPUT39), .ZN(n602) );
  NOR2_X1 U688 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U689 ( .A(KEYINPUT28), .B(n606), .Z(n607) );
  XNOR2_X1 U690 ( .A(n609), .B(n608), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n365), .A2(n706), .ZN(n710) );
  NOR2_X1 U692 ( .A1(n710), .A2(n709), .ZN(n610) );
  XNOR2_X1 U693 ( .A(n610), .B(KEYINPUT41), .ZN(n721) );
  NOR2_X1 U694 ( .A1(n622), .A2(n721), .ZN(n612) );
  INV_X1 U695 ( .A(n600), .ZN(n638) );
  NAND2_X1 U696 ( .A1(n711), .A2(KEYINPUT47), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n621), .B(KEYINPUT80), .ZN(n624) );
  INV_X1 U698 ( .A(n622), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n623), .A2(n467), .ZN(n625) );
  INV_X1 U700 ( .A(n625), .ZN(n680) );
  NAND2_X1 U701 ( .A1(n624), .A2(n680), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n625), .A2(KEYINPUT47), .ZN(n626) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT79), .ZN(n629) );
  NOR2_X2 U704 ( .A1(n630), .A2(n629), .ZN(n631) );
  INV_X1 U705 ( .A(n706), .ZN(n633) );
  NOR2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U708 ( .A(KEYINPUT109), .B(n636), .ZN(n637) );
  XOR2_X1 U709 ( .A(KEYINPUT43), .B(n637), .Z(n639) );
  AND2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n657) );
  AND2_X1 U711 ( .A1(n640), .A2(n683), .ZN(n689) );
  NOR2_X1 U712 ( .A1(n657), .A2(n689), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n642), .A2(KEYINPUT2), .ZN(n643) );
  BUF_X2 U714 ( .A(n645), .Z(n748) );
  NAND2_X1 U715 ( .A1(n739), .A2(G472), .ZN(n649) );
  XOR2_X1 U716 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(n648) );
  INV_X1 U718 ( .A(G952), .ZN(n651) );
  AND2_X1 U719 ( .A1(n651), .A2(G953), .ZN(n747) );
  NAND2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U721 ( .A(n654), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U722 ( .A(n359), .B(G119), .ZN(G21) );
  XOR2_X1 U723 ( .A(n656), .B(G110), .Z(G12) );
  XOR2_X1 U724 ( .A(n657), .B(G140), .Z(G42) );
  NAND2_X1 U725 ( .A1(n739), .A2(G475), .ZN(n661) );
  XOR2_X1 U726 ( .A(KEYINPUT94), .B(KEYINPUT59), .Z(n658) );
  XNOR2_X1 U727 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n663) );
  NAND2_X1 U728 ( .A1(n739), .A2(G210), .ZN(n668) );
  XOR2_X1 U729 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n665) );
  XOR2_X1 U730 ( .A(KEYINPUT91), .B(KEYINPUT56), .Z(n670) );
  NAND2_X1 U731 ( .A1(n435), .A2(n371), .ZN(n672) );
  XNOR2_X1 U732 ( .A(n672), .B(G104), .ZN(G6) );
  XOR2_X1 U733 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n674) );
  NAND2_X1 U734 ( .A1(n435), .A2(n683), .ZN(n673) );
  XNOR2_X1 U735 ( .A(n674), .B(n673), .ZN(n676) );
  XOR2_X1 U736 ( .A(G107), .B(KEYINPUT26), .Z(n675) );
  XNOR2_X1 U737 ( .A(n676), .B(n675), .ZN(G9) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n678) );
  NAND2_X1 U739 ( .A1(n680), .A2(n683), .ZN(n677) );
  XNOR2_X1 U740 ( .A(n678), .B(n677), .ZN(G30) );
  XNOR2_X1 U741 ( .A(G143), .B(n679), .ZN(G45) );
  NAND2_X1 U742 ( .A1(n680), .A2(n371), .ZN(n681) );
  XNOR2_X1 U743 ( .A(n681), .B(G146), .ZN(G48) );
  NAND2_X1 U744 ( .A1(n684), .A2(n371), .ZN(n682) );
  XNOR2_X1 U745 ( .A(n682), .B(G113), .ZN(G15) );
  NAND2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U747 ( .A(n685), .B(G116), .ZN(G18) );
  XOR2_X1 U748 ( .A(KEYINPUT116), .B(KEYINPUT37), .Z(n686) );
  XNOR2_X1 U749 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U750 ( .A(G125), .B(n688), .ZN(G27) );
  XNOR2_X1 U751 ( .A(G134), .B(n689), .ZN(n690) );
  XNOR2_X1 U752 ( .A(n690), .B(KEYINPUT117), .ZN(G36) );
  XOR2_X1 U753 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n704) );
  NAND2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U755 ( .A(n693), .B(KEYINPUT50), .ZN(n700) );
  NOR2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U757 ( .A(KEYINPUT49), .B(n696), .Z(n697) );
  NOR2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U759 ( .A1(n700), .A2(n699), .ZN(n702) );
  NAND2_X1 U760 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U761 ( .A(n704), .B(n703), .Z(n705) );
  NOR2_X1 U762 ( .A1(n721), .A2(n705), .ZN(n717) );
  NOR2_X1 U763 ( .A1(n365), .A2(n706), .ZN(n707) );
  XOR2_X1 U764 ( .A(KEYINPUT119), .B(n707), .Z(n708) );
  NOR2_X1 U765 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U767 ( .A1(n713), .A2(n712), .ZN(n715) );
  NOR2_X1 U768 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U770 ( .A(n718), .B(KEYINPUT52), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n723) );
  NOR2_X1 U772 ( .A1(n721), .A2(n714), .ZN(n722) );
  NOR2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n729) );
  NAND2_X1 U774 ( .A1(n748), .A2(n761), .ZN(n725) );
  INV_X1 U775 ( .A(KEYINPUT2), .ZN(n724) );
  NAND2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n727) );
  NAND2_X1 U777 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U779 ( .A1(G953), .A2(n730), .ZN(n732) );
  XNOR2_X1 U780 ( .A(KEYINPUT53), .B(KEYINPUT120), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(G75) );
  XOR2_X1 U782 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n735) );
  XNOR2_X1 U783 ( .A(n733), .B(KEYINPUT121), .ZN(n734) );
  XNOR2_X1 U784 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U785 ( .A1(n739), .A2(G469), .ZN(n736) );
  XOR2_X1 U786 ( .A(n737), .B(n736), .Z(n738) );
  NOR2_X1 U787 ( .A1(n747), .A2(n738), .ZN(G54) );
  NAND2_X1 U788 ( .A1(n743), .A2(G478), .ZN(n741) );
  XNOR2_X1 U789 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U790 ( .A1(n747), .A2(n742), .ZN(G63) );
  NAND2_X1 U791 ( .A1(n743), .A2(G217), .ZN(n745) );
  XNOR2_X1 U792 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U793 ( .A1(n747), .A2(n746), .ZN(G66) );
  NAND2_X1 U794 ( .A1(n748), .A2(n762), .ZN(n752) );
  NAND2_X1 U795 ( .A1(G953), .A2(G224), .ZN(n749) );
  XNOR2_X1 U796 ( .A(KEYINPUT61), .B(n749), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n750), .A2(G898), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n752), .A2(n751), .ZN(n758) );
  XOR2_X1 U799 ( .A(n754), .B(n753), .Z(n756) );
  NOR2_X1 U800 ( .A1(n762), .A2(G898), .ZN(n755) );
  NOR2_X1 U801 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U802 ( .A(n758), .B(n757), .ZN(G69) );
  XOR2_X1 U803 ( .A(n760), .B(n759), .Z(n765) );
  XOR2_X1 U804 ( .A(n765), .B(n761), .Z(n763) );
  NAND2_X1 U805 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U806 ( .A(n764), .B(KEYINPUT124), .ZN(n769) );
  XNOR2_X1 U807 ( .A(G227), .B(n765), .ZN(n766) );
  NAND2_X1 U808 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U809 ( .A1(G953), .A2(n767), .ZN(n768) );
  NAND2_X1 U810 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U811 ( .A(KEYINPUT125), .B(n770), .Z(G72) );
  XNOR2_X1 U812 ( .A(n771), .B(KEYINPUT126), .ZN(G24) );
  XNOR2_X1 U813 ( .A(G101), .B(n772), .ZN(G3) );
  XNOR2_X1 U814 ( .A(n773), .B(G131), .ZN(G33) );
  XNOR2_X1 U815 ( .A(G137), .B(n774), .ZN(G39) );
endmodule

