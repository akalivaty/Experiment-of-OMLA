//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(G8gat), .Z(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n207), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n208));
  XOR2_X1   g007(.A(KEYINPUT14), .B(G29gat), .Z(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(G36gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT92), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n210), .A2(new_n212), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n210), .A2(KEYINPUT92), .A3(new_n212), .A4(new_n213), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n216), .A2(KEYINPUT17), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n206), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT17), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n206), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n220), .A2(new_n223), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT18), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT93), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n225), .A2(KEYINPUT93), .A3(KEYINPUT18), .A4(new_n226), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT18), .B1(new_n225), .B2(new_n226), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n206), .B(new_n221), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n226), .B(KEYINPUT13), .Z(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G141gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G197gat), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT11), .B(G169gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n242), .B(KEYINPUT12), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n243), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n231), .A2(new_n245), .A3(new_n237), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250));
  INV_X1    g049(.A(G127gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(G134gat), .ZN(new_n252));
  INV_X1    g051(.A(G134gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(G127gat), .ZN(new_n254));
  OAI22_X1  g053(.A1(new_n250), .A2(KEYINPUT1), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G120gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G113gat), .ZN(new_n257));
  INV_X1    g056(.A(G113gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G120gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n255), .A2(new_n263), .A3(KEYINPUT70), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT70), .B1(new_n255), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n267));
  INV_X1    g066(.A(G169gat), .ZN(new_n268));
  INV_X1    g067(.A(G176gat), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT23), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n269), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(new_n268), .A3(new_n269), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(KEYINPUT23), .A3(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT24), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n283));
  INV_X1    g082(.A(G183gat), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n278), .A2(KEYINPUT68), .A3(new_n279), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n282), .A2(new_n283), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT65), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n290), .A2(new_n291), .A3(new_n280), .A4(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n270), .A2(new_n271), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n268), .A2(KEYINPUT23), .ZN(new_n294));
  NOR2_X1   g093(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(new_n293), .A3(new_n298), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n277), .A2(new_n288), .B1(new_n299), .B2(new_n267), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n284), .A2(KEYINPUT27), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT27), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G183gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n303), .A3(new_n285), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n304), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT69), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT26), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n274), .A2(new_n275), .A3(new_n308), .A4(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n307), .B1(new_n268), .B2(new_n269), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n271), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n305), .A2(new_n306), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n266), .B1(new_n300), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT70), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n261), .B1(new_n262), .B2(new_n260), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n255), .A2(new_n263), .A3(KEYINPUT70), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n299), .A2(new_n267), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n288), .A2(new_n276), .A3(new_n272), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n326), .A3(new_n315), .ZN(new_n327));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n328), .B(KEYINPUT64), .Z(new_n329));
  NAND3_X1  g128(.A1(new_n317), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT32), .ZN(new_n331));
  XOR2_X1   g130(.A(G15gat), .B(G43gat), .Z(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT71), .ZN(new_n333));
  XNOR2_X1  g132(.A(G71gat), .B(G99gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n331), .B1(KEYINPUT33), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n331), .A2(new_n338), .A3(new_n335), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n335), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(new_n330), .B2(KEYINPUT32), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(KEYINPUT72), .A3(new_n338), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n336), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n317), .A2(new_n327), .ZN(new_n346));
  INV_X1    g145(.A(new_n329), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT74), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n336), .ZN(new_n352));
  INV_X1    g151(.A(new_n344), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT72), .B1(new_n343), .B2(new_n338), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n356));
  INV_X1    g155(.A(new_n350), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n351), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(G22gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G141gat), .ZN(new_n365));
  INV_X1    g164(.A(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT81), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n371), .A3(new_n368), .ZN(new_n372));
  AND2_X1   g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT2), .ZN(new_n375));
  INV_X1    g174(.A(G155gat), .ZN(new_n376));
  INV_X1    g175(.A(G162gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n370), .A2(new_n372), .A3(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NOR3_X1   g181(.A1(KEYINPUT79), .A2(G155gat), .A3(G162gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n374), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT80), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n376), .A3(new_n377), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n373), .B1(new_n387), .B2(new_n381), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n367), .B(new_n368), .C1(new_n373), .C2(new_n375), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n380), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G211gat), .B(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G218gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT75), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(G218gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT22), .B1(new_n402), .B2(G211gat), .ZN(new_n403));
  XOR2_X1   g202(.A(G197gat), .B(G204gat), .Z(new_n404));
  OAI21_X1  g203(.A(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT22), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT75), .B(G218gat), .ZN(new_n407));
  INV_X1    g206(.A(G211gat), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n404), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n396), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n405), .A2(KEYINPUT76), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT76), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n413), .B(new_n397), .C1(new_n403), .C2(new_n404), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT77), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n417), .A3(new_n414), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n395), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT29), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n412), .A2(new_n420), .A3(new_n414), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n393), .B1(new_n421), .B2(new_n394), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n364), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n388), .A2(new_n389), .ZN(new_n424));
  AOI211_X1 g223(.A(KEYINPUT80), .B(new_n373), .C1(new_n387), .C2(new_n381), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n392), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n370), .A2(new_n372), .A3(new_n379), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(new_n405), .B2(new_n411), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n429), .A2(KEYINPUT85), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n394), .B1(new_n429), .B2(KEYINPUT85), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n394), .A3(new_n427), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n420), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n412), .A2(new_n417), .A3(new_n414), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n417), .B1(new_n412), .B2(new_n414), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n437), .A3(new_n363), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT31), .B(G50gat), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n423), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n423), .B2(new_n438), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n362), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n438), .ZN(new_n444));
  INV_X1    g243(.A(new_n422), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n363), .B1(new_n445), .B2(new_n437), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n439), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n423), .A2(new_n438), .A3(new_n440), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n361), .A3(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n350), .B(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n443), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n249), .B1(new_n359), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n443), .A2(new_n449), .A3(new_n450), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n453), .A2(KEYINPUT89), .A3(new_n351), .A4(new_n358), .ZN(new_n454));
  INV_X1    g253(.A(G226gat), .ZN(new_n455));
  INV_X1    g254(.A(G233gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(KEYINPUT29), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n326), .B2(new_n315), .ZN(new_n459));
  INV_X1    g258(.A(new_n457), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n288), .A2(new_n276), .A3(new_n272), .ZN(new_n461));
  INV_X1    g260(.A(new_n297), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(new_n295), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n463), .A2(new_n294), .B1(new_n270), .B2(new_n271), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT25), .B1(new_n464), .B2(new_n292), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n315), .B(new_n460), .C1(new_n461), .C2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OAI22_X1  g266(.A1(new_n459), .A2(new_n467), .B1(new_n435), .B2(new_n436), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT78), .ZN(new_n469));
  OAI22_X1  g268(.A1(new_n300), .A2(new_n316), .B1(KEYINPUT29), .B2(new_n457), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n416), .A2(new_n470), .A3(new_n418), .A4(new_n466), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n416), .A2(new_n418), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n466), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(KEYINPUT78), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G8gat), .B(G36gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(G64gat), .B(G92gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n472), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT30), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n475), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n478), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n481), .B(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n426), .A2(new_n321), .A3(new_n427), .A4(new_n322), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT4), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n319), .A2(new_n320), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n393), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n485), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n428), .A2(KEYINPUT3), .ZN(new_n492));
  INV_X1    g291(.A(new_n489), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n433), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n393), .A2(new_n266), .A3(new_n488), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n426), .A2(new_n427), .A3(new_n489), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT83), .ZN(new_n498));
  NAND2_X1  g297(.A1(G225gat), .A2(G233gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n491), .A2(new_n494), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT84), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n495), .A2(new_n497), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n489), .B1(new_n428), .B2(KEYINPUT3), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n504), .A2(new_n485), .B1(new_n433), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT84), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n506), .A2(new_n507), .A3(new_n498), .A4(new_n501), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n496), .A2(new_n488), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n393), .A2(new_n266), .A3(KEYINPUT4), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n494), .A2(new_n510), .A3(new_n499), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n428), .A2(new_n493), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n496), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n515), .B2(new_n500), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n509), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G1gat), .B(G29gat), .Z(new_n520));
  XNOR2_X1  g319(.A(G57gat), .B(G85gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n522), .B(new_n523), .Z(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n517), .B1(new_n503), .B2(new_n508), .ZN(new_n526));
  INV_X1    g325(.A(new_n524), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT6), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n519), .A2(KEYINPUT6), .A3(new_n524), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n484), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n452), .A2(new_n454), .A3(new_n531), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n532), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT90), .B1(new_n532), .B2(KEYINPUT35), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n355), .A2(new_n357), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n536), .A2(new_n451), .A3(KEYINPUT35), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n531), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n351), .A2(KEYINPUT36), .A3(new_n358), .A4(new_n450), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n450), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n443), .A2(new_n449), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n531), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT86), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n484), .A2(new_n525), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT40), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n506), .A2(new_n498), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT39), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(new_n500), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n527), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n514), .A2(new_n496), .A3(new_n499), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT39), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n552), .B2(new_n500), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n551), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n558), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n560), .A2(KEYINPUT40), .A3(new_n527), .A4(new_n554), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n549), .B1(new_n550), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n559), .A2(new_n561), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n564), .A2(KEYINPUT86), .A3(new_n525), .A4(new_n484), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n529), .A2(new_n530), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n478), .B1(new_n482), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(new_n569), .B2(new_n482), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT38), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT87), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n471), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n468), .A2(KEYINPUT88), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT88), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n473), .A2(new_n576), .A3(new_n474), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n471), .A2(new_n573), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT38), .B1(new_n579), .B2(KEYINPUT37), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n570), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n572), .A2(new_n483), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n546), .B1(new_n568), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n548), .B1(new_n566), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT91), .B1(new_n540), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n532), .A2(KEYINPUT35), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT90), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n539), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n532), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n248), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G71gat), .B(G78gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT94), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n600));
  AND2_X1   g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n251), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n224), .B1(new_n599), .B2(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n602), .B(G127gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT95), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G155gat), .ZN(new_n611));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n605), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n605), .B2(new_n608), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G85gat), .ZN(new_n617));
  INV_X1    g416(.A(G92gat), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT96), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(G85gat), .A3(G92gat), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n621), .A3(KEYINPUT7), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n623));
  OAI211_X1 g422(.A(KEYINPUT96), .B(new_n623), .C1(new_n617), .C2(new_n618), .ZN(new_n624));
  NAND2_X1  g423(.A1(G99gat), .A2(G106gat), .ZN(new_n625));
  AOI22_X1  g424(.A1(KEYINPUT8), .A2(new_n625), .B1(new_n617), .B2(new_n618), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n622), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  XOR2_X1   g427(.A(G99gat), .B(G106gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n221), .ZN(new_n631));
  NAND3_X1  g430(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n629), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n628), .B(new_n634), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n635), .A2(new_n223), .A3(new_n219), .ZN(new_n636));
  XNOR2_X1  g435(.A(G190gat), .B(G218gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  NOR3_X1   g438(.A1(new_n633), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n643));
  INV_X1    g442(.A(G232gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n456), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n642), .B(new_n645), .Z(new_n646));
  OAI21_X1  g445(.A(new_n639), .B1(new_n633), .B2(new_n636), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n641), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n641), .B2(new_n647), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n598), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n630), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n599), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT10), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n655));
  INV_X1    g454(.A(G230gat), .ZN(new_n656));
  OAI22_X1  g455(.A1(new_n654), .A2(new_n655), .B1(new_n656), .B2(new_n456), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n456), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n652), .A2(new_n653), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n661), .B(new_n662), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n657), .A2(new_n659), .A3(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n616), .A2(new_n650), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n593), .A2(new_n568), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT100), .B(G1gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1324gat));
  NAND2_X1  g472(.A1(new_n593), .A2(new_n670), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT16), .B(G8gat), .Z(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n484), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n484), .ZN(new_n678));
  OAI21_X1  g477(.A(G8gat), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  MUX2_X1   g479(.A(new_n677), .B(new_n680), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g480(.A(G15gat), .B1(new_n674), .B2(new_n545), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n669), .A2(G15gat), .A3(new_n542), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n593), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n675), .A2(new_n546), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n650), .A2(new_n689), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT91), .B(new_n584), .C1(new_n588), .C2(new_n589), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n586), .A2(new_n587), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n589), .A3(new_n538), .ZN(new_n693));
  INV_X1    g492(.A(new_n584), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n591), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n690), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n689), .B1(new_n590), .B2(new_n650), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n667), .B(KEYINPUT101), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(new_n616), .A3(new_n248), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G29gat), .B1(new_n702), .B2(new_n567), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n704));
  INV_X1    g503(.A(new_n616), .ZN(new_n705));
  INV_X1    g504(.A(new_n650), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n706), .A3(new_n668), .ZN(new_n707));
  AOI211_X1 g506(.A(new_n248), .B(new_n707), .C1(new_n585), .C2(new_n592), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n568), .A2(new_n207), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n704), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n708), .A2(KEYINPUT45), .A3(new_n207), .A4(new_n568), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n703), .A2(new_n711), .A3(new_n712), .ZN(G1328gat));
  OAI21_X1  g512(.A(G36gat), .B1(new_n702), .B2(new_n678), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n678), .A2(G36gat), .ZN(new_n715));
  OR3_X1    g514(.A1(new_n709), .A2(KEYINPUT46), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT46), .B1(new_n709), .B2(new_n715), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(G1329gat));
  INV_X1    g517(.A(new_n545), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n696), .A2(new_n719), .A3(new_n697), .A4(new_n701), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G43gat), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n542), .A2(G43gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n708), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT102), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n720), .A2(G43gat), .B1(new_n708), .B2(new_n722), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n727), .A2(new_n728), .A3(KEYINPUT47), .ZN(new_n729));
  AND4_X1   g528(.A1(KEYINPUT103), .A2(new_n721), .A3(KEYINPUT47), .A4(new_n723), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT103), .B1(new_n727), .B2(KEYINPUT47), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n726), .A2(new_n729), .B1(new_n730), .B2(new_n731), .ZN(G1330gat));
  NAND4_X1  g531(.A1(new_n696), .A2(new_n546), .A3(new_n697), .A4(new_n701), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G50gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT48), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n547), .A2(G50gat), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n734), .B1(new_n709), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n736), .B(new_n739), .ZN(G1331gat));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n700), .A2(new_n248), .A3(new_n616), .A4(new_n650), .ZN(new_n742));
  OR3_X1    g541(.A1(new_n590), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n590), .B2(new_n742), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n567), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(G57gat), .Z(G1332gat));
  AOI21_X1  g546(.A(new_n678), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n743), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT106), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1333gat));
  OAI21_X1  g551(.A(G71gat), .B1(new_n745), .B2(new_n545), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n542), .A2(G71gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n745), .B2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g555(.A1(new_n745), .A2(new_n547), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT107), .B(G78gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n616), .A2(new_n247), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n667), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT108), .Z(new_n762));
  AND2_X1   g561(.A1(new_n698), .A2(new_n762), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n763), .A2(new_n568), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n706), .B(new_n760), .C1(new_n540), .C2(new_n584), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n568), .A2(new_n617), .A3(new_n667), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n764), .A2(new_n617), .B1(new_n768), .B2(new_n769), .ZN(G1336gat));
  NAND4_X1  g569(.A1(new_n696), .A2(new_n484), .A3(new_n697), .A4(new_n762), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n699), .A2(G92gat), .A3(new_n678), .ZN(new_n772));
  AOI22_X1  g571(.A1(G92gat), .A2(new_n771), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1337gat));
  AND2_X1   g574(.A1(new_n763), .A2(new_n719), .ZN(new_n776));
  INV_X1    g575(.A(G99gat), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n667), .A2(new_n777), .A3(new_n535), .A4(new_n450), .ZN(new_n778));
  OAI22_X1  g577(.A1(new_n776), .A2(new_n777), .B1(new_n768), .B2(new_n778), .ZN(G1338gat));
  NOR3_X1   g578(.A1(new_n699), .A2(G106gat), .A3(new_n547), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT110), .Z(new_n781));
  AND2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n765), .A2(new_n766), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n767), .A2(KEYINPUT111), .A3(new_n781), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n696), .A2(new_n546), .A3(new_n697), .A4(new_n762), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT53), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  INV_X1    g591(.A(new_n780), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n768), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n791), .B1(new_n790), .B2(new_n794), .ZN(G1339gat));
  NAND2_X1  g594(.A1(new_n670), .A2(new_n248), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT112), .B1(new_n225), .B2(new_n226), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n233), .A2(new_n235), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n225), .A2(KEYINPUT112), .A3(new_n226), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n797), .B(new_n242), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n246), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n242), .B1(new_n800), .B2(new_n801), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT113), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n652), .A2(new_n653), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT10), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n655), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n658), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n663), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n658), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(KEYINPUT54), .A3(new_n657), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n666), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT55), .B1(new_n812), .B2(new_n814), .ZN(new_n817));
  NOR4_X1   g616(.A1(new_n806), .A2(new_n816), .A3(new_n650), .A4(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n813), .A2(KEYINPUT54), .A3(new_n657), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n664), .B1(new_n657), .B2(KEYINPUT54), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(new_n247), .A3(new_n666), .A4(new_n815), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n803), .A2(new_n667), .A3(new_n805), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n706), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n705), .B1(new_n818), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n536), .B(new_n451), .C1(new_n796), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n568), .A2(new_n678), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831), .B2(new_n248), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n567), .B1(new_n796), .B2(new_n826), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n452), .A2(new_n454), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n484), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n247), .A2(new_n258), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT114), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n832), .A2(new_n839), .ZN(G1340gat));
  AOI21_X1  g639(.A(new_n256), .B1(new_n830), .B2(new_n700), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT115), .Z(new_n842));
  NAND3_X1  g641(.A1(new_n836), .A2(new_n256), .A3(new_n667), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n831), .B2(new_n705), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n836), .A2(new_n251), .A3(new_n616), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1342gat));
  NAND2_X1  g646(.A1(new_n706), .A2(new_n678), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT116), .ZN(new_n849));
  OR4_X1    g648(.A1(G134gat), .A2(new_n834), .A3(new_n835), .A4(new_n849), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n831), .B2(new_n650), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  INV_X1    g653(.A(new_n825), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n816), .A2(new_n650), .A3(new_n817), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n805), .A3(new_n803), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n616), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n669), .A2(new_n247), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT121), .B(new_n568), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n719), .A2(new_n547), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n833), .A2(KEYINPUT121), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n248), .A2(G141gat), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n864), .A2(KEYINPUT122), .A3(new_n678), .A4(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n861), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n833), .B2(KEYINPUT121), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n858), .A2(new_n859), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n567), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n868), .A2(new_n871), .A3(new_n678), .A4(new_n865), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n866), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n828), .A2(new_n719), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT117), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n547), .B1(new_n796), .B2(new_n826), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n824), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n803), .A2(KEYINPUT118), .A3(new_n667), .A4(new_n805), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n822), .A2(KEYINPUT119), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n817), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n247), .A2(new_n666), .A3(new_n815), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n883), .B(new_n884), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n818), .B1(new_n890), .B2(new_n650), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n796), .B1(new_n891), .B2(new_n616), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(new_n546), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n247), .B(new_n881), .C1(new_n893), .C2(new_n880), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT58), .B1(new_n894), .B2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n875), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n875), .B2(new_n895), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(new_n881), .C1(new_n893), .C2(new_n880), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n880), .B1(new_n892), .B2(new_n546), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n880), .B(new_n546), .C1(new_n858), .C2(new_n859), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n877), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT120), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(new_n905), .A3(new_n247), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n868), .A2(new_n871), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n484), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n906), .A2(G141gat), .B1(new_n908), .B2(new_n865), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n897), .A2(new_n898), .B1(new_n899), .B2(new_n909), .ZN(G1344gat));
  NAND2_X1  g709(.A1(new_n366), .A2(KEYINPUT59), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(new_n908), .B2(new_n667), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n893), .A2(new_n880), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT57), .B1(new_n870), .B2(new_n547), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n915), .A2(KEYINPUT59), .A3(new_n667), .A4(new_n877), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n905), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n668), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n918), .B2(KEYINPUT59), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n912), .B1(new_n919), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g719(.A(G155gat), .B1(new_n917), .B2(new_n705), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n908), .A2(new_n376), .A3(new_n616), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n917), .B2(new_n650), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n849), .A2(G162gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n907), .B2(new_n925), .ZN(G1347gat));
  NAND3_X1  g725(.A1(new_n827), .A2(new_n484), .A3(new_n567), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(new_n268), .A3(new_n248), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n870), .A2(new_n568), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n835), .A2(new_n678), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n247), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n928), .B1(new_n933), .B2(new_n268), .ZN(G1348gat));
  OAI21_X1  g733(.A(new_n269), .B1(new_n931), .B2(new_n668), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT124), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n927), .A2(new_n463), .A3(new_n699), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n927), .B2(new_n705), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n616), .A2(new_n301), .A3(new_n303), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n931), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n932), .A2(new_n285), .A3(new_n706), .ZN(new_n943));
  OAI21_X1  g742(.A(G190gat), .B1(new_n927), .B2(new_n650), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  NOR4_X1   g749(.A1(new_n870), .A2(new_n678), .A3(new_n568), .A4(new_n867), .ZN(new_n951));
  AOI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n247), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n719), .A2(new_n678), .A3(new_n568), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n915), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n247), .A2(G197gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1352gat));
  OAI21_X1  g756(.A(G204gat), .B1(new_n954), .B2(new_n699), .ZN(new_n958));
  INV_X1    g757(.A(G204gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n951), .A2(new_n959), .A3(new_n667), .ZN(new_n960));
  AND2_X1   g759(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n961));
  NOR2_X1   g760(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n958), .B(new_n963), .C1(new_n961), .C2(new_n960), .ZN(G1353gat));
  NAND4_X1  g763(.A1(new_n913), .A2(new_n616), .A3(new_n914), .A4(new_n953), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G211gat), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n966), .A2(KEYINPUT63), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(KEYINPUT63), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n408), .A3(new_n616), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT127), .Z(new_n970));
  NAND3_X1  g769(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(G1354gat));
  AOI21_X1  g770(.A(G218gat), .B1(new_n951), .B2(new_n706), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n650), .A2(new_n407), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n955), .B2(new_n973), .ZN(G1355gat));
endmodule


