//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n187));
  NOR2_X1   g001(.A1(G475), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT71), .A4(KEYINPUT16), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT71), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(new_n191), .B2(KEYINPUT16), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n189), .B(new_n194), .C1(new_n195), .C2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n200));
  OR3_X1    g014(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(new_n196), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n189), .B1(new_n202), .B2(new_n194), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT90), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G237), .ZN(new_n205));
  INV_X1    g019(.A(G953), .ZN(new_n206));
  AND4_X1   g020(.A1(G143), .A2(new_n205), .A3(new_n206), .A4(G214), .ZN(new_n207));
  NOR2_X1   g021(.A1(G237), .A2(G953), .ZN(new_n208));
  AOI21_X1  g022(.A(G143), .B1(new_n208), .B2(G214), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n205), .A2(new_n206), .A3(G214), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n208), .A2(G143), .A3(G214), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(new_n211), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n216), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT17), .A3(G131), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n194), .B1(new_n195), .B2(new_n197), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT90), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(new_n198), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n204), .A2(new_n221), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G125), .B(G140), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(new_n189), .ZN(new_n228));
  OAI211_X1 g042(.A(KEYINPUT18), .B(G131), .C1(new_n207), .C2(new_n209), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT18), .A2(G131), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n214), .A2(new_n216), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT87), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n228), .A2(KEYINPUT87), .A3(new_n229), .A4(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G113), .B(G122), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT89), .B(G104), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n226), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT91), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT91), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n226), .A2(new_n242), .A3(new_n236), .A4(new_n239), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(new_n227), .B(KEYINPUT19), .Z(new_n245));
  OR2_X1    g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n210), .A2(new_n247), .A3(new_n217), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n210), .A2(new_n217), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT88), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n246), .A2(new_n223), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n239), .B1(new_n251), .B2(new_n236), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n187), .B(new_n188), .C1(new_n244), .C2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n239), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n236), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n241), .A2(new_n243), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n188), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT92), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n258), .A3(KEYINPUT20), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n213), .A2(G128), .ZN(new_n260));
  XOR2_X1   g074(.A(new_n260), .B(KEYINPUT13), .Z(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT64), .B(G128), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(G134), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G116), .B(G122), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n260), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n265), .B(new_n268), .C1(G134), .C2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT9), .B(G234), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(G217), .A3(new_n206), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G134), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n269), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT14), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n266), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G116), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n279), .A2(G122), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n267), .B1(new_n280), .B2(KEYINPUT14), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n266), .A2(new_n267), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n278), .A2(new_n281), .B1(new_n282), .B2(KEYINPUT94), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(KEYINPUT94), .B2(new_n282), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n270), .B(new_n274), .C1(new_n276), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT95), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n276), .A2(new_n284), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT95), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n270), .A4(new_n274), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n270), .B1(new_n276), .B2(new_n284), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n273), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n286), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G478), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(KEYINPUT15), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n296), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n292), .B2(new_n293), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT92), .B(new_n301), .C1(new_n256), .C2(new_n257), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT93), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n226), .A2(new_n303), .A3(new_n236), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n226), .A2(new_n236), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n239), .B1(new_n305), .B2(KEYINPUT93), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n304), .A2(new_n306), .B1(new_n241), .B2(new_n243), .ZN(new_n307));
  OAI21_X1  g121(.A(G475), .B1(new_n307), .B2(G902), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n259), .A2(new_n300), .A3(new_n302), .A4(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G221), .B1(new_n271), .B2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n206), .A2(G227), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(KEYINPUT75), .ZN(new_n312));
  XNOR2_X1  g126(.A(G110), .B(G140), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n189), .A2(G143), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n213), .A2(G146), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .A4(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n316), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G128), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n315), .B2(KEYINPUT1), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n324));
  INV_X1    g138(.A(G104), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(G107), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n267), .A2(KEYINPUT3), .A3(G104), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n267), .B2(G104), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(KEYINPUT77), .A3(G107), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n328), .A2(new_n329), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n325), .A2(G107), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n267), .A2(G104), .ZN(new_n335));
  OAI21_X1  g149(.A(G101), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n323), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n326), .A2(new_n327), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n331), .A2(new_n332), .ZN(new_n341));
  OAI21_X1  g155(.A(G101), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n342), .A2(KEYINPUT4), .A3(new_n333), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n344), .B(G101), .C1(new_n340), .C2(new_n341), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT0), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(new_n321), .ZN(new_n347));
  NOR2_X1   g161(.A1(KEYINPUT0), .A2(G128), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n319), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n315), .B(new_n316), .C1(new_n346), .C2(new_n321), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n339), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n317), .B1(G143), .B2(new_n189), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n319), .B1(new_n262), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n354), .B1(new_n356), .B2(new_n318), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n333), .A2(new_n358), .A3(new_n336), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n333), .B2(new_n336), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT80), .B(new_n357), .C1(new_n359), .C2(new_n360), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n353), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT11), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n275), .B2(G137), .ZN(new_n367));
  INV_X1    g181(.A(G137), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(KEYINPUT11), .A3(G134), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n275), .A2(G137), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G131), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n367), .A2(new_n369), .A3(new_n215), .A4(new_n370), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n365), .A2(new_n375), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n374), .B(new_n353), .C1(new_n363), .C2(new_n364), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n314), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n314), .B1(new_n365), .B2(new_n375), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n333), .A2(new_n336), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n356), .A3(new_n318), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n375), .B1(new_n381), .B2(new_n337), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT12), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  AOI211_X1 g198(.A(G469), .B(G902), .C1(new_n378), .C2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n352), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n342), .A2(KEYINPUT4), .A3(new_n333), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n386), .A2(new_n387), .B1(new_n337), .B2(new_n338), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n380), .A2(KEYINPUT79), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n333), .A2(new_n358), .A3(new_n336), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT80), .B1(new_n391), .B2(new_n357), .ZN(new_n392));
  INV_X1    g206(.A(new_n364), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n375), .B(new_n388), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n383), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n314), .B(KEYINPUT76), .Z(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n374), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n379), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n400), .A3(G469), .ZN(new_n401));
  INV_X1    g215(.A(G469), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(new_n293), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n310), .B1(new_n385), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n206), .A2(G952), .ZN(new_n407));
  NAND2_X1  g221(.A1(G234), .A2(G237), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(G902), .A3(G953), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT21), .B(G898), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G214), .B1(G237), .B2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT65), .ZN(new_n420));
  INV_X1    g234(.A(G113), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT2), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT2), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G113), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G116), .B(G119), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G119), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G116), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n279), .A2(G119), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT2), .B(G113), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n420), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(new_n432), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n425), .A2(new_n426), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT65), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT81), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n387), .A4(new_n345), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT82), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n429), .B2(KEYINPUT5), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT5), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT5), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n444), .A2(new_n428), .A3(KEYINPUT82), .A4(G116), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n442), .A2(new_n443), .A3(G113), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n436), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n359), .B2(new_n360), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n440), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n341), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n329), .B1(new_n451), .B2(new_n328), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n434), .A2(new_n437), .B1(new_n452), .B2(new_n344), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n439), .B1(new_n453), .B2(new_n387), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n419), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT65), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT65), .B1(new_n435), .B2(new_n436), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n345), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT81), .B1(new_n458), .B2(new_n343), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n459), .A2(new_n418), .A3(new_n449), .A4(new_n440), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n192), .B1(new_n349), .B2(new_n350), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n356), .A2(new_n318), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n462), .B1(new_n192), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n206), .A2(G224), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n464), .B(new_n465), .Z(new_n466));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n467), .B(new_n419), .C1(new_n450), .C2(new_n454), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n461), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n418), .B(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT84), .B1(new_n446), .B2(new_n436), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT85), .ZN(new_n474));
  INV_X1    g288(.A(new_n380), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n446), .A2(KEYINPUT84), .A3(new_n436), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n473), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n476), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n478), .A2(new_n472), .A3(new_n380), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT85), .B1(new_n448), .B2(new_n475), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n471), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n465), .A2(KEYINPUT7), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n465), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(new_n464), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n463), .A2(new_n192), .ZN(new_n486));
  INV_X1    g300(.A(new_n462), .ZN(new_n487));
  AND4_X1   g301(.A1(new_n486), .A2(new_n487), .A3(new_n482), .A4(new_n484), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n460), .A2(new_n481), .A3(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n490), .A2(new_n293), .ZN(new_n491));
  OAI21_X1  g305(.A(G210), .B1(G237), .B2(G902), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n469), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(new_n469), .B2(new_n491), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n417), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n309), .A2(new_n406), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G234), .ZN(new_n497));
  OAI21_X1  g311(.A(G217), .B1(new_n497), .B2(G902), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT69), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n321), .A2(KEYINPUT64), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT64), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G128), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n502), .A3(G119), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n428), .A2(G128), .ZN(new_n504));
  INV_X1    g318(.A(G110), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT24), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G110), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n503), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT70), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n503), .A2(new_n509), .A3(new_n512), .A4(new_n504), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT23), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n428), .B2(G128), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n504), .B(new_n516), .C1(new_n503), .C2(new_n515), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G110), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n514), .B(new_n518), .C1(new_n199), .C2(new_n203), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n227), .A2(new_n189), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n517), .A2(G110), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n509), .B1(new_n503), .B2(new_n504), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n223), .B(new_n520), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n206), .A2(G221), .A3(G234), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT72), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT22), .B(G137), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n519), .A2(new_n523), .A3(new_n528), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT25), .B1(new_n532), .B2(new_n293), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n519), .A2(new_n523), .A3(new_n528), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n528), .B1(new_n519), .B2(new_n523), .ZN(new_n535));
  OAI211_X1 g349(.A(KEYINPUT25), .B(new_n293), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n499), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT73), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT73), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n540), .B(new_n499), .C1(new_n533), .C2(new_n537), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n499), .A2(G902), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n532), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT74), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n539), .A2(KEYINPUT74), .A3(new_n541), .A4(new_n543), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT32), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n208), .A2(G210), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT27), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT26), .B(G101), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n275), .A2(G137), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n368), .A2(G134), .ZN(new_n556));
  OAI21_X1  g370(.A(G131), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n373), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n356), .B2(new_n318), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n372), .A2(new_n373), .B1(new_n349), .B2(new_n350), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n438), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT28), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT28), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n438), .B1(new_n559), .B2(new_n560), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n374), .A2(new_n351), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n373), .A2(new_n557), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n463), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n566), .A2(new_n568), .A3(new_n434), .A4(new_n437), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n564), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT67), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n563), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n438), .A2(new_n559), .A3(new_n560), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n566), .A2(new_n568), .B1(new_n434), .B2(new_n437), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT28), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT67), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT30), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT30), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n566), .B2(new_n568), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n438), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT66), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n554), .B1(new_n582), .B2(KEYINPUT31), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n569), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n582), .A2(KEYINPUT31), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT30), .B1(new_n559), .B2(new_n560), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n566), .A2(new_n568), .A3(new_n579), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n573), .B1(new_n589), .B2(new_n438), .ZN(new_n590));
  INV_X1    g404(.A(new_n585), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n583), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n554), .A2(new_n577), .B1(new_n586), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(G472), .A2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n549), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n554), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n572), .A2(new_n576), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n581), .A2(new_n569), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT29), .B1(new_n599), .B2(new_n554), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n570), .A2(new_n563), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n597), .A2(KEYINPUT29), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G472), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n586), .A2(new_n592), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n597), .B1(new_n572), .B2(new_n576), .ZN(new_n608));
  OAI211_X1 g422(.A(KEYINPUT32), .B(new_n594), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n596), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT68), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT68), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n596), .A2(new_n606), .A3(new_n609), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n496), .A2(new_n548), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  NAND2_X1  g430(.A1(new_n469), .A2(new_n491), .ZN(new_n617));
  INV_X1    g431(.A(new_n492), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n469), .A2(new_n491), .A3(new_n492), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n469), .A2(new_n491), .A3(KEYINPUT96), .A4(new_n492), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n623), .A2(new_n415), .ZN(new_n624));
  INV_X1    g438(.A(new_n414), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n290), .B2(new_n273), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n292), .A2(new_n627), .B1(new_n628), .B2(new_n285), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n295), .A2(G902), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n629), .A2(new_n630), .B1(new_n295), .B2(new_n294), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n253), .A2(new_n258), .A3(KEYINPUT20), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n308), .A2(new_n302), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n626), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n586), .A2(new_n592), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n571), .B(KEYINPUT28), .C1(new_n573), .C2(new_n574), .ZN(new_n638));
  INV_X1    g452(.A(new_n563), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n570), .A2(new_n571), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n554), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(G472), .ZN(new_n644));
  OAI22_X1  g458(.A1(new_n643), .A2(new_n644), .B1(new_n593), .B2(new_n595), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n406), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n636), .A2(new_n548), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  AND2_X1   g463(.A1(new_n308), .A2(new_n302), .ZN(new_n650));
  INV_X1    g464(.A(new_n300), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n259), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n626), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n548), .A3(new_n646), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NOR2_X1   g470(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n524), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n542), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n539), .A2(new_n541), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n645), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n496), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  INV_X1    g479(.A(new_n310), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n395), .A2(new_n396), .B1(new_n379), .B2(new_n399), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n403), .B1(new_n667), .B2(G469), .ZN(new_n668));
  INV_X1    g482(.A(new_n314), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n399), .B2(new_n394), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n394), .A2(new_n383), .A3(new_n669), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n402), .B(new_n293), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n666), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n673), .A2(new_n622), .A3(new_n624), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n614), .A2(new_n674), .A3(new_n660), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n410), .B1(new_n412), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n652), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XOR2_X1   g494(.A(new_n677), .B(KEYINPUT39), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT40), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT98), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n493), .A2(new_n494), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n651), .B1(new_n633), .B2(new_n634), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n590), .A2(new_n554), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n565), .A2(new_n569), .A3(new_n554), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n293), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n596), .A2(new_n609), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n661), .A2(new_n696), .A3(new_n415), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n690), .A2(new_n691), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n685), .A2(new_n686), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n213), .ZN(G45));
  AOI211_X1 g514(.A(new_n631), .B(new_n677), .C1(new_n650), .C2(new_n259), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n614), .A2(new_n674), .A3(new_n660), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  OAI21_X1  g517(.A(new_n293), .B1(new_n670), .B2(new_n671), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT99), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n672), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n704), .A2(KEYINPUT99), .A3(G469), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n666), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n636), .A2(new_n548), .A3(new_n614), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND4_X1  g526(.A1(new_n653), .A2(new_n548), .A3(new_n614), .A4(new_n709), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT100), .B(G116), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G18));
  INV_X1    g529(.A(new_n309), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n614), .A2(new_n716), .A3(new_n660), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n623), .A2(new_n415), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n687), .B2(new_n620), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n709), .A2(new_n625), .A3(new_n719), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  AOI21_X1  g536(.A(new_n300), .B1(new_n650), .B2(new_n259), .ZN(new_n723));
  INV_X1    g537(.A(new_n544), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n554), .B1(new_n570), .B2(new_n563), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n595), .B1(new_n637), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT101), .B1(new_n643), .B2(new_n644), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT101), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n728), .B(G472), .C1(new_n593), .C2(G902), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n719), .A2(new_n723), .A3(new_n724), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n707), .A2(new_n708), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n625), .A3(new_n310), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT102), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n414), .B(new_n666), .C1(new_n707), .C2(new_n708), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n622), .A2(new_n624), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n691), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n730), .A2(new_n724), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT102), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n735), .A2(new_n737), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  NAND2_X1  g556(.A1(new_n709), .A2(new_n719), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n631), .B1(new_n650), .B2(new_n259), .ZN(new_n744));
  INV_X1    g558(.A(new_n677), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n730), .A3(new_n660), .A4(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT103), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n727), .A2(new_n729), .ZN(new_n748));
  INV_X1    g562(.A(new_n726), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n660), .A3(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n632), .B(new_n745), .C1(new_n633), .C2(new_n634), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT103), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n719), .A4(new_n709), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n747), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  NAND3_X1  g570(.A1(new_n619), .A2(new_n621), .A3(new_n415), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n406), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n548), .A2(new_n614), .A3(new_n701), .A4(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n593), .A2(new_n595), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(KEYINPUT105), .A3(KEYINPUT32), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n609), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n763), .A2(new_n765), .A3(new_n606), .A4(new_n596), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n766), .A2(new_n724), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(KEYINPUT42), .A3(new_n701), .A4(new_n758), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  AND3_X1   g584(.A1(new_n548), .A2(new_n614), .A3(new_n758), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n678), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NAND3_X1  g587(.A1(new_n650), .A2(new_n259), .A3(new_n632), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT43), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT43), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n660), .A2(new_n645), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(KEYINPUT44), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n757), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n667), .A2(KEYINPUT45), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n667), .A2(KEYINPUT45), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(G469), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n404), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n784), .B1(new_n789), .B2(KEYINPUT46), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n385), .B1(new_n789), .B2(KEYINPUT46), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(KEYINPUT106), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n310), .A3(new_n681), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n783), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(new_n368), .ZN(G39));
  NOR4_X1   g611(.A1(new_n548), .A2(new_n614), .A3(new_n751), .A4(new_n757), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n794), .A2(KEYINPUT47), .A3(new_n310), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT47), .B1(new_n794), .B2(new_n310), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT107), .B(G140), .Z(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(G42));
  INV_X1    g617(.A(new_n750), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n493), .A2(new_n494), .A3(new_n416), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n709), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n777), .A2(new_n410), .A3(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n777), .A2(new_n410), .A3(new_n738), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n690), .A2(new_n416), .A3(new_n709), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT50), .ZN(new_n815));
  INV_X1    g629(.A(new_n696), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n807), .A2(new_n548), .A3(new_n410), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n650), .A2(new_n259), .A3(new_n631), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n811), .B(new_n815), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n799), .A2(new_n800), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n732), .A2(new_n666), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n757), .B(new_n812), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n819), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n820), .B1(new_n819), .B2(new_n823), .ZN(new_n825));
  OAI221_X1 g639(.A(new_n407), .B1(new_n817), .B2(new_n635), .C1(new_n812), .C2(new_n743), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n767), .B1(new_n809), .B2(new_n810), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n824), .A2(new_n825), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n635), .A2(new_n652), .ZN(new_n833));
  INV_X1    g647(.A(new_n495), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n548), .A2(new_n833), .A3(new_n834), .A4(new_n646), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n615), .A2(new_n835), .A3(new_n663), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n406), .A2(new_n757), .A3(new_n677), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n804), .A2(new_n837), .A3(new_n838), .A4(new_n744), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n744), .A2(new_n730), .A3(new_n660), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n673), .A2(new_n805), .A3(new_n745), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT111), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n661), .B(new_n309), .C1(new_n611), .C2(new_n613), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n839), .A2(new_n842), .B1(new_n843), .B2(new_n837), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n769), .A2(new_n836), .A3(new_n844), .A4(new_n772), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n539), .A2(new_n541), .A3(new_n659), .A4(new_n745), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n816), .A2(new_n406), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n737), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n850), .A2(new_n702), .ZN(new_n851));
  AND4_X1   g665(.A1(KEYINPUT52), .A2(new_n851), .A3(new_n755), .A4(new_n679), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n754), .A2(new_n747), .B1(new_n675), .B2(new_n678), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(new_n853), .B2(new_n851), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n845), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT110), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n734), .A2(new_n740), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n710), .B(new_n713), .C1(new_n717), .C2(new_n720), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n546), .A2(new_n547), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n613), .B2(new_n611), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n861), .B(new_n709), .C1(new_n636), .C2(new_n653), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n741), .A2(new_n721), .A3(new_n862), .A4(KEYINPUT110), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n832), .B1(new_n855), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n859), .A2(new_n863), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n851), .A2(new_n755), .A3(new_n679), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n853), .A2(KEYINPUT52), .A3(new_n851), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n867), .A2(new_n872), .A3(new_n845), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n832), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT54), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT54), .B1(new_n873), .B2(new_n832), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n852), .A2(new_n854), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n836), .A2(new_n844), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n857), .A2(new_n858), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n761), .A2(new_n768), .B1(new_n678), .B2(new_n771), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT53), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT113), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n769), .A2(new_n836), .A3(new_n844), .A4(new_n772), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n741), .A2(new_n721), .A3(new_n862), .A4(KEYINPUT53), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n872), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n876), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n875), .A2(new_n889), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n831), .A2(new_n890), .B1(G952), .B2(G953), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n774), .A2(new_n544), .A3(new_n416), .A4(new_n666), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT108), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT49), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n892), .A2(new_n893), .B1(new_n894), .B2(new_n732), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n893), .B2(new_n892), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT109), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n732), .A2(new_n894), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n690), .A2(new_n816), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n891), .B1(new_n897), .B2(new_n899), .ZN(G75));
  AND3_X1   g714(.A1(new_n872), .A2(new_n885), .A3(new_n886), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n886), .B1(new_n872), .B2(new_n885), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n865), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(G210), .A2(G902), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT56), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n461), .A2(new_n468), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT115), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n466), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n206), .A2(G952), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n905), .B2(new_n909), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT116), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n905), .A2(new_n909), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT116), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n917), .A3(new_n910), .A4(new_n913), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(G51));
  XNOR2_X1  g733(.A(new_n403), .B(KEYINPUT57), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n876), .A2(new_n888), .A3(KEYINPUT117), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT117), .B1(new_n876), .B2(new_n888), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n378), .A2(new_n384), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n882), .A2(new_n887), .B1(new_n873), .B2(new_n832), .ZN(new_n928));
  OR3_X1    g742(.A1(new_n928), .A2(new_n293), .A3(new_n787), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n912), .B1(new_n927), .B2(new_n929), .ZN(G54));
  NAND4_X1  g744(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n931), .A2(new_n256), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n256), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n912), .ZN(G60));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n875), .B2(new_n889), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n913), .B1(new_n937), .B2(new_n629), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n923), .A2(new_n924), .ZN(new_n939));
  INV_X1    g753(.A(new_n936), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n629), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n939), .B2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT60), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n531), .B(new_n530), .C1(new_n928), .C2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n944), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n903), .A2(new_n658), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n913), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT118), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n949), .A3(new_n913), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT61), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n944), .B1(new_n888), .B2(new_n865), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n912), .B1(new_n952), .B2(new_n658), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n953), .B(new_n945), .C1(new_n949), .C2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n951), .A2(new_n955), .ZN(G66));
  INV_X1    g770(.A(G224), .ZN(new_n957));
  OAI21_X1  g771(.A(G953), .B1(new_n413), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n867), .A2(new_n836), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT119), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT119), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n867), .A2(new_n961), .A3(new_n836), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n958), .B1(new_n963), .B2(G953), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n907), .B1(G898), .B2(new_n206), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(G69));
  XNOR2_X1  g780(.A(new_n589), .B(new_n245), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n783), .A2(new_n795), .ZN(new_n968));
  INV_X1    g782(.A(new_n771), .ZN(new_n969));
  INV_X1    g783(.A(new_n833), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n970), .A2(KEYINPUT120), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(KEYINPUT120), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n681), .A3(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n801), .B(new_n968), .C1(new_n969), .C2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n853), .A2(new_n702), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n699), .B2(new_n976), .ZN(new_n977));
  OR3_X1    g791(.A1(new_n699), .A2(new_n976), .A3(new_n975), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n967), .B1(new_n979), .B2(G953), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT121), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(KEYINPUT121), .B(new_n967), .C1(new_n979), .C2(G953), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n968), .A2(KEYINPUT122), .A3(new_n702), .A4(new_n853), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT122), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n796), .B2(new_n976), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n880), .A2(KEYINPUT123), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n880), .A2(KEYINPUT123), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n767), .A2(new_n737), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n795), .A2(new_n990), .ZN(new_n991));
  AND4_X1   g805(.A1(new_n801), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n987), .A2(new_n206), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n967), .B1(G900), .B2(G953), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n982), .A2(new_n983), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n206), .B1(G227), .B2(G900), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT124), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n996), .B(new_n999), .ZN(G72));
  INV_X1    g814(.A(new_n692), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n979), .A2(new_n962), .A3(new_n960), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT63), .Z(new_n1004));
  AOI21_X1  g818(.A(new_n1001), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n866), .A2(new_n874), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n590), .A2(new_n554), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1001), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1005), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n987), .A2(new_n960), .A3(new_n962), .A4(new_n992), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1011), .A2(new_n1004), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1007), .B(KEYINPUT125), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1010), .B(new_n913), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1014), .B1(new_n1011), .B2(new_n1004), .ZN(new_n1016));
  OAI21_X1  g830(.A(KEYINPUT126), .B1(new_n1016), .B2(new_n912), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n1009), .A2(new_n1015), .A3(new_n1017), .ZN(G57));
endmodule


