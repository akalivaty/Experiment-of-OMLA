//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT80), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT9), .B(G234), .ZN(new_n190));
  OAI21_X1  g004(.A(G221), .B1(new_n190), .B2(G902), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G469), .ZN(new_n193));
  INV_X1    g007(.A(G902), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT0), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT0), .B(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT78), .B(G101), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G104), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n207), .A2(new_n209), .A3(new_n210), .A4(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n213), .A3(new_n210), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n214), .A2(KEYINPUT4), .B1(new_n215), .B2(G101), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n215), .A2(KEYINPUT4), .A3(G101), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n206), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(G137), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT11), .A3(G134), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(G137), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n221), .A2(new_n223), .A3(new_n227), .A4(new_n224), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n210), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n208), .A2(G107), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n214), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n202), .B1(KEYINPUT1), .B2(new_n197), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n203), .A2(new_n197), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(KEYINPUT10), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT10), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n203), .A2(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n242), .A2(new_n235), .B1(new_n197), .B2(new_n203), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n214), .A2(new_n233), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n240), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n218), .A2(new_n230), .A3(new_n239), .A4(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G110), .B(G140), .ZN(new_n247));
  INV_X1    g061(.A(G227), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G953), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n247), .B(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT79), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n234), .A2(new_n238), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n243), .A2(new_n244), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT12), .B1(new_n256), .B2(new_n229), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT12), .ZN(new_n258));
  AOI211_X1 g072(.A(new_n258), .B(new_n230), .C1(new_n254), .C2(new_n255), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT79), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n246), .B2(new_n251), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n253), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n218), .A2(new_n245), .A3(new_n239), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n229), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n251), .B1(new_n265), .B2(new_n246), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n193), .B(new_n194), .C1(new_n263), .C2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n193), .A2(new_n194), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n246), .B1(new_n257), .B2(new_n259), .ZN(new_n269));
  INV_X1    g083(.A(new_n252), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n269), .A2(new_n250), .B1(new_n270), .B2(new_n265), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n268), .B1(new_n271), .B2(G469), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n192), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n274));
  AND2_X1   g088(.A1(KEYINPUT65), .A2(G119), .ZN(new_n275));
  NOR2_X1   g089(.A1(KEYINPUT65), .A2(G119), .ZN(new_n276));
  OAI21_X1  g090(.A(G116), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT2), .B(G113), .ZN(new_n278));
  NOR2_X1   g092(.A1(G116), .A2(G119), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n278), .B1(new_n277), .B2(new_n280), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n274), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n280), .ZN(new_n284));
  INV_X1    g098(.A(new_n278), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(KEYINPUT66), .A3(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n283), .B(new_n288), .C1(new_n216), .C2(new_n217), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n284), .A2(KEYINPUT5), .ZN(new_n291));
  INV_X1    g105(.A(G116), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(KEYINPUT5), .ZN(new_n293));
  OR2_X1    g107(.A1(KEYINPUT65), .A2(G119), .ZN(new_n294));
  NAND2_X1  g108(.A1(KEYINPUT65), .A2(G119), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT81), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n293), .A2(new_n294), .A3(new_n298), .A4(new_n295), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(G113), .A3(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n286), .B(new_n234), .C1(new_n291), .C2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n289), .A2(new_n290), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G110), .B(G122), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n303), .B(KEYINPUT83), .Z(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n290), .B1(new_n289), .B2(new_n301), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n289), .A2(new_n301), .A3(new_n303), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT6), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT84), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n206), .A2(G125), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(G125), .B2(new_n243), .ZN(new_n312));
  INV_X1    g126(.A(G953), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G224), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n312), .B(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n308), .A2(KEYINPUT6), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT84), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n316), .B(new_n317), .C1(new_n306), .C2(new_n305), .ZN(new_n318));
  OR3_X1    g132(.A1(new_n305), .A2(KEYINPUT6), .A3(new_n306), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n310), .A2(new_n315), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G210), .B1(G237), .B2(G902), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(KEYINPUT7), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n312), .B(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n323), .A2(new_n308), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n303), .B(KEYINPUT8), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n291), .A2(new_n300), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n244), .A2(new_n286), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT85), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n291), .B1(new_n300), .B2(new_n328), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n300), .A2(new_n328), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n282), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI221_X1 g145(.A(new_n325), .B1(new_n326), .B2(new_n327), .C1(new_n331), .C2(new_n244), .ZN(new_n332));
  AOI21_X1  g146(.A(G902), .B1(new_n324), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n320), .A2(new_n321), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n321), .B1(new_n320), .B2(new_n333), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n189), .B(new_n273), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n338));
  XNOR2_X1  g152(.A(G113), .B(G122), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(new_n208), .ZN(new_n340));
  INV_X1    g154(.A(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G140), .ZN(new_n342));
  INV_X1    g156(.A(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G125), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT76), .ZN(new_n345));
  OR3_X1    g159(.A1(new_n343), .A2(KEYINPUT76), .A3(G125), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT19), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT86), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT86), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n345), .A2(new_n346), .A3(new_n350), .A4(KEYINPUT19), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n348), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n349), .A2(new_n199), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n344), .A2(KEYINPUT16), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n343), .A2(KEYINPUT76), .A3(G125), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n352), .B2(KEYINPUT76), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT16), .ZN(new_n359));
  OAI211_X1 g173(.A(G146), .B(new_n356), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(G237), .A2(G953), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G143), .A3(G214), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(G143), .B1(new_n361), .B2(G214), .ZN(new_n364));
  OAI21_X1  g178(.A(G131), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(G214), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n201), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n227), .A3(new_n362), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n354), .A2(new_n360), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n362), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(KEYINPUT18), .A3(G131), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n352), .A2(new_n199), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n347), .B2(new_n199), .ZN(new_n374));
  NAND2_X1  g188(.A1(KEYINPUT18), .A2(G131), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n367), .A2(new_n362), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n340), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT17), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n365), .A2(new_n379), .A3(new_n368), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n359), .B1(new_n345), .B2(new_n346), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n199), .B1(new_n381), .B2(new_n355), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n371), .A2(KEYINPUT17), .A3(G131), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n380), .A2(new_n382), .A3(new_n360), .A4(new_n383), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n384), .A2(new_n377), .A3(new_n340), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n338), .B1(new_n378), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(G475), .A2(G902), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n377), .A3(new_n340), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n360), .A2(new_n369), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n372), .A2(new_n376), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n389), .A2(new_n354), .B1(new_n390), .B2(new_n374), .ZN(new_n391));
  OAI211_X1 g205(.A(KEYINPUT87), .B(new_n388), .C1(new_n391), .C2(new_n340), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n387), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n388), .B1(new_n391), .B2(new_n340), .ZN(new_n394));
  NOR3_X1   g208(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n393), .A2(KEYINPUT20), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n340), .B1(new_n384), .B2(new_n377), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n194), .B1(new_n385), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G475), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(G234), .A2(G237), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(G952), .A3(new_n313), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT21), .B(G898), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(G902), .A3(G953), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT88), .B1(new_n201), .B2(G128), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT88), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n197), .A3(G143), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n201), .A2(G128), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n412), .A2(new_n220), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n220), .B1(new_n412), .B2(new_n413), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n408), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n292), .A2(G122), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n292), .A2(G122), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n418), .A2(new_n419), .A3(new_n212), .ZN(new_n420));
  INV_X1    g234(.A(G122), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n421), .A2(KEYINPUT14), .A3(G116), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(new_n417), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT90), .B1(new_n419), .B2(KEYINPUT14), .ZN(new_n424));
  OAI211_X1 g238(.A(KEYINPUT90), .B(KEYINPUT14), .C1(new_n421), .C2(G116), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n423), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n420), .B1(new_n427), .B2(G107), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n410), .B1(new_n197), .B2(G143), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n201), .A2(KEYINPUT88), .A3(G128), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n413), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G134), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n412), .A2(new_n220), .A3(new_n413), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(KEYINPUT89), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n416), .A2(new_n428), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT13), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n413), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n412), .ZN(new_n438));
  OAI21_X1  g252(.A(G134), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n212), .B1(new_n418), .B2(new_n419), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n439), .B(new_n433), .C1(new_n440), .C2(new_n420), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G217), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n190), .A2(new_n443), .A3(G953), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT91), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n435), .A2(new_n441), .A3(new_n444), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n442), .A2(KEYINPUT91), .A3(new_n445), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n194), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G478), .B1(KEYINPUT92), .B2(KEYINPUT15), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(KEYINPUT92), .B2(KEYINPUT15), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n451), .A2(new_n453), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n401), .A2(new_n407), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n283), .A2(new_n288), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n220), .A2(G137), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n222), .A2(G134), .ZN(new_n462));
  OAI21_X1  g276(.A(G131), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n228), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n238), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n226), .A2(new_n228), .B1(new_n198), .B2(new_n205), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT30), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n238), .B2(new_n464), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT67), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n229), .A2(new_n206), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n469), .B2(new_n471), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n459), .B(new_n467), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT26), .B(G101), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT69), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(G210), .A3(new_n361), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n475), .B(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n361), .A2(G210), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n478), .A2(new_n481), .A3(new_n483), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n238), .A2(new_n464), .B1(new_n229), .B2(new_n206), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n458), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n474), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT70), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT70), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n474), .A2(new_n491), .A3(new_n488), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(KEYINPUT31), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT31), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n474), .A2(new_n494), .A3(new_n488), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT71), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n474), .A2(KEYINPUT71), .A3(new_n488), .A4(new_n494), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n458), .A2(new_n487), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT72), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT72), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n503), .B(KEYINPUT28), .C1(new_n458), .C2(new_n487), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n458), .B(new_n487), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT28), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n485), .A2(new_n486), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n493), .A2(new_n499), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(G472), .A2(G902), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT32), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n505), .A2(new_n507), .A3(new_n509), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT73), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT73), .A4(new_n509), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n509), .B1(new_n474), .B2(new_n500), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(KEYINPUT29), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n500), .A2(new_n501), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n503), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT74), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n500), .A2(KEYINPUT72), .A3(new_n501), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT74), .B1(new_n502), .B2(new_n504), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n507), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n509), .A2(KEYINPUT29), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n194), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G472), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n512), .A2(KEYINPUT32), .A3(new_n513), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n516), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n313), .A2(G221), .A3(G234), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT22), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(G137), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n382), .A2(new_n360), .ZN(new_n539));
  OAI21_X1  g353(.A(G128), .B1(new_n275), .B2(new_n276), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n540), .B(KEYINPUT23), .C1(G119), .C2(G128), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n197), .B1(new_n275), .B2(new_n276), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT23), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G110), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT75), .ZN(new_n547));
  NOR2_X1   g361(.A1(G119), .A2(G128), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n294), .A2(new_n295), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n549), .B2(G128), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT24), .B(G110), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n540), .B1(G119), .B2(G128), .ZN(new_n553));
  INV_X1    g367(.A(new_n551), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(KEYINPUT75), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n539), .A2(new_n546), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G110), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n541), .A2(new_n558), .A3(new_n544), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n550), .A2(new_n551), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n360), .A3(new_n373), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n557), .A2(new_n562), .A3(KEYINPUT77), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT77), .B1(new_n557), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n538), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n557), .A2(new_n562), .A3(KEYINPUT77), .ZN(new_n566));
  INV_X1    g380(.A(new_n538), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT25), .B1(new_n569), .B2(G902), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n443), .B1(G234), .B2(new_n194), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n565), .A2(new_n572), .A3(new_n194), .A4(new_n568), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n552), .A2(new_n555), .B1(new_n545), .B2(G110), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n360), .A2(new_n373), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n575), .A2(new_n539), .B1(new_n576), .B2(new_n561), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n538), .B1(new_n577), .B2(KEYINPUT77), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n557), .A2(new_n562), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT77), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n566), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n578), .B1(new_n582), .B2(new_n538), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n571), .A2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n574), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n337), .A2(new_n457), .A3(new_n535), .A4(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n587), .B(new_n207), .Z(G3));
  INV_X1    g402(.A(new_n187), .ZN(new_n589));
  INV_X1    g403(.A(new_n335), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n320), .A2(new_n321), .A3(new_n333), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n393), .A2(KEYINPUT20), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n394), .A2(new_n395), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n399), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n449), .A2(new_n597), .A3(new_n450), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT93), .B1(new_n442), .B2(new_n445), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT93), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n600), .B(new_n444), .C1(new_n435), .C2(new_n441), .ZN(new_n601));
  OAI211_X1 g415(.A(KEYINPUT33), .B(new_n448), .C1(new_n599), .C2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G478), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G902), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n598), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n451), .A2(new_n603), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n596), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n592), .A2(new_n407), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n512), .A2(new_n194), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G472), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n612), .A2(new_n586), .A3(new_n273), .A4(new_n514), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  AOI21_X1  g430(.A(new_n400), .B1(new_n455), .B2(new_n454), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n386), .A2(new_n392), .A3(new_n395), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT94), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n386), .A2(new_n620), .A3(new_n392), .A4(new_n395), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n593), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n592), .A2(new_n407), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n613), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT95), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT35), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G107), .ZN(G9));
  NOR2_X1   g443(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n579), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n584), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n572), .B1(new_n583), .B2(new_n194), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n573), .A2(new_n571), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n574), .A2(KEYINPUT96), .A3(new_n632), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n456), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G472), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n512), .B2(new_n194), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n513), .B2(new_n512), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n337), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  NAND2_X1  g459(.A1(new_n267), .A2(new_n272), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n191), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n637), .B2(new_n638), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n535), .A2(new_n648), .A3(new_n592), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n403), .B1(new_n406), .B2(G900), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n617), .A2(new_n623), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT97), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n197), .ZN(G30));
  NAND2_X1  g469(.A1(new_n590), .A2(new_n591), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT38), .Z(new_n657));
  NAND2_X1  g471(.A1(new_n637), .A2(new_n638), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n455), .A2(new_n454), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n596), .A2(new_n187), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT98), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n474), .A2(new_n491), .A3(new_n488), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n491), .B1(new_n474), .B2(new_n488), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n510), .A2(new_n506), .ZN(new_n666));
  AOI21_X1  g480(.A(G902), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(new_n640), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n516), .A2(new_n534), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n650), .B(KEYINPUT39), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n273), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT40), .ZN(new_n673));
  OR4_X1    g487(.A1(new_n657), .A2(new_n662), .A3(new_n670), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  OAI211_X1 g489(.A(new_n607), .B(new_n650), .C1(new_n396), .C2(new_n400), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n596), .A2(KEYINPUT99), .A3(new_n607), .A4(new_n650), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(new_n535), .A3(new_n592), .A4(new_n648), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  NOR2_X1   g496(.A1(new_n260), .A2(new_n262), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n270), .A2(new_n261), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n266), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(G469), .B1(new_n685), .B2(G902), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n267), .A3(new_n191), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n267), .A3(KEYINPUT100), .A4(new_n191), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n535), .A3(new_n586), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n610), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT41), .B(G113), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  AND3_X1   g509(.A1(new_n592), .A2(new_n407), .A3(new_n624), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n574), .A2(new_n585), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n512), .A2(KEYINPUT32), .A3(new_n513), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT32), .B1(new_n512), .B2(new_n513), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n697), .B1(new_n700), .B2(new_n533), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n696), .A2(new_n701), .A3(new_n702), .A4(new_n691), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT101), .B1(new_n692), .B2(new_n625), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT102), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NAND2_X1  g521(.A1(new_n639), .A2(new_n535), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n709));
  INV_X1    g523(.A(new_n687), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n592), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n710), .B(new_n187), .C1(new_n334), .C2(new_n335), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT103), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n708), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n714), .B(G119), .Z(G21));
  AND3_X1   g529(.A1(new_n689), .A2(new_n407), .A3(new_n690), .ZN(new_n716));
  INV_X1    g530(.A(new_n513), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n530), .A2(KEYINPUT104), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n528), .A2(new_n529), .A3(new_n719), .A4(new_n507), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n510), .A3(new_n720), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n665), .A2(KEYINPUT31), .B1(new_n497), .B2(new_n498), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n717), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n723), .A2(new_n641), .A3(new_n697), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n660), .B1(new_n590), .B2(new_n591), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n716), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NOR2_X1   g541(.A1(new_n723), .A2(new_n641), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n658), .A3(new_n678), .A4(new_n679), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n711), .B2(new_n713), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n341), .ZN(G27));
  XNOR2_X1  g545(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n334), .A2(new_n335), .A3(new_n589), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n535), .A2(new_n734), .A3(new_n273), .A4(new_n586), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n678), .A2(new_n679), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n590), .A2(new_n591), .A3(new_n187), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n647), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(KEYINPUT42), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n701), .A2(new_n680), .A3(new_n739), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NOR2_X1   g559(.A1(new_n735), .A2(new_n653), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT106), .B(G134), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G36));
  NAND2_X1  g562(.A1(new_n401), .A2(new_n607), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT108), .Z(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n750), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT107), .Z(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n642), .B1(new_n637), .B2(new_n638), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(KEYINPUT44), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT44), .B1(new_n755), .B2(new_n756), .ZN(new_n760));
  OAI21_X1  g574(.A(G469), .B1(new_n271), .B2(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(KEYINPUT45), .B2(new_n271), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n268), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n267), .B1(new_n763), .B2(KEYINPUT46), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n191), .B(new_n671), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n760), .A2(new_n738), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  OAI21_X1  g583(.A(new_n191), .B1(new_n764), .B2(new_n765), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT47), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n700), .A2(new_n533), .A3(new_n697), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n771), .A2(new_n736), .A3(new_n738), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n343), .ZN(G42));
  NAND2_X1  g588(.A1(new_n734), .A2(new_n710), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n775), .A2(KEYINPUT118), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n403), .B1(new_n775), .B2(KEYINPUT118), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n755), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n701), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT48), .Z(new_n781));
  AND4_X1   g595(.A1(new_n586), .A2(new_n776), .A3(new_n670), .A4(new_n777), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n609), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n728), .A2(new_n586), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n403), .B(new_n784), .C1(new_n752), .C2(new_n754), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n711), .A2(new_n713), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT119), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n313), .A2(G952), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n787), .B2(KEYINPUT119), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n781), .A2(new_n783), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n686), .A2(new_n267), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n191), .B1(new_n792), .B2(KEYINPUT116), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(KEYINPUT116), .B2(new_n792), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n771), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n785), .A2(new_n795), .A3(new_n734), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT117), .Z(new_n797));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n728), .A2(new_n658), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n778), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n596), .A2(new_n607), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n800), .B1(new_n782), .B2(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n657), .A2(new_n589), .A3(new_n710), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n785), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n797), .A2(new_n798), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n802), .A3(new_n796), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n791), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n587), .A2(new_n643), .A3(new_n726), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n692), .ZN(new_n814));
  INV_X1    g628(.A(new_n610), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n656), .A2(new_n189), .A3(new_n407), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n613), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n608), .A2(KEYINPUT110), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n596), .A2(new_n819), .A3(new_n607), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n401), .A2(new_n822), .A3(new_n659), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n401), .B2(new_n659), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n814), .A2(new_n815), .B1(new_n817), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n714), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n705), .A2(new_n813), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n535), .A2(new_n648), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n399), .A2(new_n650), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n832), .B(new_n659), .C1(new_n593), .C2(new_n622), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n831), .A3(new_n734), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n535), .A2(new_n648), .A3(new_n833), .A4(new_n734), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT112), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n734), .A2(new_n273), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n735), .A2(new_n653), .B1(new_n729), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n744), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n829), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n574), .A2(new_n632), .A3(new_n650), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n844), .B2(new_n647), .ZN(new_n845));
  INV_X1    g659(.A(new_n635), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(KEYINPUT113), .A3(new_n273), .A4(new_n650), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n725), .A2(new_n669), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n681), .B(new_n848), .C1(new_n653), .C2(new_n649), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT114), .B1(new_n849), .B2(new_n730), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n651), .B(KEYINPUT97), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n830), .B(new_n592), .C1(new_n851), .C2(new_n680), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n799), .A2(new_n736), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n786), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n852), .A2(new_n854), .A3(new_n855), .A4(new_n848), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT52), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n849), .A2(new_n858), .A3(new_n730), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n842), .B(KEYINPUT53), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n826), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n188), .B1(new_n590), .B2(new_n591), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n647), .A2(new_n697), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n642), .A2(new_n862), .A3(new_n407), .A4(new_n863), .ZN(new_n864));
  OAI22_X1  g678(.A1(new_n861), .A2(new_n864), .B1(new_n692), .B2(new_n610), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n865), .A2(new_n812), .A3(new_n714), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n839), .B1(new_n834), .B2(new_n836), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n705), .A3(new_n867), .A4(new_n744), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n850), .A2(new_n856), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n858), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n850), .A2(KEYINPUT52), .A3(new_n856), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n811), .B(new_n860), .C1(new_n872), .C2(KEYINPUT53), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n850), .A2(KEYINPUT52), .A3(new_n856), .ZN(new_n876));
  OAI211_X1 g690(.A(KEYINPUT53), .B(new_n842), .C1(new_n876), .C2(new_n857), .ZN(new_n877));
  INV_X1    g691(.A(new_n859), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n868), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n879), .B2(KEYINPUT53), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT54), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n842), .B1(new_n876), .B2(new_n857), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(KEYINPUT115), .A3(new_n811), .A4(new_n860), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n810), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(G952), .B2(G953), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n792), .B(KEYINPUT49), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n889), .A2(new_n188), .A3(new_n192), .A4(new_n749), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n657), .A2(new_n890), .A3(new_n586), .A4(new_n670), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n891), .ZN(G75));
  AOI21_X1  g706(.A(new_n194), .B1(new_n885), .B2(new_n860), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(G210), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n310), .A2(new_n318), .A3(new_n319), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n315), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT55), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n894), .B2(new_n895), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n313), .A2(G952), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT120), .Z(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(G51));
  NAND2_X1  g718(.A1(new_n873), .A2(KEYINPUT121), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n885), .A2(new_n906), .A3(new_n811), .A4(new_n860), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n860), .B1(new_n872), .B2(KEYINPUT53), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n268), .B(KEYINPUT57), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n266), .B2(new_n263), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n893), .A2(new_n762), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n901), .B1(new_n913), .B2(new_n914), .ZN(G54));
  NAND2_X1  g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT122), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n893), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n386), .A2(new_n392), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n918), .A2(new_n919), .B1(G952), .B2(new_n313), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n919), .B2(new_n918), .ZN(G60));
  AND2_X1   g735(.A1(new_n598), .A2(new_n602), .ZN(new_n922));
  XNOR2_X1  g736(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n603), .A2(new_n194), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n903), .B1(new_n910), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n875), .A2(new_n886), .A3(new_n881), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n922), .B1(new_n928), .B2(new_n925), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI211_X1 g745(.A(KEYINPUT124), .B(new_n922), .C1(new_n928), .C2(new_n925), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(G63));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT60), .Z(new_n935));
  NAND2_X1  g749(.A1(new_n908), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n631), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n902), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT61), .B1(new_n938), .B2(KEYINPUT125), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n569), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n940), .B(new_n902), .C1(new_n937), .C2(new_n936), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G66));
  NAND2_X1  g756(.A1(new_n829), .A2(new_n313), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT126), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n313), .B1(new_n405), .B2(G224), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n896), .B1(G898), .B2(new_n313), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n946), .B(new_n947), .Z(G69));
  OAI21_X1  g762(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT127), .Z(new_n951));
  XNOR2_X1  g765(.A(new_n949), .B(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n725), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n766), .A2(new_n779), .A3(new_n953), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n773), .A2(new_n746), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n852), .A2(new_n854), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n955), .A2(new_n768), .A3(new_n744), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n313), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n248), .A2(G900), .A3(G953), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n952), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n674), .A2(new_n956), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n773), .B1(new_n962), .B2(KEYINPUT62), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(KEYINPUT62), .B2(new_n962), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n701), .A2(new_n826), .A3(new_n671), .A4(new_n739), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n768), .A2(new_n313), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n961), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n960), .B1(new_n967), .B2(new_n952), .ZN(G72));
  NAND2_X1  g782(.A1(G472), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT63), .Z(new_n970));
  NAND4_X1  g784(.A1(new_n768), .A2(new_n705), .A3(new_n866), .A4(new_n965), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n964), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n474), .A2(new_n500), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n509), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n970), .B1(new_n957), .B2(new_n829), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n973), .A2(new_n509), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n901), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n665), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n880), .B(new_n970), .C1(new_n978), .C2(new_n521), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n974), .A2(new_n977), .A3(new_n979), .ZN(G57));
endmodule


